magic
tech scmos
timestamp 1394680314
<< m1p >>
use CELL  1
transform -1 0 1885 0 1 1740
box 0 0 6 6
use CELL  2
transform 1 0 1792 0 1 1908
box 0 0 6 6
use CELL  3
transform 1 0 1910 0 1 1668
box 0 0 6 6
use CELL  4
transform 1 0 1731 0 1 1704
box 0 0 6 6
use CELL  5
transform 1 0 1793 0 1 1848
box 0 0 6 6
use CELL  6
transform 1 0 1929 0 1 1704
box 0 0 6 6
use CELL  7
transform 1 0 1942 0 1 1812
box 0 0 6 6
use CELL  8
transform 1 0 1943 0 1 1752
box 0 0 6 6
use CELL  9
transform 1 0 1738 0 -1 1830
box 0 0 6 6
use CELL  10
transform 1 0 1801 0 1 1932
box 0 0 6 6
use CELL  11
transform 1 0 1947 0 1 1716
box 0 0 6 6
use CELL  12
transform 1 0 1866 0 1 1920
box 0 0 6 6
use CELL  13
transform -1 0 1785 0 1 1776
box 0 0 6 6
use CELL  14
transform 1 0 1921 0 1 1812
box 0 0 6 6
use CELL  15
transform 1 0 1816 0 -1 1950
box 0 0 6 6
use CELL  16
transform 1 0 1767 0 -1 1794
box 0 0 6 6
use CELL  17
transform 1 0 1813 0 1 1692
box 0 0 6 6
use CELL  18
transform 1 0 1846 0 1 1812
box 0 0 6 6
use CELL  19
transform 1 0 1799 0 1 1692
box 0 0 6 6
use CELL  20
transform -1 0 1923 0 -1 1782
box 0 0 6 6
use CELL  21
transform 1 0 1852 0 1 1920
box 0 0 6 6
use CELL  22
transform -1 0 1941 0 1 1836
box 0 0 6 6
use CELL  23
transform 1 0 1839 0 1 1776
box 0 0 6 6
use CELL  24
transform -1 0 1752 0 -1 1782
box 0 0 6 6
use CELL  25
transform 1 0 1836 0 1 1932
box 0 0 6 6
use CELL  26
transform 1 0 1792 0 1 1932
box 0 0 6 6
use CELL  27
transform -1 0 1734 0 -1 1674
box 0 0 6 6
use CELL  28
transform 1 0 1887 0 -1 1878
box 0 0 6 6
use CELL  29
transform 1 0 1814 0 1 1836
box 0 0 6 6
use CELL  30
transform 1 0 1762 0 1 1920
box 0 0 6 6
use CELL  31
transform 1 0 1794 0 -1 1650
box 0 0 6 6
use CELL  32
transform 1 0 1791 0 -1 1818
box 0 0 6 6
use CELL  33
transform 1 0 1792 0 1 1920
box 0 0 6 6
use CELL  34
transform 1 0 1829 0 1 1920
box 0 0 6 6
use CELL  35
transform 1 0 1845 0 1 1920
box 0 0 6 6
use CELL  36
transform -1 0 1976 0 1 1776
box 0 0 6 6
use CELL  37
transform 1 0 1924 0 1 1776
box 0 0 6 6
use CELL  38
transform -1 0 1848 0 -1 1854
box 0 0 6 6
use CELL  39
transform -1 0 1746 0 1 1812
box 0 0 6 6
use CELL  40
transform -1 0 1922 0 -1 1758
box 0 0 6 6
use CELL  41
transform 1 0 1903 0 1 1920
box 0 0 6 6
use CELL  42
transform 1 0 1734 0 1 1872
box 0 0 6 6
use CELL  43
transform 1 0 1860 0 1 1704
box 0 0 6 6
use CELL  44
transform -1 0 1957 0 1 1728
box 0 0 6 6
use CELL  45
transform 1 0 1821 0 1 1872
box 0 0 6 6
use CELL  46
transform -1 0 1788 0 -1 1890
box 0 0 6 6
use CELL  47
transform 1 0 1761 0 1 1824
box 0 0 6 6
use CELL  48
transform 1 0 1771 0 1 1704
box 0 0 6 6
use CELL  49
transform 1 0 1852 0 1 1836
box 0 0 6 6
use CELL  50
transform -1 0 1793 0 1 1728
box 0 0 6 6
use CELL  51
transform -1 0 1833 0 1 1656
box 0 0 6 6
use CELL  52
transform -1 0 1875 0 -1 1722
box 0 0 6 6
use CELL  53
transform 1 0 1753 0 1 1656
box 0 0 6 6
use CELL  54
transform 1 0 1799 0 1 1704
box 0 0 6 6
use CELL  55
transform -1 0 1959 0 1 1800
box 0 0 6 6
use CELL  56
transform -1 0 1938 0 1 1800
box 0 0 6 6
use CELL  57
transform 1 0 1882 0 1 1704
box 0 0 6 6
use CELL  58
transform 1 0 1755 0 1 1920
box 0 0 6 6
use CELL  59
transform -1 0 1799 0 1 1860
box 0 0 6 6
use CELL  60
transform 1 0 1859 0 1 1908
box 0 0 6 6
use CELL  61
transform -1 0 1747 0 -1 1950
box 0 0 6 6
use CELL  62
transform -1 0 1913 0 1 1800
box 0 0 6 6
use CELL  63
transform -1 0 1946 0 -1 1854
box 0 0 6 6
use CELL  64
transform -1 0 2022 0 1 1812
box 0 0 6 6
use CELL  65
transform 1 0 1769 0 1 1920
box 0 0 6 6
use CELL  66
transform 1 0 1916 0 -1 1734
box 0 0 6 6
use CELL  67
transform 1 0 1808 0 1 1824
box 0 0 6 6
use CELL  68
transform 1 0 1896 0 1 1908
box 0 0 6 6
use CELL  69
transform 1 0 1894 0 1 1896
box 0 0 6 6
use CELL  70
transform 1 0 1893 0 1 1884
box 0 0 6 6
use CELL  71
transform 1 0 1741 0 1 1884
box 0 0 6 6
use CELL  72
transform 1 0 1908 0 1 1704
box 0 0 6 6
use CELL  73
transform -1 0 1843 0 1 1800
box 0 0 6 6
use CELL  74
transform -1 0 1973 0 1 1764
box 0 0 6 6
use CELL  75
transform 1 0 1795 0 1 1668
box 0 0 6 6
use CELL  76
transform 1 0 1802 0 1 1668
box 0 0 6 6
use CELL  77
transform 1 0 1758 0 1 1668
box 0 0 6 6
use CELL  78
transform -1 0 1741 0 1 1740
box 0 0 6 6
use CELL  79
transform -1 0 1824 0 -1 1758
box 0 0 6 6
use CELL  80
transform 1 0 1834 0 1 1668
box 0 0 6 6
use CELL  81
transform 1 0 1776 0 1 1908
box 0 0 6 6
use CELL  82
transform 1 0 1741 0 1 1848
box 0 0 6 6
use CELL  83
transform 1 0 1901 0 1 1704
box 0 0 6 6
use CELL  84
transform -1 0 1789 0 1 1788
box 0 0 6 6
use CELL  85
transform -1 0 1761 0 -1 1878
box 0 0 6 6
use CELL  86
transform -1 0 1869 0 -1 1794
box 0 0 6 6
use CELL  87
transform 1 0 1872 0 1 1824
box 0 0 6 6
use CELL  88
transform 1 0 1796 0 1 1752
box 0 0 6 6
use CELL  89
transform -1 0 1734 0 1 1788
box 0 0 6 6
use CELL  90
transform 1 0 1693 0 -1 1902
box 0 0 6 6
use CELL  91
transform 1 0 1956 0 1 1776
box 0 0 6 6
use CELL  92
transform 1 0 1946 0 1 1764
box 0 0 6 6
use CELL  93
transform 1 0 1887 0 1 1896
box 0 0 6 6
use CELL  94
transform -1 0 1971 0 1 1740
box 0 0 6 6
use CELL  95
transform 1 0 1922 0 1 1704
box 0 0 6 6
use CELL  96
transform 1 0 1922 0 1 1692
box 0 0 6 6
use CELL  97
transform 1 0 1904 0 1 1680
box 0 0 6 6
use CELL  98
transform 1 0 1836 0 1 1740
box 0 0 6 6
use CELL  99
transform -1 0 1692 0 -1 1902
box 0 0 6 6
use CELL  100
transform -1 0 1959 0 1 1860
box 0 0 6 6
use CELL  101
transform -1 0 1920 0 1 1860
box 0 0 6 6
use CELL  102
transform 1 0 1821 0 1 1848
box 0 0 6 6
use CELL  103
transform -1 0 1830 0 1 1644
box 0 0 6 6
use CELL  104
transform 1 0 1941 0 -1 1806
box 0 0 6 6
use CELL  105
transform -1 0 1801 0 -1 1950
box 0 0 6 6
use CELL  106
transform 1 0 1758 0 1 1752
box 0 0 6 6
use CELL  107
transform -1 0 1978 0 -1 1830
box 0 0 6 6
use CELL  108
transform 1 0 1983 0 1 1800
box 0 0 6 6
use CELL  109
transform 1 0 1866 0 1 1908
box 0 0 6 6
use CELL  110
transform 1 0 1946 0 1 1824
box 0 0 6 6
use CELL  111
transform 1 0 1801 0 1 1908
box 0 0 6 6
use CELL  112
transform 1 0 1925 0 -1 1830
box 0 0 6 6
use CELL  113
transform 1 0 1749 0 1 1740
box 0 0 6 6
use CELL  114
transform -1 0 2008 0 -1 1794
box 0 0 6 6
use CELL  115
transform -1 0 1939 0 1 1776
box 0 0 6 6
use CELL  116
transform 1 0 1974 0 1 1800
box 0 0 6 6
use CELL  117
transform -1 0 1754 0 -1 1950
box 0 0 6 6
use CELL  118
transform 1 0 1871 0 1 1896
box 0 0 6 6
use CELL  119
transform 1 0 1864 0 1 1896
box 0 0 6 6
use CELL  120
transform 1 0 1765 0 1 1740
box 0 0 6 6
use CELL  121
transform 1 0 1755 0 1 1860
box 0 0 6 6
use CELL  122
transform 1 0 1768 0 1 1824
box 0 0 6 6
use CELL  123
transform 1 0 1790 0 1 1896
box 0 0 6 6
use CELL  124
transform 1 0 1779 0 1 1836
box 0 0 6 6
use CELL  125
transform 1 0 1933 0 1 1812
box 0 0 6 6
use CELL  126
transform -1 0 1945 0 1 1788
box 0 0 6 6
use CELL  127
transform 1 0 1909 0 1 1752
box 0 0 6 6
use CELL  128
transform 1 0 1756 0 1 1740
box 0 0 6 6
use CELL  129
transform -1 0 1977 0 1 1812
box 0 0 6 6
use CELL  130
transform 1 0 1926 0 1 1716
box 0 0 6 6
use CELL  131
transform 1 0 1847 0 -1 1878
box 0 0 6 6
use CELL  132
transform 1 0 1832 0 -1 1758
box 0 0 6 6
use CELL  133
transform 1 0 1867 0 1 1704
box 0 0 6 6
use CELL  134
transform 1 0 1802 0 1 1872
box 0 0 6 6
use CELL  135
transform 1 0 1854 0 1 1788
box 0 0 6 6
use CELL  136
transform 1 0 1785 0 1 1716
box 0 0 6 6
use CELL  137
transform -1 0 1768 0 1 1872
box 0 0 6 6
use CELL  138
transform 1 0 1817 0 1 1884
box 0 0 6 6
use CELL  139
transform 1 0 1756 0 -1 1806
box 0 0 6 6
use CELL  140
transform -1 0 1866 0 1 1776
box 0 0 6 6
use CELL  141
transform 1 0 1866 0 1 1872
box 0 0 6 6
use CELL  142
transform -1 0 1950 0 1 1728
box 0 0 6 6
use CELL  143
transform -1 0 1862 0 -1 1806
box 0 0 6 6
use CELL  144
transform -1 0 1839 0 1 1884
box 0 0 6 6
use CELL  145
transform 1 0 1792 0 1 1716
box 0 0 6 6
use CELL  146
transform -1 0 1761 0 1 1848
box 0 0 6 6
use CELL  147
transform 1 0 1811 0 1 1668
box 0 0 6 6
use CELL  148
transform 1 0 1967 0 1 1800
box 0 0 6 6
use CELL  149
transform 1 0 1870 0 1 1884
box 0 0 6 6
use CELL  150
transform -1 0 1853 0 1 1824
box 0 0 6 6
use CELL  151
transform -1 0 1780 0 1 1752
box 0 0 6 6
use CELL  152
transform -1 0 1829 0 1 1836
box 0 0 6 6
use CELL  153
transform 1 0 1754 0 1 1680
box 0 0 6 6
use CELL  154
transform -1 0 1734 0 1 1740
box 0 0 6 6
use CELL  155
transform -1 0 1966 0 -1 1866
box 0 0 6 6
use CELL  156
transform 1 0 1784 0 1 1680
box 0 0 6 6
use CELL  157
transform -1 0 1915 0 -1 1746
box 0 0 6 6
use CELL  158
transform 1 0 1762 0 1 1932
box 0 0 6 6
use CELL  159
transform 1 0 1940 0 1 1776
box 0 0 6 6
use CELL  160
transform 1 0 1755 0 1 1932
box 0 0 6 6
use CELL  161
transform -1 0 1717 0 -1 1830
box 0 0 6 6
use CELL  162
transform 1 0 1896 0 1 1932
box 0 0 6 6
use CELL  163
transform -1 0 1835 0 1 1824
box 0 0 6 6
use CELL  164
transform 1 0 1828 0 1 1872
box 0 0 6 6
use CELL  165
transform -1 0 1734 0 -1 1662
box 0 0 6 6
use CELL  166
transform -1 0 1815 0 -1 1950
box 0 0 6 6
use CELL  167
transform -1 0 1745 0 1 1764
box 0 0 6 6
use CELL  168
transform 1 0 1794 0 -1 1734
box 0 0 6 6
use CELL  169
transform 1 0 1865 0 1 1848
box 0 0 6 6
use CELL  170
transform -1 0 1955 0 -1 1818
box 0 0 6 6
use CELL  171
transform -1 0 1915 0 1 1884
box 0 0 6 6
use CELL  172
transform 1 0 1963 0 -1 1782
box 0 0 6 6
use CELL  173
transform 1 0 1849 0 1 1848
box 0 0 6 6
use CELL  174
transform 1 0 1814 0 1 1872
box 0 0 6 6
use CELL  175
transform 1 0 1990 0 1 1800
box 0 0 6 6
use CELL  176
transform 1 0 1781 0 1 1872
box 0 0 6 6
use CELL  177
transform -1 0 1984 0 -1 1830
box 0 0 6 6
use CELL  178
transform 1 0 1769 0 1 1860
box 0 0 6 6
use CELL  179
transform 1 0 1780 0 1 1728
box 0 0 6 6
use CELL  180
transform 1 0 1898 0 1 1776
box 0 0 6 6
use CELL  181
transform -1 0 1784 0 1 1800
box 0 0 6 6
use CELL  182
transform 1 0 1859 0 1 1872
box 0 0 6 6
use CELL  183
transform 1 0 1909 0 1 1764
box 0 0 6 6
use CELL  184
transform 1 0 1789 0 1 1884
box 0 0 6 6
use CELL  185
transform 1 0 1764 0 1 1884
box 0 0 6 6
use CELL  186
transform 1 0 1762 0 1 1860
box 0 0 6 6
use CELL  187
transform -1 0 1964 0 1 1824
box 0 0 6 6
use CELL  188
transform -1 0 1743 0 1 1776
box 0 0 6 6
use CELL  189
transform 1 0 1990 0 1 1812
box 0 0 6 6
use CELL  190
transform 1 0 1932 0 -1 1686
box 0 0 6 6
use CELL  191
transform 1 0 1902 0 1 1752
box 0 0 6 6
use CELL  192
transform 1 0 1884 0 1 1860
box 0 0 6 6
use CELL  193
transform 1 0 1865 0 1 1860
box 0 0 6 6
use CELL  194
transform -1 0 1931 0 1 1800
box 0 0 6 6
use CELL  195
transform 1 0 1853 0 1 1860
box 0 0 6 6
use CELL  196
transform 1 0 1745 0 -1 1830
box 0 0 6 6
use CELL  197
transform 1 0 1741 0 1 1872
box 0 0 6 6
use CELL  198
transform 1 0 1932 0 -1 1866
box 0 0 6 6
use CELL  199
transform 1 0 1900 0 1 1884
box 0 0 6 6
use CELL  200
transform -1 0 1913 0 1 1728
box 0 0 6 6
use CELL  201
transform 1 0 1775 0 1 1824
box 0 0 6 6
use CELL  202
transform 1 0 1847 0 1 1788
box 0 0 6 6
use CELL  203
transform -1 0 1827 0 1 1860
box 0 0 6 6
use CELL  204
transform 1 0 1781 0 -1 1854
box 0 0 6 6
use CELL  205
transform 1 0 1862 0 1 1716
box 0 0 6 6
use CELL  206
transform 1 0 1876 0 1 1752
box 0 0 6 6
use CELL  207
transform 1 0 1840 0 1 1788
box 0 0 6 6
use CELL  208
transform 1 0 1846 0 1 1860
box 0 0 6 6
use CELL  209
transform -1 0 1808 0 1 1860
box 0 0 6 6
use CELL  210
transform -1 0 1819 0 1 1764
box 0 0 6 6
use CELL  211
transform -1 0 1737 0 1 1824
box 0 0 6 6
use CELL  212
transform 1 0 1877 0 1 1860
box 0 0 6 6
use CELL  213
transform 1 0 2030 0 -1 1818
box 0 0 6 6
use CELL  214
transform 1 0 1895 0 -1 1806
box 0 0 6 6
use CELL  215
transform 1 0 1796 0 1 1884
box 0 0 6 6
use CELL  216
transform -1 0 1754 0 -1 1770
box 0 0 6 6
use CELL  217
transform 1 0 1853 0 1 1776
box 0 0 6 6
use CELL  218
transform 1 0 1958 0 1 1788
box 0 0 6 6
use CELL  219
transform 1 0 1936 0 1 1704
box 0 0 6 6
use CELL  220
transform 1 0 1932 0 1 1824
box 0 0 6 6
use CELL  221
transform 1 0 1892 0 1 1848
box 0 0 6 6
use CELL  222
transform -1 0 1737 0 1 1680
box 0 0 6 6
use CELL  223
transform 1 0 2004 0 1 1812
box 0 0 6 6
use CELL  224
transform 1 0 1773 0 1 1884
box 0 0 6 6
use CELL  225
transform 1 0 1804 0 -1 1662
box 0 0 6 6
use CELL  226
transform -1 0 1730 0 -1 1830
box 0 0 6 6
use CELL  227
transform 1 0 1828 0 1 1812
box 0 0 6 6
use CELL  228
transform 1 0 1849 0 1 1800
box 0 0 6 6
use CELL  229
transform 1 0 1824 0 1 1728
box 0 0 6 6
use CELL  230
transform -1 0 1957 0 1 1740
box 0 0 6 6
use CELL  231
transform 1 0 1798 0 1 1812
box 0 0 6 6
use CELL  232
transform 1 0 1769 0 1 1848
box 0 0 6 6
use CELL  233
transform -1 0 1717 0 -1 1854
box 0 0 6 6
use CELL  234
transform 1 0 1876 0 1 1812
box 0 0 6 6
use CELL  235
transform 1 0 1899 0 1 1860
box 0 0 6 6
use CELL  236
transform -1 0 1736 0 1 1764
box 0 0 6 6
use CELL  237
transform 1 0 1770 0 1 1764
box 0 0 6 6
use CELL  238
transform -1 0 1888 0 1 1776
box 0 0 6 6
use CELL  239
transform -1 0 1759 0 1 1776
box 0 0 6 6
use CELL  240
transform -1 0 1773 0 1 1752
box 0 0 6 6
use CELL  241
transform 1 0 1923 0 1 1764
box 0 0 6 6
use CELL  242
transform 1 0 1825 0 1 1752
box 0 0 6 6
use CELL  243
transform 1 0 1949 0 1 1776
box 0 0 6 6
use CELL  244
transform 1 0 1843 0 1 1740
box 0 0 6 6
use CELL  245
transform 1 0 1822 0 1 1740
box 0 0 6 6
use CELL  246
transform 1 0 1728 0 -1 1782
box 0 0 6 6
use CELL  247
transform -1 0 1971 0 -1 1794
box 0 0 6 6
use CELL  248
transform 1 0 1848 0 1 1764
box 0 0 6 6
use CELL  249
transform -1 0 1894 0 -1 1746
box 0 0 6 6
use CELL  250
transform 1 0 1905 0 1 1776
box 0 0 6 6
use CELL  251
transform 1 0 1860 0 1 1752
box 0 0 6 6
use CELL  252
transform 1 0 1876 0 1 1836
box 0 0 6 6
use CELL  253
transform -1 0 1978 0 1 1788
box 0 0 6 6
use CELL  254
transform 1 0 1840 0 1 1872
box 0 0 6 6
use CELL  255
transform -1 0 1860 0 1 1824
box 0 0 6 6
use CELL  256
transform 1 0 1829 0 1 1716
box 0 0 6 6
use CELL  257
transform 1 0 1876 0 1 1716
box 0 0 6 6
use CELL  258
transform 1 0 1841 0 1 1764
box 0 0 6 6
use CELL  259
transform 1 0 1900 0 1 1716
box 0 0 6 6
use CELL  260
transform 1 0 1912 0 1 1716
box 0 0 6 6
use CELL  261
transform 1 0 1919 0 1 1716
box 0 0 6 6
use CELL  262
transform 1 0 1801 0 1 1728
box 0 0 6 6
use CELL  263
transform -1 0 1873 0 1 1740
box 0 0 6 6
use CELL  264
transform 1 0 1894 0 1 1704
box 0 0 6 6
use CELL  265
transform -1 0 1798 0 1 1764
box 0 0 6 6
use CELL  266
transform -1 0 1840 0 -1 1662
box 0 0 6 6
use CELL  267
transform -1 0 1845 0 1 1752
box 0 0 6 6
use CELL  268
transform -1 0 1743 0 -1 1794
box 0 0 6 6
use CELL  269
transform 1 0 1738 0 1 1680
box 0 0 6 6
use CELL  270
transform -1 0 1894 0 1 1752
box 0 0 6 6
use CELL  271
transform -1 0 1777 0 1 1728
box 0 0 6 6
use CELL  272
transform 1 0 1770 0 1 1680
box 0 0 6 6
use CELL  273
transform 1 0 1801 0 1 1800
box 0 0 6 6
use CELL  274
transform -1 0 1885 0 -1 1830
box 0 0 6 6
use CELL  275
transform 1 0 1807 0 1 1836
box 0 0 6 6
use CELL  276
transform 1 0 1812 0 1 1680
box 0 0 6 6
use CELL  277
transform -1 0 1743 0 1 1752
box 0 0 6 6
use CELL  278
transform 1 0 1828 0 1 1680
box 0 0 6 6
use CELL  279
transform 1 0 1859 0 1 1680
box 0 0 6 6
use CELL  280
transform 1 0 1878 0 1 1680
box 0 0 6 6
use CELL  281
transform 1 0 1897 0 1 1680
box 0 0 6 6
use CELL  282
transform 1 0 1911 0 1 1680
box 0 0 6 6
use CELL  283
transform 1 0 1925 0 1 1680
box 0 0 6 6
use CELL  284
transform -1 0 1768 0 1 1848
box 0 0 6 6
use CELL  285
transform 1 0 1930 0 -1 1758
box 0 0 6 6
use CELL  286
transform 1 0 1834 0 -1 1770
box 0 0 6 6
use CELL  287
transform 1 0 1826 0 1 1884
box 0 0 6 6
use CELL  288
transform 1 0 1863 0 1 1884
box 0 0 6 6
use CELL  289
transform -1 0 1771 0 1 1836
box 0 0 6 6
use CELL  290
transform -1 0 1768 0 -1 1950
box 0 0 6 6
use CELL  291
transform -1 0 1936 0 1 1740
box 0 0 6 6
use CELL  292
transform 1 0 1820 0 1 1704
box 0 0 6 6
use CELL  293
transform 1 0 1815 0 1 1896
box 0 0 6 6
use CELL  294
transform 1 0 1762 0 1 1704
box 0 0 6 6
use CELL  295
transform 1 0 1778 0 1 1704
box 0 0 6 6
use CELL  296
transform 1 0 1792 0 1 1704
box 0 0 6 6
use CELL  297
transform -1 0 1777 0 1 1716
box 0 0 6 6
use CELL  298
transform 1 0 1781 0 -1 1758
box 0 0 6 6
use CELL  299
transform -1 0 1763 0 1 1884
box 0 0 6 6
use CELL  300
transform -1 0 1840 0 -1 1902
box 0 0 6 6
use CELL  301
transform 1 0 1813 0 1 1716
box 0 0 6 6
use CELL  302
transform 1 0 1923 0 1 1752
box 0 0 6 6
use CELL  303
transform 1 0 1873 0 1 1872
box 0 0 6 6
use CELL  304
transform -1 0 1762 0 1 1812
box 0 0 6 6
use CELL  305
transform 1 0 1880 0 1 1872
box 0 0 6 6
use CELL  306
transform 1 0 1789 0 -1 1950
box 0 0 6 6
use CELL  307
transform 1 0 1951 0 1 1788
box 0 0 6 6
use CELL  308
transform 1 0 1820 0 1 1716
box 0 0 6 6
use CELL  309
transform -1 0 1933 0 -1 1794
box 0 0 6 6
use CELL  310
transform 1 0 1778 0 1 1716
box 0 0 6 6
use CELL  311
transform -1 0 1771 0 1 1776
box 0 0 6 6
use CELL  312
transform -1 0 1900 0 1 1836
box 0 0 6 6
use CELL  313
transform 1 0 1806 0 1 1716
box 0 0 6 6
use CELL  314
transform -1 0 1881 0 -1 1782
box 0 0 6 6
use CELL  315
transform -1 0 1862 0 1 1848
box 0 0 6 6
use CELL  316
transform -1 0 1723 0 -1 1830
box 0 0 6 6
use CELL  317
transform -1 0 1752 0 1 1656
box 0 0 6 6
use CELL  318
transform 1 0 1762 0 1 1716
box 0 0 6 6
use CELL  319
transform 1 0 1723 0 -1 1770
box 0 0 6 6
use CELL  320
transform 1 0 1762 0 1 1728
box 0 0 6 6
use CELL  321
transform 1 0 1742 0 1 1836
box 0 0 6 6
use CELL  322
transform -1 0 1790 0 -1 1818
box 0 0 6 6
use CELL  323
transform 1 0 1781 0 1 1860
box 0 0 6 6
use CELL  324
transform 1 0 1803 0 -1 1746
box 0 0 6 6
use CELL  325
transform 1 0 1977 0 -1 1782
box 0 0 6 6
use CELL  326
transform 1 0 1939 0 1 1824
box 0 0 6 6
use CELL  327
transform 1 0 1806 0 1 1704
box 0 0 6 6
use CELL  328
transform 1 0 1912 0 1 1836
box 0 0 6 6
use CELL  329
transform 1 0 1859 0 -1 1734
box 0 0 6 6
use CELL  330
transform 1 0 1866 0 1 1680
box 0 0 6 6
use CELL  331
transform 1 0 1932 0 1 1764
box 0 0 6 6
use CELL  332
transform 1 0 1783 0 1 1896
box 0 0 6 6
use CELL  333
transform 1 0 1867 0 1 1764
box 0 0 6 6
use CELL  334
transform 1 0 1799 0 1 1896
box 0 0 6 6
use CELL  335
transform 1 0 1827 0 1 1896
box 0 0 6 6
use CELL  336
transform 1 0 1850 0 1 1896
box 0 0 6 6
use CELL  337
transform 1 0 2023 0 -1 1818
box 0 0 6 6
use CELL  338
transform 1 0 1857 0 1 1896
box 0 0 6 6
use CELL  339
transform 1 0 1805 0 1 1680
box 0 0 6 6
use CELL  340
transform 1 0 1852 0 1 1680
box 0 0 6 6
use CELL  341
transform 1 0 1864 0 1 1836
box 0 0 6 6
use CELL  342
transform -1 0 1710 0 1 1824
box 0 0 6 6
use CELL  343
transform 1 0 1958 0 -1 1746
box 0 0 6 6
use CELL  344
transform 1 0 1798 0 -1 1686
box 0 0 6 6
use CELL  345
transform 1 0 1749 0 -1 1806
box 0 0 6 6
use CELL  346
transform 1 0 1880 0 1 1896
box 0 0 6 6
use CELL  347
transform -1 0 1887 0 -1 1770
box 0 0 6 6
use CELL  348
transform 1 0 1820 0 1 1692
box 0 0 6 6
use CELL  349
transform 1 0 1817 0 1 1908
box 0 0 6 6
use CELL  350
transform -1 0 1798 0 -1 1806
box 0 0 6 6
use CELL  351
transform 1 0 1762 0 1 1692
box 0 0 6 6
use CELL  352
transform 1 0 1778 0 1 1692
box 0 0 6 6
use CELL  353
transform 1 0 1806 0 1 1692
box 0 0 6 6
use CELL  354
transform 1 0 1853 0 1 1704
box 0 0 6 6
use CELL  355
transform 1 0 1958 0 -1 1734
box 0 0 6 6
use CELL  356
transform 1 0 1867 0 1 1692
box 0 0 6 6
use CELL  357
transform 1 0 1894 0 1 1692
box 0 0 6 6
use CELL  358
transform 1 0 1908 0 1 1692
box 0 0 6 6
use CELL  359
transform 1 0 1755 0 1 1716
box 0 0 6 6
use CELL  360
transform 1 0 1878 0 1 1788
box 0 0 6 6
use CELL  361
transform -1 0 1930 0 -1 1854
box 0 0 6 6
use CELL  362
transform 1 0 1829 0 1 1740
box 0 0 6 6
use CELL  363
transform 1 0 1939 0 1 1764
box 0 0 6 6
use CELL  364
transform 1 0 1903 0 1 1836
box 0 0 6 6
use CELL  365
transform 1 0 1885 0 1 1788
box 0 0 6 6
use CELL  366
transform -1 0 1966 0 1 1764
box 0 0 6 6
use CELL  367
transform 1 0 1742 0 1 1740
box 0 0 6 6
use CELL  368
transform 1 0 1769 0 1 1908
box 0 0 6 6
use CELL  369
transform 1 0 1783 0 1 1908
box 0 0 6 6
use CELL  370
transform 1 0 1704 0 -1 1782
box 0 0 6 6
use CELL  371
transform 1 0 1836 0 1 1908
box 0 0 6 6
use CELL  372
transform -1 0 1734 0 -1 1842
box 0 0 6 6
use CELL  373
transform 1 0 1782 0 -1 1950
box 0 0 6 6
use CELL  374
transform 1 0 1882 0 1 1908
box 0 0 6 6
use CELL  375
transform 1 0 1811 0 1 1656
box 0 0 6 6
use CELL  376
transform 1 0 1785 0 -1 1770
box 0 0 6 6
use CELL  377
transform 1 0 1819 0 1 1680
box 0 0 6 6
use CELL  378
transform 1 0 1774 0 1 1740
box 0 0 6 6
use CELL  379
transform 1 0 1745 0 1 1680
box 0 0 6 6
use CELL  380
transform 1 0 1740 0 -1 1806
box 0 0 6 6
use CELL  381
transform 1 0 1761 0 1 1680
box 0 0 6 6
use CELL  382
transform 1 0 1777 0 1 1680
box 0 0 6 6
use CELL  383
transform 1 0 1865 0 1 1668
box 0 0 6 6
use CELL  384
transform -1 0 1777 0 -1 1806
box 0 0 6 6
use CELL  385
transform 1 0 1791 0 1 1680
box 0 0 6 6
use CELL  386
transform 1 0 1874 0 -1 1770
box 0 0 6 6
use CELL  387
transform -1 0 1754 0 1 1860
box 0 0 6 6
use CELL  388
transform 1 0 1772 0 -1 1842
box 0 0 6 6
use CELL  389
transform -1 0 1895 0 -1 1782
box 0 0 6 6
use CELL  390
transform 1 0 1808 0 1 1728
box 0 0 6 6
use CELL  391
transform 1 0 1815 0 1 1728
box 0 0 6 6
use CELL  392
transform -1 0 1803 0 1 1776
box 0 0 6 6
use CELL  393
transform 1 0 1831 0 1 1728
box 0 0 6 6
use CELL  394
transform 1 0 1880 0 1 1728
box 0 0 6 6
use CELL  395
transform 1 0 1856 0 -1 1890
box 0 0 6 6
use CELL  396
transform 1 0 1817 0 1 1920
box 0 0 6 6
use CELL  397
transform 1 0 1885 0 1 1680
box 0 0 6 6
use CELL  398
transform -1 0 1766 0 1 1788
box 0 0 6 6
use CELL  399
transform 1 0 1918 0 1 1680
box 0 0 6 6
use CELL  400
transform 1 0 1738 0 1 1692
box 0 0 6 6
use CELL  401
transform -1 0 1913 0 -1 1830
box 0 0 6 6
use CELL  402
transform 1 0 1738 0 1 1704
box 0 0 6 6
use CELL  403
transform 1 0 1853 0 1 1692
box 0 0 6 6
use CELL  404
transform 1 0 1923 0 -1 1866
box 0 0 6 6
use CELL  405
transform -1 0 1946 0 -1 1722
box 0 0 6 6
use CELL  406
transform 1 0 1803 0 1 1884
box 0 0 6 6
use CELL  407
transform 1 0 1738 0 1 1716
box 0 0 6 6
use CELL  408
transform 1 0 1755 0 1 1908
box 0 0 6 6
use CELL  409
transform 1 0 1864 0 1 1812
box 0 0 6 6
use CELL  410
transform -1 0 1754 0 -1 1854
box 0 0 6 6
use CELL  411
transform 1 0 1842 0 1 1884
box 0 0 6 6
use CELL  412
transform -1 0 1852 0 1 1776
box 0 0 6 6
use CELL  413
transform -1 0 1929 0 1 1740
box 0 0 6 6
use CELL  414
transform -1 0 1871 0 1 1800
box 0 0 6 6
use CELL  415
transform 1 0 1792 0 1 1692
box 0 0 6 6
use CELL  416
transform 1 0 1852 0 1 1908
box 0 0 6 6
use CELL  417
transform 1 0 1917 0 1 1848
box 0 0 6 6
use CELL  418
transform 1 0 1849 0 -1 1890
box 0 0 6 6
use CELL  419
transform -1 0 1949 0 1 1704
box 0 0 6 6
use CELL  420
transform -1 0 1922 0 -1 1746
box 0 0 6 6
use CELL  421
transform 1 0 1800 0 1 1836
box 0 0 6 6
use CELL  422
transform -1 0 1710 0 -1 1854
box 0 0 6 6
use CELL  423
transform 1 0 1748 0 1 1884
box 0 0 6 6
use CELL  424
transform 1 0 1748 0 1 1896
box 0 0 6 6
use CELL  425
transform -1 0 1943 0 1 1740
box 0 0 6 6
use CELL  426
transform 1 0 1769 0 -1 1902
box 0 0 6 6
use CELL  427
transform -1 0 1802 0 1 1824
box 0 0 6 6
use CELL  428
transform 1 0 1762 0 1 1908
box 0 0 6 6
use CELL  429
transform 1 0 1748 0 1 1908
box 0 0 6 6
use CELL  430
transform 1 0 1884 0 1 1668
box 0 0 6 6
use CELL  431
transform 1 0 1858 0 1 1668
box 0 0 6 6
use CELL  432
transform -1 0 1851 0 1 1836
box 0 0 6 6
use CELL  433
transform -1 0 1885 0 1 1884
box 0 0 6 6
use CELL  434
transform 1 0 1872 0 1 1668
box 0 0 6 6
use CELL  435
transform 1 0 1939 0 1 1860
box 0 0 6 6
use CELL  436
transform 1 0 1825 0 1 1668
box 0 0 6 6
use CELL  437
transform -1 0 1921 0 1 1788
box 0 0 6 6
use CELL  438
transform 1 0 1811 0 1 1752
box 0 0 6 6
use CELL  439
transform -1 0 1939 0 1 1716
box 0 0 6 6
use CELL  440
transform 1 0 1891 0 1 1824
box 0 0 6 6
use CELL  441
transform 1 0 1788 0 1 1668
box 0 0 6 6
use CELL  442
transform 1 0 1774 0 1 1668
box 0 0 6 6
use CELL  443
transform 1 0 1781 0 1 1668
box 0 0 6 6
use CELL  444
transform 1 0 1828 0 -1 1866
box 0 0 6 6
use CELL  445
transform 1 0 1964 0 1 1812
box 0 0 6 6
use CELL  446
transform 1 0 1793 0 1 1872
box 0 0 6 6
use CELL  447
transform 1 0 1749 0 1 1668
box 0 0 6 6
use CELL  448
transform 1 0 1867 0 1 1752
box 0 0 6 6
use CELL  449
transform 1 0 1734 0 1 1860
box 0 0 6 6
use CELL  450
transform 1 0 1912 0 1 1872
box 0 0 6 6
use CELL  451
transform -1 0 1911 0 -1 1878
box 0 0 6 6
use CELL  452
transform 1 0 1782 0 1 1656
box 0 0 6 6
use CELL  453
transform 1 0 1741 0 1 1896
box 0 0 6 6
use CELL  454
transform -1 0 1820 0 1 1848
box 0 0 6 6
use CELL  455
transform 1 0 1741 0 1 1908
box 0 0 6 6
use CELL  456
transform -1 0 1896 0 -1 1770
box 0 0 6 6
use CELL  457
transform 1 0 1749 0 1 1836
box 0 0 6 6
use CELL  458
transform -1 0 1722 0 -1 1770
box 0 0 6 6
use CELL  459
transform -1 0 1945 0 1 1680
box 0 0 6 6
use CELL  460
transform 1 0 1808 0 1 1908
box 0 0 6 6
use CELL  461
transform -1 0 1734 0 -1 1758
box 0 0 6 6
use CELL  462
transform 1 0 1783 0 1 1920
box 0 0 6 6
use CELL  463
transform 1 0 1801 0 1 1920
box 0 0 6 6
use CELL  464
transform 1 0 1836 0 1 1920
box 0 0 6 6
use CELL  465
transform 1 0 1889 0 1 1908
box 0 0 6 6
use CELL  466
transform -1 0 1750 0 1 1752
box 0 0 6 6
use CELL  467
transform 1 0 1809 0 -1 1866
box 0 0 6 6
use CELL  468
transform 1 0 1751 0 -1 1758
box 0 0 6 6
use CELL  469
transform 1 0 1873 0 1 1908
box 0 0 6 6
use CELL  470
transform -1 0 1925 0 -1 1842
box 0 0 6 6
use CELL  471
transform 1 0 1845 0 1 1908
box 0 0 6 6
use CELL  472
transform -1 0 1816 0 -1 1746
box 0 0 6 6
use CELL  473
transform 1 0 1829 0 1 1908
box 0 0 6 6
use CELL  474
transform -1 0 1754 0 1 1872
box 0 0 6 6
use CELL  475
transform 1 0 1829 0 1 1704
box 0 0 6 6
use CELL  476
transform -1 0 1932 0 1 1836
box 0 0 6 6
use CELL  477
transform 1 0 1923 0 -1 1734
box 0 0 6 6
use CELL  478
transform 1 0 1763 0 1 1812
box 0 0 6 6
use CELL  479
transform 1 0 1776 0 1 1788
box 0 0 6 6
use CELL  480
transform 1 0 1769 0 1 1872
box 0 0 6 6
use CELL  481
transform 1 0 1983 0 1 1812
box 0 0 6 6
use CELL  482
transform -1 0 1759 0 1 1788
box 0 0 6 6
use CELL  483
transform -1 0 1908 0 1 1764
box 0 0 6 6
use CELL  484
transform 1 0 1931 0 1 1848
box 0 0 6 6
use CELL  485
transform 1 0 1785 0 1 1800
box 0 0 6 6
use CELL  486
transform 1 0 1813 0 1 1704
box 0 0 6 6
use CELL  487
transform 1 0 1915 0 1 1704
box 0 0 6 6
use CELL  488
transform 1 0 1843 0 1 1896
box 0 0 6 6
use CELL  489
transform 1 0 1716 0 1 1860
box 0 0 6 6
use CELL  490
transform 1 0 1860 0 1 1692
box 0 0 6 6
use CELL  491
transform 1 0 1802 0 1 1944
box 0 0 6 6
use CELL  492
transform 1 0 1755 0 1 1704
box 0 0 6 6
use CELL  493
transform -1 0 1758 0 -1 1830
box 0 0 6 6
use CELL  494
transform 1 0 1776 0 1 1896
box 0 0 6 6
use CELL  495
transform 1 0 1833 0 1 1848
box 0 0 6 6
use CELL  496
transform 1 0 1734 0 1 1932
box 0 0 6 6
use CELL  497
transform 1 0 1741 0 1 1932
box 0 0 6 6
use CELL  498
transform -1 0 1880 0 1 1848
box 0 0 6 6
use CELL  499
transform 1 0 1748 0 1 1932
box 0 0 6 6
use CELL  500
transform -1 0 1942 0 1 1752
box 0 0 6 6
use CELL  501
transform -1 0 1803 0 1 1656
box 0 0 6 6
use CELL  502
transform 1 0 1889 0 1 1920
box 0 0 6 6
use CELL  503
transform 1 0 1873 0 1 1920
box 0 0 6 6
use CELL  504
transform 1 0 1859 0 1 1920
box 0 0 6 6
use CELL  505
transform -1 0 1761 0 -1 1770
box 0 0 6 6
use CELL  506
transform -1 0 1889 0 1 1848
box 0 0 6 6
use CELL  507
transform -1 0 1844 0 1 1836
box 0 0 6 6
use CELL  508
transform 1 0 1873 0 1 1932
box 0 0 6 6
use CELL  509
transform 1 0 1734 0 -1 1854
box 0 0 6 6
use CELL  510
transform 1 0 1776 0 1 1920
box 0 0 6 6
use CELL  511
transform 1 0 1755 0 1 1944
box 0 0 6 6
use CELL  512
transform -1 0 1892 0 1 1884
box 0 0 6 6
use CELL  513
transform 1 0 1799 0 1 1716
box 0 0 6 6
use CELL  514
transform -1 0 1747 0 1 1860
box 0 0 6 6
use CELL  515
transform -1 0 1744 0 1 1728
box 0 0 6 6
use CELL  516
transform 1 0 1748 0 1 1920
box 0 0 6 6
use CELL  517
transform 1 0 1734 0 1 1920
box 0 0 6 6
use CELL  518
transform 1 0 1903 0 1 1932
box 0 0 6 6
use CELL  519
transform 1 0 1728 0 1 1800
box 0 0 6 6
use CELL  520
transform 1 0 1997 0 1 1800
box 0 0 6 6
use CELL  521
transform 1 0 1889 0 1 1932
box 0 0 6 6
use CELL  522
transform 1 0 1882 0 1 1932
box 0 0 6 6
use CELL  523
transform -1 0 1861 0 1 1764
box 0 0 6 6
use CELL  524
transform 1 0 1808 0 1 1920
box 0 0 6 6
use CELL  525
transform 1 0 1769 0 1 1932
box 0 0 6 6
use CELL  526
transform 1 0 1776 0 1 1932
box 0 0 6 6
use CELL  527
transform 1 0 1783 0 1 1932
box 0 0 6 6
use CELL  528
transform -1 0 1960 0 1 1716
box 0 0 6 6
use CELL  529
transform 1 0 1802 0 1 1848
box 0 0 6 6
use CELL  530
transform 1 0 1917 0 1 1668
box 0 0 6 6
use CELL  531
transform 1 0 1916 0 1 1764
box 0 0 6 6
use CELL  532
transform 1 0 1924 0 1 1668
box 0 0 6 6
use CELL  533
transform 1 0 1937 0 -1 1734
box 0 0 6 6
use CELL  534
transform 1 0 1953 0 1 1764
box 0 0 6 6
use CELL  535
transform 1 0 1758 0 1 1836
box 0 0 6 6
use CELL  536
transform 1 0 1903 0 1 1908
box 0 0 6 6
use CELL  537
transform 1 0 1746 0 -1 1650
box 0 0 6 6
use CELL  538
transform 1 0 1988 0 1 1788
box 0 0 6 6
use CELL  539
transform -1 0 2001 0 1 1788
box 0 0 6 6
use CELL  540
transform 1 0 1965 0 1 1824
box 0 0 6 6
use CELL  541
transform 1 0 1734 0 1 1884
box 0 0 6 6
use CELL  542
transform 1 0 1944 0 1 1740
box 0 0 6 6
use CELL  543
transform 1 0 1919 0 1 1872
box 0 0 6 6
use CELL  544
transform 1 0 1997 0 1 1812
box 0 0 6 6
use CELL  545
transform 1 0 1734 0 1 1896
box 0 0 6 6
use CELL  546
transform 1 0 1901 0 1 1896
box 0 0 6 6
use CELL  547
transform 1 0 1734 0 1 1908
box 0 0 6 6
use CELL  548
transform 1 0 1731 0 1 1692
box 0 0 6 6
use CELL  549
transform -1 0 1936 0 1 1728
box 0 0 6 6
use CELL  550
transform 1 0 1755 0 1 1692
box 0 0 6 6
use CELL  551
transform 1 0 1771 0 1 1692
box 0 0 6 6
use CELL  552
transform 1 0 1785 0 1 1692
box 0 0 6 6
use CELL  553
transform -1 0 1740 0 -1 1950
box 0 0 6 6
use CELL  554
transform -1 0 1812 0 1 1896
box 0 0 6 6
use CELL  555
transform -1 0 1752 0 1 1788
box 0 0 6 6
use CELL  556
transform -1 0 1901 0 1 1752
box 0 0 6 6
use CELL  557
transform 1 0 1762 0 -1 1902
box 0 0 6 6
use CELL  558
transform 1 0 1829 0 1 1692
box 0 0 6 6
use CELL  559
transform 1 0 1755 0 1 1896
box 0 0 6 6
use CELL  560
transform -1 0 1795 0 1 1740
box 0 0 6 6
use CELL  561
transform 1 0 1882 0 1 1692
box 0 0 6 6
use CELL  562
transform 1 0 1901 0 1 1692
box 0 0 6 6
use CELL  563
transform -1 0 1891 0 -1 1842
box 0 0 6 6
use CELL  564
transform 1 0 1810 0 1 1884
box 0 0 6 6
use CELL  565
transform 1 0 1882 0 1 1920
box 0 0 6 6
use CELL  566
transform 1 0 1896 0 1 1920
box 0 0 6 6
use CELL  567
transform 1 0 1818 0 1 1668
box 0 0 6 6
use CELL  568
transform 1 0 1817 0 1 1932
box 0 0 6 6
use CELL  569
transform 1 0 1735 0 1 1668
box 0 0 6 6
use CELL  570
transform 1 0 1742 0 1 1668
box 0 0 6 6
use CELL  571
transform 1 0 1785 0 1 1704
box 0 0 6 6
use CELL  572
transform 1 0 1981 0 1 1788
box 0 0 6 6
use CELL  573
transform -1 0 1778 0 1 1776
box 0 0 6 6
use CELL  574
transform 1 0 1915 0 1 1692
box 0 0 6 6
use CELL  575
transform 1 0 1741 0 1 1920
box 0 0 6 6
use CELL  576
transform 1 0 1946 0 1 1860
box 0 0 6 6
use CELL  577
transform 1 0 1942 0 1 1836
box 0 0 6 6
use CELL  578
transform -1 0 1761 0 1 1728
box 0 0 6 6
use CELL  579
transform -1 0 1755 0 1 1812
box 0 0 6 6
use CELL  580
transform 1 0 1808 0 1 1932
box 0 0 6 6
use CELL  581
transform 1 0 1829 0 1 1932
box 0 0 6 6
use CELL  582
transform 1 0 1852 0 1 1932
box 0 0 6 6
use CELL  583
transform 1 0 1859 0 1 1932
box 0 0 6 6
use CELL  584
transform 1 0 1866 0 1 1932
box 0 0 6 6
use CELL  585
transform 1 0 1845 0 1 1932
box 0 0 6 6
use CELL  586
transform 1 0 1735 0 1 1836
box 0 0 6 6
use CELL  587
transform 1 0 1767 0 1 1668
box 0 0 6 6
use CELL  588
transform 1 0 1910 0 1 1848
box 0 0 6 6
use CELL  589
transform 1 0 1731 0 1 1728
box 0 0 6 6
use CELL  590
transform 1 0 1838 0 1 1728
box 0 0 6 6
use CELL  591
transform -1 0 1847 0 -1 1662
box 0 0 6 6
use CELL  592
transform 1 0 1731 0 1 1716
box 0 0 6 6
use CELL  593
transform -1 0 1902 0 1 1872
box 0 0 6 6
use CELL  594
transform -1 0 1966 0 1 1800
box 0 0 6 6
use CELL  595
transform -1 0 1904 0 -1 1830
box 0 0 6 6
use CELL  596
transform 1 0 1929 0 1 1692
box 0 0 6 6
use CELL  597
transform 1 0 1825 0 -1 1794
box 0 0 6 6
use CELL  598
transform 1 0 1903 0 1 1668
box 0 0 6 6
use CELL  599
transform 1 0 1891 0 1 1668
box 0 0 6 6
use CELL  600
transform 1 0 1796 0 1 1740
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 1871 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 1832 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 1826 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 1746 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 1746 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 1743 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 1743 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 1745 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 1842 0 1 1932
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 1842 0 1 1920
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 1842 0 1 1908
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 1840 0 1 1896
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 1839 0 1 1884
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 1856 0 1 1872
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 1859 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 1788 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 1767 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 1764 0 1 1752
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 1762 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 1768 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 1768 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 1768 0 1 1704
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 1768 0 1 1692
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 1767 0 1 1680
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 1764 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 1759 0 1 1656
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 1887 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 1873 0 1 1752
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 1873 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 1952 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 2010 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 1980 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 1978 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 1946 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 1929 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 1728 0 1 1680
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 1728 0 1 1692
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 1728 0 1 1704
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 1728 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 1728 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 1890 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 1889 0 1 1848
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 1891 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 1913 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 1977 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 1947 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 1945 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 1911 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 1899 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 1882 0 1 1752
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 1885 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 1877 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 1888 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 1879 0 1 1704
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 1879 0 1 1692
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 1802 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 1794 0 1 1656
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 1933 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 1938 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 1835 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 1835 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 1888 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 1862 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 1860 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 1840 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 1837 0 1 1872
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 1823 0 1 1884
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 1821 0 1 1896
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 1823 0 1 1908
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 1823 0 1 1920
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 1823 0 1 1932
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 1900 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 1901 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 1906 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 1888 0 1 1704
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 1888 0 1 1692
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 1891 0 1 1680
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 1897 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 1771 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 1831 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 1825 0 1 1680
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 1826 0 1 1692
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 1826 0 1 1704
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 1826 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 1755 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 1751 0 1 1680
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 1752 0 1 1692
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 1752 0 1 1704
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 1752 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 1752 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 1961 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 1885 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 1873 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 1880 0 1 1848
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 1874 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 1936 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 1909 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 1920 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 1859 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 1850 0 1 1704
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 1850 0 1 1692
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 1849 0 1 1680
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 1855 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 1810 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 1798 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 1795 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 1791 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 1798 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-109
transform 1 0 1793 0 1 1752
box 0 0 3 6
use FEEDTHRU  F-110
transform 1 0 1786 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-111
transform 1 0 1777 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-112
transform 1 0 1813 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-113
transform 1 0 1787 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-114
transform 1 0 1797 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-115
transform 1 0 1799 0 1 1848
box 0 0 3 6
use FEEDTHRU  F-116
transform 1 0 1799 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-117
transform 1 0 1799 0 1 1872
box 0 0 3 6
use FEEDTHRU  F-118
transform 1 0 1734 0 1 1752
box 0 0 3 6
use FEEDTHRU  F-119
transform 1 0 1736 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-120
transform 1 0 1734 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-121
transform 1 0 1734 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-122
transform 1 0 1768 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-123
transform 1 0 1778 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-124
transform 1 0 1754 0 1 1884
box 0 0 3 6
use FEEDTHRU  F-125
transform 1 0 1891 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-126
transform 1 0 1824 0 1 1656
box 0 0 3 6
use FEEDTHRU  F-127
transform 1 0 1814 0 1 1932
box 0 0 3 6
use FEEDTHRU  F-128
transform 1 0 1814 0 1 1920
box 0 0 3 6
use FEEDTHRU  F-129
transform 1 0 1814 0 1 1908
box 0 0 3 6
use FEEDTHRU  F-130
transform 1 0 1812 0 1 1896
box 0 0 3 6
use FEEDTHRU  F-131
transform 1 0 1948 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-132
transform 1 0 1950 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-133
transform 1 0 1980 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-134
transform 1 0 1811 0 1 1848
box 0 0 3 6
use FEEDTHRU  F-135
transform 1 0 1818 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-136
transform 1 0 1811 0 1 1872
box 0 0 3 6
use FEEDTHRU  F-137
transform 1 0 1770 0 1 1884
box 0 0 3 6
use FEEDTHRU  F-138
transform 1 0 1838 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-139
transform 1 0 1904 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-140
transform 1 0 1831 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-141
transform 1 0 1830 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-142
transform 1 0 1831 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-143
transform 1 0 1828 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-144
transform 1 0 1819 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-145
transform 1 0 1827 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-146
transform 1 0 1828 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-147
transform 1 0 1808 0 1 1752
box 0 0 3 6
use FEEDTHRU  F-148
transform 1 0 1824 0 1 1896
box 0 0 3 6
use FEEDTHRU  F-149
transform 1 0 1826 0 1 1908
box 0 0 3 6
use FEEDTHRU  F-150
transform 1 0 1826 0 1 1920
box 0 0 3 6
use FEEDTHRU  F-151
transform 1 0 1826 0 1 1932
box 0 0 3 6
use FEEDTHRU  F-152
transform 1 0 1805 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-153
transform 1 0 1822 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-154
transform 1 0 1819 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-155
transform 1 0 1816 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-156
transform 1 0 1824 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-157
transform 1 0 1868 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-158
transform 1 0 1894 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-159
transform 1 0 1913 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-160
transform 1 0 1930 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-161
transform 1 0 1825 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-162
transform 1 0 1822 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-163
transform 1 0 1822 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-164
transform 1 0 1821 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-165
transform 1 0 1819 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-166
transform 1 0 1819 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-167
transform 1 0 1805 0 1 1752
box 0 0 3 6
use FEEDTHRU  F-168
transform 1 0 1825 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-169
transform 1 0 1836 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-170
transform 1 0 1837 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-171
transform 1 0 1846 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-172
transform 1 0 1861 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-173
transform 1 0 1790 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-174
transform 1 0 1791 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-175
transform 1 0 1830 0 1 1848
box 0 0 3 6
use FEEDTHRU  F-176
transform 1 0 1837 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-177
transform 1 0 1790 0 1 1872
box 0 0 3 6
use FEEDTHRU  F-178
transform 1 0 1779 0 1 1884
box 0 0 3 6
use FEEDTHRU  F-179
transform 1 0 1796 0 1 1896
box 0 0 3 6
use FEEDTHRU  F-180
transform 1 0 1798 0 1 1908
box 0 0 3 6
use FEEDTHRU  F-181
transform 1 0 1798 0 1 1920
box 0 0 3 6
use FEEDTHRU  F-182
transform 1 0 1798 0 1 1932
box 0 0 3 6
use FEEDTHRU  F-183
transform 1 0 1932 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-184
transform 1 0 1937 0 1 1848
box 0 0 3 6
use FEEDTHRU  F-185
transform 1 0 1929 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-186
transform 1 0 1925 0 1 1872
box 0 0 3 6
use FEEDTHRU  F-187
transform 1 0 1906 0 1 1884
box 0 0 3 6
use FEEDTHRU  F-188
transform 1 0 1792 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-189
transform 1 0 1785 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-190
transform 1 0 1900 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-191
transform 1 0 1907 0 1 1848
box 0 0 3 6
use FEEDTHRU  F-192
transform 1 0 1908 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-193
transform 1 0 1893 0 1 1872
box 0 0 3 6
use FEEDTHRU  F-194
transform 1 0 1876 0 1 1884
box 0 0 3 6
use FEEDTHRU  F-195
transform 1 0 1877 0 1 1896
box 0 0 3 6
use FEEDTHRU  F-196
transform 1 0 1879 0 1 1908
box 0 0 3 6
use FEEDTHRU  F-197
transform 1 0 1879 0 1 1920
box 0 0 3 6
use FEEDTHRU  F-198
transform 1 0 1879 0 1 1932
box 0 0 3 6
use FEEDTHRU  F-199
transform 1 0 1903 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-200
transform 1 0 1866 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-201
transform 1 0 1858 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-202
transform 1 0 1902 0 1 1872
box 0 0 3 6
use FEEDTHRU  F-203
transform 1 0 1911 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-204
transform 1 0 1844 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-205
transform 1 0 1847 0 1 1704
box 0 0 3 6
use FEEDTHRU  F-206
transform 1 0 1847 0 1 1692
box 0 0 3 6
use FEEDTHRU  F-207
transform 1 0 1846 0 1 1680
box 0 0 3 6
use FEEDTHRU  F-208
transform 1 0 1852 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-209
transform 1 0 1876 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-210
transform 1 0 1769 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-211
transform 1 0 1765 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-212
transform 1 0 1775 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-213
transform 1 0 1922 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-214
transform 1 0 1870 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-215
transform 1 0 1813 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-216
transform 1 0 1810 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-217
transform 1 0 1809 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-218
transform 1 0 1807 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-219
transform 1 0 1913 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-220
transform 1 0 1789 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-221
transform 1 0 1776 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-222
transform 1 0 1912 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-223
transform 1 0 1782 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-224
transform 1 0 1850 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-225
transform 1 0 1841 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-226
transform 1 0 1844 0 1 1704
box 0 0 3 6
use FEEDTHRU  F-227
transform 1 0 1844 0 1 1692
box 0 0 3 6
use FEEDTHRU  F-228
transform 1 0 1843 0 1 1680
box 0 0 3 6
use FEEDTHRU  F-229
transform 1 0 1849 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-230
transform 1 0 1856 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-231
transform 1 0 1865 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-232
transform 1 0 1846 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-233
transform 1 0 1840 0 1 1680
box 0 0 3 6
use FEEDTHRU  F-234
transform 1 0 1841 0 1 1692
box 0 0 3 6
use FEEDTHRU  F-235
transform 1 0 1841 0 1 1704
box 0 0 3 6
use FEEDTHRU  F-236
transform 1 0 1847 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-237
transform 1 0 1874 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-238
transform 1 0 1849 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-239
transform 1 0 1857 0 1 1752
box 0 0 3 6
use FEEDTHRU  F-240
transform 1 0 1864 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-241
transform 1 0 1872 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-242
transform 1 0 1875 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-243
transform 1 0 1886 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-244
transform 1 0 1906 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-245
transform 1 0 1869 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-246
transform 1 0 1870 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-247
transform 1 0 1871 0 1 1848
box 0 0 3 6
use FEEDTHRU  F-248
transform 1 0 1871 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-249
transform 1 0 1861 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-250
transform 1 0 1906 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-251
transform 1 0 1789 0 1 1932
box 0 0 3 6
use FEEDTHRU  F-252
transform 1 0 1789 0 1 1920
box 0 0 3 6
use FEEDTHRU  F-253
transform 1 0 1789 0 1 1908
box 0 0 3 6
use FEEDTHRU  F-254
transform 1 0 1895 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-255
transform 1 0 1909 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-256
transform 1 0 1787 0 1 1872
box 0 0 3 6
use FEEDTHRU  F-257
transform 1 0 1858 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-258
transform 1 0 1854 0 1 1752
box 0 0 3 6
use FEEDTHRU  F-259
transform 1 0 1861 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-260
transform 1 0 1869 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-261
transform 1 0 1872 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-262
transform 1 0 1883 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-263
transform 1 0 1900 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-264
transform 1 0 1863 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-265
transform 1 0 1808 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-266
transform 1 0 1866 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-267
transform 1 0 1869 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-268
transform 1 0 1871 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-269
transform 1 0 1912 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-270
transform 1 0 1860 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-271
transform 1 0 1861 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-272
transform 1 0 1862 0 1 1848
box 0 0 3 6
use FEEDTHRU  F-273
transform 1 0 1862 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-274
transform 1 0 1853 0 1 1872
box 0 0 3 6
use FEEDTHRU  F-275
transform 1 0 1843 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-276
transform 1 0 1814 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-277
transform 1 0 1820 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-278
transform 1 0 1808 0 1 1848
box 0 0 3 6
use FEEDTHRU  F-279
transform 1 0 1815 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-280
transform 1 0 1808 0 1 1872
box 0 0 3 6
use FEEDTHRU  F-281
transform 1 0 1930 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-282
transform 1 0 1773 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-283
transform 1 0 1762 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-284
transform 1 0 1781 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-285
transform 1 0 1758 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-286
transform 1 0 1755 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-287
transform 1 0 1834 0 1 1872
box 0 0 3 6
use FEEDTHRU  F-288
transform 1 0 1843 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-289
transform 1 0 1839 0 1 1848
box 0 0 3 6
use FEEDTHRU  F-290
transform 1 0 1904 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-291
transform 1 0 1897 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-292
transform 1 0 1852 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-293
transform 1 0 1831 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-294
transform 1 0 1834 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-295
transform 1 0 1833 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-296
transform 1 0 1822 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-297
transform 1 0 1802 0 1 1752
box 0 0 3 6
use FEEDTHRU  F-298
transform 1 0 1816 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-299
transform 1 0 1821 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-300
transform 1 0 1880 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-301
transform 1 0 1834 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-302
transform 1 0 1827 0 1 1848
box 0 0 3 6
use FEEDTHRU  F-303
transform 1 0 1829 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-304
transform 1 0 1823 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-305
transform 1 0 1858 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-306
transform 1 0 1843 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-307
transform 1 0 1851 0 1 1752
box 0 0 3 6
use FEEDTHRU  F-308
transform 1 0 1779 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-309
transform 1 0 1794 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-310
transform 1 0 1904 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-311
transform 1 0 1939 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-312
transform 1 0 1922 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-313
transform 1 0 1909 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-314
transform 1 0 1914 0 1 1776
box 0 0 3 6
use FEEDTHRU  F-315
transform 1 0 1896 0 1 1764
box 0 0 3 6
use FEEDTHRU  F-316
transform 1 0 1885 0 1 1752
box 0 0 3 6
use FEEDTHRU  F-317
transform 1 0 1903 0 1 1740
box 0 0 3 6
use FEEDTHRU  F-318
transform 1 0 1898 0 1 1728
box 0 0 3 6
use FEEDTHRU  F-319
transform 1 0 1891 0 1 1716
box 0 0 3 6
use FEEDTHRU  F-320
transform 1 0 1891 0 1 1704
box 0 0 3 6
use FEEDTHRU  F-321
transform 1 0 1891 0 1 1692
box 0 0 3 6
use FEEDTHRU  F-322
transform 1 0 1894 0 1 1680
box 0 0 3 6
use FEEDTHRU  F-323
transform 1 0 1900 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-324
transform 1 0 1904 0 1 1848
box 0 0 3 6
use FEEDTHRU  F-325
transform 1 0 1905 0 1 1860
box 0 0 3 6
use FEEDTHRU  F-326
transform 1 0 1825 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-327
transform 1 0 1840 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-328
transform 1 0 1909 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-329
transform 1 0 1955 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-330
transform 1 0 2013 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-331
transform 1 0 1882 0 1 1836
box 0 0 3 6
use FEEDTHRU  F-332
transform 1 0 1888 0 1 1824
box 0 0 3 6
use FEEDTHRU  F-333
transform 1 0 1927 0 1 1812
box 0 0 3 6
use FEEDTHRU  F-334
transform 1 0 1901 0 1 1800
box 0 0 3 6
use FEEDTHRU  F-335
transform 1 0 1891 0 1 1788
box 0 0 3 6
use FEEDTHRU  F-336
transform 1 0 1895 0 1 1776
box 0 0 3 6
<< end >>
