magic
tech scmos
timestamp 1394680307
<< m1p >>
use CELL  1
transform 1 0 291 0 1 264
box 0 0 6 6
use CELL  2
transform -1 0 249 0 1 276
box 0 0 6 6
use CELL  3
transform -1 0 310 0 -1 282
box 0 0 6 6
use CELL  4
transform -1 0 269 0 1 252
box 0 0 6 6
use CELL  5
transform -1 0 318 0 1 264
box 0 0 6 6
use CELL  6
transform 1 0 279 0 -1 294
box 0 0 6 6
use CELL  7
transform -1 0 257 0 1 264
box 0 0 6 6
use CELL  8
transform -1 0 277 0 1 276
box 0 0 6 6
use CELL  9
transform 1 0 271 0 -1 318
box 0 0 6 6
use CELL  10
transform -1 0 294 0 -1 258
box 0 0 6 6
use CELL  11
transform -1 0 262 0 1 288
box 0 0 6 6
use CELL  12
transform 1 0 256 0 -1 222
box 0 0 6 6
use CELL  13
transform -1 0 234 0 -1 258
box 0 0 6 6
use CELL  14
transform -1 0 252 0 1 240
box 0 0 6 6
use CELL  15
transform 1 0 273 0 1 300
box 0 0 6 6
use CELL  16
transform -1 0 260 0 1 204
box 0 0 6 6
use CELL  17
transform -1 0 246 0 1 216
box 0 0 6 6
use CELL  18
transform 1 0 252 0 1 300
box 0 0 6 6
use CELL  19
transform 1 0 259 0 1 300
box 0 0 6 6
use CELL  20
transform -1 0 246 0 -1 210
box 0 0 6 6
use CELL  21
transform -1 0 293 0 -1 306
box 0 0 6 6
use CELL  22
transform -1 0 299 0 -1 294
box 0 0 6 6
use CELL  23
transform 1 0 272 0 1 216
box 0 0 6 6
use CELL  24
transform -1 0 276 0 1 288
box 0 0 6 6
use CELL  25
transform -1 0 285 0 1 216
box 0 0 6 6
use CELL  26
transform -1 0 266 0 1 240
box 0 0 6 6
use CELL  27
transform -1 0 312 0 1 228
box 0 0 6 6
use CELL  28
transform -1 0 311 0 1 264
box 0 0 6 6
use CELL  29
transform -1 0 292 0 1 216
box 0 0 6 6
use CELL  30
transform -1 0 271 0 1 216
box 0 0 6 6
use CELL  31
transform -1 0 306 0 1 288
box 0 0 6 6
use CELL  32
transform 1 0 266 0 1 300
box 0 0 6 6
use CELL  33
transform -1 0 246 0 1 252
box 0 0 6 6
use CELL  34
transform -1 0 240 0 1 228
box 0 0 6 6
use CELL  35
transform 1 0 240 0 -1 294
box 0 0 6 6
use CELL  36
transform -1 0 240 0 1 276
box 0 0 6 6
use CELL  37
transform -1 0 285 0 1 252
box 0 0 6 6
use CELL  38
transform -1 0 301 0 1 240
box 0 0 6 6
use CELL  39
transform -1 0 308 0 1 240
box 0 0 6 6
use CELL  40
transform -1 0 291 0 1 228
box 0 0 6 6
use CELL  41
transform 1 0 261 0 1 204
box 0 0 6 6
use CELL  42
transform -1 0 305 0 1 228
box 0 0 6 6
use CELL  43
transform -1 0 286 0 1 300
box 0 0 6 6
use CELL  44
transform -1 0 241 0 1 264
box 0 0 6 6
use CELL  45
transform -1 0 345 0 1 276
box 0 0 6 6
use CELL  46
transform -1 0 262 0 1 252
box 0 0 6 6
use CELL  47
transform 1 0 272 0 -1 270
box 0 0 6 6
use CELL  48
transform 1 0 295 0 -1 258
box 0 0 6 6
use CELL  49
transform -1 0 259 0 1 240
box 0 0 6 6
use CELL  50
transform 1 0 313 0 1 228
box 0 0 6 6
use CELL  51
transform 1 0 247 0 -1 210
box 0 0 6 6
use CELL  52
transform -1 0 250 0 1 264
box 0 0 6 6
use CELL  53
transform -1 0 278 0 1 252
box 0 0 6 6
use CELL  54
transform -1 0 317 0 1 240
box 0 0 6 6
use CELL  55
transform 1 0 265 0 1 312
box 0 0 6 6
use CELL  56
transform -1 0 234 0 1 264
box 0 0 6 6
use CELL  57
transform 1 0 278 0 1 276
box 0 0 6 6
use CELL  58
transform -1 0 256 0 1 276
box 0 0 6 6
use CELL  59
transform -1 0 308 0 1 252
box 0 0 6 6
use CELL  60
transform -1 0 324 0 1 240
box 0 0 6 6
use CELL  61
transform -1 0 247 0 1 228
box 0 0 6 6
use CELL  62
transform -1 0 324 0 1 276
box 0 0 6 6
use CELL  63
transform 1 0 258 0 1 312
box 0 0 6 6
use CELL  64
transform 1 0 250 0 -1 234
box 0 0 6 6
use CELL  65
transform -1 0 253 0 1 216
box 0 0 6 6
use CELL  66
transform 1 0 279 0 1 264
box 0 0 6 6
use CELL  67
transform 1 0 297 0 1 276
box 0 0 6 6
use CELL  68
transform -1 0 269 0 1 288
box 0 0 6 6
use CELL  69
transform -1 0 331 0 1 240
box 0 0 6 6
use CELL  70
transform -1 0 255 0 -1 294
box 0 0 6 6
use CELL  71
transform 1 0 307 0 1 288
box 0 0 6 6
use CELL  72
transform -1 0 255 0 -1 258
box 0 0 6 6
use CELL  73
transform -1 0 331 0 1 276
box 0 0 6 6
use CELL  74
transform -1 0 268 0 1 228
box 0 0 6 6
use CELL  75
transform -1 0 317 0 1 276
box 0 0 6 6
use CELL  76
transform -1 0 268 0 1 276
box 0 0 6 6
use CELL  77
transform -1 0 273 0 1 240
box 0 0 6 6
use CELL  78
transform -1 0 284 0 1 228
box 0 0 6 6
use CELL  79
transform -1 0 274 0 1 204
box 0 0 6 6
use CELL  80
transform -1 0 281 0 1 204
box 0 0 6 6
use CELL  81
transform -1 0 294 0 -1 246
box 0 0 6 6
use CELL  82
transform -1 0 275 0 1 228
box 0 0 6 6
use CELL  83
transform -1 0 296 0 1 276
box 0 0 6 6
use CELL  84
transform -1 0 269 0 1 264
box 0 0 6 6
use CELL  85
transform -1 0 292 0 1 288
box 0 0 6 6
use CELL  86
transform -1 0 322 0 1 252
box 0 0 6 6
use CELL  87
transform -1 0 315 0 1 252
box 0 0 6 6
use CELL  88
transform 1 0 332 0 -1 282
box 0 0 6 6
use CELL  89
transform -1 0 304 0 1 264
box 0 0 6 6
use CELL  90
transform -1 0 298 0 1 228
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 285 0 1 264
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 284 0 1 276
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 276 0 1 288
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 256 0 1 276
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 257 0 1 264
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 234 0 1 252
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 253 0 1 216
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 256 0 1 228
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 247 0 1 228
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 246 0 1 252
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 287 0 1 276
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 275 0 1 228
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 308 0 1 240
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 240 0 1 240
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 243 0 1 240
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 269 0 1 264
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 268 0 1 276
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 259 0 1 228
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 262 0 1 216
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 279 0 1 240
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 269 0 1 252
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 282 0 1 240
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 285 0 1 240
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 237 0 1 252
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 241 0 1 264
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 240 0 1 276
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 246 0 1 288
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 240 0 1 300
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 260 0 1 264
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 259 0 1 276
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 285 0 1 252
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 288 0 1 264
box 0 0 3 6
<< end >>
