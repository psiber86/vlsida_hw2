magic
tech scmos
timestamp 1395743065
<< m1p >>
use CELL  1
transform 1 0 102 0 1 46
box 0 0 6 6
use CELL  2
transform -1 0 179 0 1 120
box 0 0 6 6
use CELL  3
transform 1 0 167 0 1 196
box 0 0 6 6
use CELL  4
transform 1 0 90 0 -1 227
box 0 0 6 6
use CELL  5
transform -1 0 112 0 1 221
box 0 0 6 6
use CELL  6
transform -1 0 146 0 -1 68
box 0 0 6 6
use CELL  7
transform -1 0 96 0 1 196
box 0 0 6 6
use CELL  8
transform -1 0 102 0 1 62
box 0 0 6 6
use CELL  9
transform -1 0 186 0 1 120
box 0 0 6 6
use CELL  10
transform 1 0 201 0 1 161
box 0 0 6 6
use CELL  11
transform -1 0 170 0 1 120
box 0 0 6 6
use CELL  12
transform 1 0 176 0 1 196
box 0 0 6 6
use CELL  13
transform -1 0 90 0 1 161
box 0 0 6 6
use CELL  14
transform -1 0 171 0 1 161
box 0 0 6 6
use CELL  15
transform -1 0 155 0 1 196
box 0 0 6 6
use CELL  16
transform -1 0 139 0 1 62
box 0 0 6 6
use CELL  17
transform 1 0 183 0 1 196
box 0 0 6 6
use CELL  18
transform -1 0 105 0 1 221
box 0 0 6 6
use CELL  19
transform 1 0 160 0 1 221
box 0 0 6 6
use CELL  20
transform 1 0 97 0 -1 126
box 0 0 6 6
use CELL  21
transform -1 0 109 0 -1 68
box 0 0 6 6
use CELL  22
transform 1 0 190 0 1 196
box 0 0 6 6
use CELL  23
transform -1 0 169 0 1 89
box 0 0 6 6
use CELL  24
transform -1 0 158 0 1 120
box 0 0 6 6
use CELL  25
transform -1 0 151 0 1 221
box 0 0 6 6
use CELL  26
transform -1 0 104 0 1 161
box 0 0 6 6
use CELL  27
transform -1 0 137 0 1 196
box 0 0 6 6
use CELL  28
transform -1 0 200 0 -1 167
box 0 0 6 6
use CELL  29
transform -1 0 130 0 1 221
box 0 0 6 6
use CELL  30
transform -1 0 102 0 1 89
box 0 0 6 6
use CELL  31
transform -1 0 111 0 1 161
box 0 0 6 6
use CELL  32
transform -1 0 130 0 1 62
box 0 0 6 6
use CELL  33
transform -1 0 141 0 1 161
box 0 0 6 6
use CELL  34
transform -1 0 109 0 1 89
box 0 0 6 6
use CELL  35
transform -1 0 96 0 1 120
box 0 0 6 6
use CELL  36
transform -1 0 151 0 1 89
box 0 0 6 6
use CELL  37
transform -1 0 160 0 1 221
box 0 0 6 6
use CELL  38
transform -1 0 110 0 1 196
box 0 0 6 6
use CELL  39
transform -1 0 90 0 1 89
box 0 0 6 6
use CELL  40
transform -1 0 97 0 1 161
box 0 0 6 6
use CELL  41
transform -1 0 103 0 1 196
box 0 0 6 6
use CELL  42
transform -1 0 186 0 1 161
box 0 0 6 6
use CELL  43
transform -1 0 178 0 1 89
box 0 0 6 6
use CELL  44
transform -1 0 110 0 1 120
box 0 0 6 6
use CELL  45
transform -1 0 193 0 1 161
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 121 0 1 62
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 130 0 1 89
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 149 0 1 120
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 144 0 1 161
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 125 0 1 196
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 171 0 1 161
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 161 0 1 196
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 164 0 1 196
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 151 0 1 221
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 96 0 1 221
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 121 0 1 221
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 116 0 1 196
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 118 0 1 221
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 122 0 1 196
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 169 0 1 89
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 170 0 1 120
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 118 0 1 62
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 115 0 1 62
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 127 0 1 89
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 125 0 1 120
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 161 0 1 120
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 157 0 1 89
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 156 0 1 161
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 153 0 1 161
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 129 0 1 161
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 173 0 1 196
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 160 0 1 89
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 139 0 1 221
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 142 0 1 221
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 126 0 1 161
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 116 0 1 120
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 115 0 1 89
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 177 0 1 161
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 130 0 1 221
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 146 0 1 196
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 124 0 1 89
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 122 0 1 120
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 141 0 1 161
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 146 0 1 120
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 130 0 1 62
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 142 0 1 89
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 143 0 1 196
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 158 0 1 120
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 139 0 1 89
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 137 0 1 120
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 123 0 1 161
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 121 0 1 89
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 134 0 1 120
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 132 0 1 161
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 128 0 1 196
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 174 0 1 161
box 0 0 3 6
<< metal1 >>
rect 100 53 117 54
rect 103 55 123 56
rect 104 57 120 58
rect 125 57 138 58
rect 128 59 132 60
rect 97 69 120 70
rect 97 71 126 72
rect 100 73 105 74
rect 107 73 141 74
rect 128 75 147 76
rect 116 77 129 78
rect 88 79 117 80
rect 134 79 168 80
rect 144 81 171 82
rect 131 83 144 84
rect 122 85 132 86
rect 85 87 123 88
rect 149 87 159 88
rect 161 87 165 88
rect 85 96 139 97
rect 104 98 144 99
rect 105 100 148 101
rect 108 102 150 103
rect 122 104 136 105
rect 123 106 126 107
rect 126 108 129 109
rect 131 108 151 109
rect 161 108 174 109
rect 156 110 163 111
rect 176 110 182 111
rect 167 112 178 113
rect 164 114 169 115
rect 158 116 166 117
rect 140 118 160 119
rect 85 127 95 128
rect 88 129 106 130
rect 91 131 124 132
rect 95 133 134 134
rect 98 135 131 136
rect 106 137 127 138
rect 108 139 136 140
rect 117 141 128 142
rect 124 143 139 144
rect 139 145 160 146
rect 142 147 148 148
rect 145 149 151 150
rect 156 149 172 150
rect 157 151 185 152
rect 162 153 166 154
rect 154 155 167 156
rect 172 155 178 156
rect 175 157 189 158
rect 178 159 196 160
rect 88 168 92 169
rect 95 168 125 169
rect 99 170 128 171
rect 98 172 118 173
rect 102 174 131 175
rect 109 176 143 177
rect 108 178 148 179
rect 126 180 146 181
rect 129 182 134 183
rect 123 184 133 185
rect 139 184 145 185
rect 150 184 155 185
rect 157 184 170 185
rect 166 186 173 187
rect 162 188 172 189
rect 165 190 169 191
rect 175 190 185 191
rect 174 192 192 193
rect 178 194 189 195
rect 98 203 130 204
rect 94 205 98 206
rect 108 205 127 206
rect 119 207 124 208
rect 117 209 123 210
rect 131 209 148 210
rect 135 211 154 212
rect 140 213 156 214
rect 144 215 159 216
rect 143 217 147 218
rect 152 217 166 218
rect 162 219 169 220
rect 174 219 195 220
rect 97 228 101 229
rect 107 228 120 229
rect 110 230 123 231
rect 125 230 132 231
rect 128 232 144 233
rect 140 234 150 235
rect 152 234 156 235
<< metal2 >>
rect 100 53 101 63
rect 116 53 117 63
rect 103 51 104 56
rect 122 55 123 63
rect 104 57 105 63
rect 119 57 120 63
rect 125 57 126 63
rect 137 57 138 63
rect 128 59 129 63
rect 131 59 132 63
rect 97 67 98 70
rect 119 67 120 70
rect 97 71 98 90
rect 125 71 126 90
rect 100 67 101 74
rect 104 73 105 90
rect 107 73 108 90
rect 140 73 141 90
rect 128 67 129 76
rect 146 75 147 90
rect 116 67 117 78
rect 128 77 129 90
rect 88 79 89 90
rect 116 79 117 90
rect 134 67 135 80
rect 167 79 168 90
rect 144 67 145 82
rect 170 81 171 90
rect 131 67 132 84
rect 143 83 144 90
rect 122 67 123 86
rect 131 85 132 90
rect 85 87 86 90
rect 122 87 123 90
rect 149 87 150 90
rect 158 87 159 90
rect 161 87 162 90
rect 164 87 165 90
rect 85 94 86 97
rect 138 96 139 121
rect 104 94 105 99
rect 143 94 144 99
rect 105 100 106 121
rect 147 100 148 121
rect 108 102 109 121
rect 149 94 150 103
rect 116 94 117 105
rect 117 104 118 121
rect 122 94 123 105
rect 135 104 136 121
rect 123 106 124 121
rect 125 94 126 107
rect 126 108 127 121
rect 128 94 129 109
rect 131 94 132 109
rect 150 108 151 121
rect 161 94 162 109
rect 173 94 174 109
rect 156 110 157 121
rect 162 110 163 121
rect 170 94 171 111
rect 171 110 172 121
rect 176 94 177 111
rect 181 110 182 121
rect 167 94 168 113
rect 177 112 178 121
rect 164 94 165 115
rect 168 114 169 121
rect 158 94 159 117
rect 165 116 166 121
rect 140 94 141 119
rect 159 118 160 121
rect 85 127 86 162
rect 94 125 95 128
rect 88 129 89 162
rect 105 125 106 130
rect 91 125 92 132
rect 123 125 124 132
rect 95 133 96 162
rect 133 133 134 162
rect 98 125 99 136
rect 130 135 131 162
rect 106 137 107 162
rect 126 125 127 138
rect 108 125 109 140
rect 135 125 136 140
rect 117 125 118 142
rect 127 141 128 162
rect 124 143 125 162
rect 138 125 139 144
rect 139 145 140 162
rect 159 125 160 146
rect 142 147 143 162
rect 147 125 148 148
rect 145 149 146 162
rect 150 125 151 150
rect 156 125 157 150
rect 171 125 172 150
rect 157 151 158 162
rect 184 151 185 162
rect 162 125 163 154
rect 165 125 166 154
rect 154 155 155 162
rect 166 155 167 162
rect 172 155 173 162
rect 177 125 178 156
rect 175 157 176 162
rect 188 157 189 162
rect 178 159 179 162
rect 195 159 196 162
rect 88 166 89 169
rect 91 168 92 197
rect 95 166 96 169
rect 124 166 125 169
rect 99 166 100 171
rect 127 166 128 171
rect 98 172 99 197
rect 117 172 118 197
rect 102 166 103 175
rect 130 166 131 175
rect 105 176 106 197
rect 106 166 107 177
rect 109 166 110 177
rect 142 166 143 177
rect 108 178 109 197
rect 147 178 148 197
rect 126 180 127 197
rect 145 166 146 181
rect 129 182 130 197
rect 133 166 134 183
rect 123 184 124 197
rect 132 184 133 197
rect 139 166 140 185
rect 144 184 145 197
rect 150 184 151 197
rect 154 166 155 185
rect 157 166 158 185
rect 169 166 170 185
rect 166 166 167 187
rect 172 166 173 187
rect 162 188 163 197
rect 171 188 172 197
rect 165 190 166 197
rect 168 190 169 197
rect 175 166 176 191
rect 184 166 185 191
rect 174 192 175 197
rect 191 192 192 197
rect 178 166 179 195
rect 188 166 189 195
rect 91 203 92 222
rect 91 201 92 204
rect 98 201 99 204
rect 129 201 130 204
rect 94 205 95 222
rect 97 205 98 222
rect 108 201 109 206
rect 126 201 127 206
rect 119 207 120 222
rect 123 201 124 208
rect 117 201 118 210
rect 122 209 123 222
rect 131 209 132 222
rect 147 201 148 210
rect 135 201 136 212
rect 153 201 154 212
rect 140 213 141 222
rect 155 213 156 222
rect 144 201 145 216
rect 158 215 159 222
rect 143 217 144 222
rect 146 217 147 222
rect 152 217 153 222
rect 165 201 166 218
rect 162 201 163 220
rect 168 201 169 220
rect 174 201 175 220
rect 194 201 195 220
rect 97 226 98 229
rect 100 226 101 229
rect 107 226 108 229
rect 119 226 120 229
rect 110 226 111 231
rect 122 226 123 231
rect 125 226 126 231
rect 131 226 132 231
rect 128 226 129 233
rect 143 226 144 233
rect 140 226 141 235
rect 149 226 150 235
rect 152 226 153 235
rect 155 226 156 235
<< via >>
rect 100 53 101 54
rect 116 53 117 54
rect 103 55 104 56
rect 122 55 123 56
rect 104 57 105 58
rect 119 57 120 58
rect 125 57 126 58
rect 137 57 138 58
rect 128 59 129 60
rect 131 59 132 60
rect 97 69 98 70
rect 119 69 120 70
rect 97 71 98 72
rect 125 71 126 72
rect 100 73 101 74
rect 104 73 105 74
rect 107 73 108 74
rect 140 73 141 74
rect 128 75 129 76
rect 146 75 147 76
rect 116 77 117 78
rect 128 77 129 78
rect 88 79 89 80
rect 116 79 117 80
rect 134 79 135 80
rect 167 79 168 80
rect 144 81 145 82
rect 170 81 171 82
rect 131 83 132 84
rect 143 83 144 84
rect 122 85 123 86
rect 131 85 132 86
rect 85 87 86 88
rect 122 87 123 88
rect 149 87 150 88
rect 158 87 159 88
rect 161 87 162 88
rect 164 87 165 88
rect 85 96 86 97
rect 138 96 139 97
rect 104 98 105 99
rect 143 98 144 99
rect 105 100 106 101
rect 147 100 148 101
rect 108 102 109 103
rect 149 102 150 103
rect 122 104 123 105
rect 135 104 136 105
rect 123 106 124 107
rect 125 106 126 107
rect 126 108 127 109
rect 128 108 129 109
rect 131 108 132 109
rect 150 108 151 109
rect 161 108 162 109
rect 173 108 174 109
rect 156 110 157 111
rect 162 110 163 111
rect 176 110 177 111
rect 181 110 182 111
rect 167 112 168 113
rect 177 112 178 113
rect 164 114 165 115
rect 168 114 169 115
rect 158 116 159 117
rect 165 116 166 117
rect 140 118 141 119
rect 159 118 160 119
rect 85 127 86 128
rect 94 127 95 128
rect 88 129 89 130
rect 105 129 106 130
rect 91 131 92 132
rect 123 131 124 132
rect 95 133 96 134
rect 133 133 134 134
rect 98 135 99 136
rect 130 135 131 136
rect 106 137 107 138
rect 126 137 127 138
rect 108 139 109 140
rect 135 139 136 140
rect 117 141 118 142
rect 127 141 128 142
rect 124 143 125 144
rect 138 143 139 144
rect 139 145 140 146
rect 159 145 160 146
rect 142 147 143 148
rect 147 147 148 148
rect 145 149 146 150
rect 150 149 151 150
rect 156 149 157 150
rect 171 149 172 150
rect 157 151 158 152
rect 184 151 185 152
rect 162 153 163 154
rect 165 153 166 154
rect 154 155 155 156
rect 166 155 167 156
rect 172 155 173 156
rect 177 155 178 156
rect 175 157 176 158
rect 188 157 189 158
rect 178 159 179 160
rect 195 159 196 160
rect 88 168 89 169
rect 91 168 92 169
rect 95 168 96 169
rect 124 168 125 169
rect 99 170 100 171
rect 127 170 128 171
rect 98 172 99 173
rect 117 172 118 173
rect 102 174 103 175
rect 130 174 131 175
rect 109 176 110 177
rect 142 176 143 177
rect 108 178 109 179
rect 147 178 148 179
rect 126 180 127 181
rect 145 180 146 181
rect 129 182 130 183
rect 133 182 134 183
rect 123 184 124 185
rect 132 184 133 185
rect 139 184 140 185
rect 144 184 145 185
rect 150 184 151 185
rect 154 184 155 185
rect 157 184 158 185
rect 169 184 170 185
rect 166 186 167 187
rect 172 186 173 187
rect 162 188 163 189
rect 171 188 172 189
rect 165 190 166 191
rect 168 190 169 191
rect 175 190 176 191
rect 184 190 185 191
rect 174 192 175 193
rect 191 192 192 193
rect 178 194 179 195
rect 188 194 189 195
rect 98 203 99 204
rect 129 203 130 204
rect 94 205 95 206
rect 97 205 98 206
rect 108 205 109 206
rect 126 205 127 206
rect 119 207 120 208
rect 123 207 124 208
rect 117 209 118 210
rect 122 209 123 210
rect 131 209 132 210
rect 147 209 148 210
rect 135 211 136 212
rect 153 211 154 212
rect 140 213 141 214
rect 155 213 156 214
rect 144 215 145 216
rect 158 215 159 216
rect 143 217 144 218
rect 146 217 147 218
rect 152 217 153 218
rect 165 217 166 218
rect 162 219 163 220
rect 168 219 169 220
rect 174 219 175 220
rect 194 219 195 220
rect 97 228 98 229
rect 100 228 101 229
rect 107 228 108 229
rect 119 228 120 229
rect 110 230 111 231
rect 122 230 123 231
rect 125 230 126 231
rect 131 230 132 231
rect 128 232 129 233
rect 143 232 144 233
rect 140 234 141 235
rect 149 234 150 235
rect 152 234 153 235
rect 155 234 156 235
<< end >>
