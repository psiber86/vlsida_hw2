magic
tech scmos
timestamp 1395743089
<< m1p >>
use CELL  1
transform -1 0 2938 0 1 5009
box 0 0 6 6
use CELL  2
transform 1 0 2893 0 1 3775
box 0 0 6 6
use CELL  3
transform -1 0 3603 0 1 6554
box 0 0 6 6
use CELL  4
transform -1 0 2931 0 1 5920
box 0 0 6 6
use CELL  5
transform -1 0 3829 0 1 5318
box 0 0 6 6
use CELL  6
transform -1 0 2923 0 1 4345
box 0 0 6 6
use CELL  7
transform -1 0 3794 0 1 4068
box 0 0 6 6
use CELL  8
transform 1 0 3059 0 1 4658
box 0 0 6 6
use CELL  9
transform -1 0 2936 0 1 8510
box 0 0 6 6
use CELL  10
transform -1 0 3891 0 1 5009
box 0 0 6 6
use CELL  11
transform -1 0 3707 0 1 7849
box 0 0 6 6
use CELL  12
transform -1 0 2933 0 1 1990
box 0 0 6 6
use CELL  13
transform 1 0 2981 0 -1 7395
box 0 0 6 6
use CELL  14
transform -1 0 2925 0 1 6261
box 0 0 6 6
use CELL  15
transform 1 0 3879 0 1 3452
box 0 0 6 6
use CELL  16
transform 1 0 3415 0 1 2667
box 0 0 6 6
use CELL  17
transform -1 0 3681 0 1 7632
box 0 0 6 6
use CELL  18
transform -1 0 3880 0 1 4068
box 0 0 6 6
use CELL  19
transform -1 0 2981 0 1 8510
box 0 0 6 6
use CELL  20
transform 1 0 2862 0 -1 5015
box 0 0 6 6
use CELL  21
transform -1 0 3660 0 1 7389
box 0 0 6 6
use CELL  22
transform -1 0 3638 0 1 7632
box 0 0 6 6
use CELL  23
transform 1 0 3613 0 -1 8102
box 0 0 6 6
use CELL  24
transform -1 0 3773 0 1 3153
box 0 0 6 6
use CELL  25
transform -1 0 2917 0 -1 2217
box 0 0 6 6
use CELL  26
transform 1 0 3247 0 -1 1511
box 0 0 6 6
use CELL  27
transform -1 0 3599 0 1 7849
box 0 0 6 6
use CELL  28
transform -1 0 3409 0 1 8315
box 0 0 6 6
use CELL  29
transform -1 0 3012 0 1 1630
box 0 0 6 6
use CELL  30
transform -1 0 2985 0 1 1783
box 0 0 6 6
use CELL  31
transform -1 0 2963 0 1 3452
box 0 0 6 6
use CELL  32
transform -1 0 3421 0 1 8315
box 0 0 6 6
use CELL  33
transform -1 0 3197 0 1 3153
box 0 0 6 6
use CELL  34
transform -1 0 2924 0 1 5318
box 0 0 6 6
use CELL  35
transform -1 0 3072 0 1 6554
box 0 0 6 6
use CELL  36
transform -1 0 3833 0 1 3775
box 0 0 6 6
use CELL  37
transform -1 0 2969 0 1 6261
box 0 0 6 6
use CELL  38
transform -1 0 3077 0 1 5617
box 0 0 6 6
use CELL  39
transform -1 0 3046 0 1 5009
box 0 0 6 6
use CELL  40
transform 1 0 3028 0 1 1434
box 0 0 6 6
use CELL  41
transform 1 0 2911 0 -1 5015
box 0 0 6 6
use CELL  42
transform -1 0 3749 0 1 3452
box 0 0 6 6
use CELL  43
transform -1 0 2910 0 -1 2930
box 0 0 6 6
use CELL  44
transform -1 0 2886 0 -1 7855
box 0 0 6 6
use CELL  45
transform -1 0 2916 0 1 7389
box 0 0 6 6
use CELL  46
transform -1 0 3023 0 1 5318
box 0 0 6 6
use CELL  47
transform -1 0 3775 0 1 4345
box 0 0 6 6
use CELL  48
transform -1 0 3563 0 1 7389
box 0 0 6 6
use CELL  49
transform -1 0 3574 0 1 1783
box 0 0 6 6
use CELL  50
transform 1 0 3511 0 -1 8321
box 0 0 6 6
use CELL  51
transform -1 0 3791 0 1 6261
box 0 0 6 6
use CELL  52
transform -1 0 2932 0 -1 2673
box 0 0 6 6
use CELL  53
transform -1 0 3786 0 1 6821
box 0 0 6 6
use CELL  54
transform 1 0 3666 0 -1 7395
box 0 0 6 6
use CELL  55
transform 1 0 3909 0 1 4345
box 0 0 6 6
use CELL  56
transform -1 0 3713 0 -1 5324
box 0 0 6 6
use CELL  57
transform -1 0 3422 0 1 8510
box 0 0 6 6
use CELL  58
transform -1 0 3001 0 1 5617
box 0 0 6 6
use CELL  59
transform 1 0 2924 0 -1 8102
box 0 0 6 6
use CELL  60
transform 1 0 2906 0 -1 1996
box 0 0 6 6
use CELL  61
transform -1 0 3073 0 1 6261
box 0 0 6 6
use CELL  62
transform -1 0 3029 0 1 8315
box 0 0 6 6
use CELL  63
transform -1 0 3128 0 1 3452
box 0 0 6 6
use CELL  64
transform -1 0 3554 0 1 8096
box 0 0 6 6
use CELL  65
transform 1 0 3185 0 1 6821
box 0 0 6 6
use CELL  66
transform -1 0 3071 0 1 3153
box 0 0 6 6
use CELL  67
transform -1 0 3178 0 1 2454
box 0 0 6 6
use CELL  68
transform 1 0 3620 0 1 1990
box 0 0 6 6
use CELL  69
transform -1 0 2945 0 1 4658
box 0 0 6 6
use CELL  70
transform 1 0 2964 0 1 5920
box 0 0 6 6
use CELL  71
transform -1 0 3670 0 1 6554
box 0 0 6 6
use CELL  72
transform -1 0 3053 0 1 8734
box 0 0 6 6
use CELL  73
transform -1 0 2995 0 1 3775
box 0 0 6 6
use CELL  74
transform -1 0 3776 0 1 7389
box 0 0 6 6
use CELL  75
transform -1 0 2960 0 -1 2673
box 0 0 6 6
use CELL  76
transform -1 0 3531 0 1 2211
box 0 0 6 6
use CELL  77
transform -1 0 3819 0 1 3775
box 0 0 6 6
use CELL  78
transform -1 0 2908 0 1 4658
box 0 0 6 6
use CELL  79
transform -1 0 2920 0 1 2667
box 0 0 6 6
use CELL  80
transform -1 0 3460 0 1 8315
box 0 0 6 6
use CELL  81
transform -1 0 2976 0 1 4068
box 0 0 6 6
use CELL  82
transform 1 0 3095 0 -1 5623
box 0 0 6 6
use CELL  83
transform -1 0 3868 0 1 6261
box 0 0 6 6
use CELL  84
transform -1 0 3081 0 1 5920
box 0 0 6 6
use CELL  85
transform -1 0 3994 0 1 5920
box 0 0 6 6
use CELL  86
transform -1 0 3035 0 1 5318
box 0 0 6 6
use CELL  87
transform -1 0 3846 0 1 3452
box 0 0 6 6
use CELL  88
transform -1 0 3862 0 1 5617
box 0 0 6 6
use CELL  89
transform -1 0 3950 0 1 4345
box 0 0 6 6
use CELL  90
transform 1 0 3694 0 -1 7855
box 0 0 6 6
use CELL  91
transform -1 0 2887 0 1 4658
box 0 0 6 6
use CELL  92
transform -1 0 3631 0 1 7632
box 0 0 6 6
use CELL  93
transform 1 0 3855 0 -1 6267
box 0 0 6 6
use CELL  94
transform -1 0 3861 0 -1 6560
box 0 0 6 6
use CELL  95
transform 1 0 3877 0 1 5920
box 0 0 6 6
use CELL  96
transform -1 0 3092 0 1 7389
box 0 0 6 6
use CELL  97
transform -1 0 2922 0 1 1505
box 0 0 6 6
use CELL  98
transform -1 0 3898 0 1 5009
box 0 0 6 6
use CELL  99
transform -1 0 3629 0 1 2667
box 0 0 6 6
use CELL  100
transform 1 0 3799 0 1 6821
box 0 0 6 6
use CELL  101
transform 1 0 3689 0 1 7632
box 0 0 6 6
use CELL  102
transform -1 0 3059 0 1 7632
box 0 0 6 6
use CELL  103
transform -1 0 2974 0 1 7632
box 0 0 6 6
use CELL  104
transform -1 0 3357 0 1 6554
box 0 0 6 6
use CELL  105
transform -1 0 2977 0 1 4345
box 0 0 6 6
use CELL  106
transform -1 0 2957 0 1 1505
box 0 0 6 6
use CELL  107
transform -1 0 3873 0 -1 3781
box 0 0 6 6
use CELL  108
transform -1 0 3828 0 1 6261
box 0 0 6 6
use CELL  109
transform 1 0 3487 0 1 1783
box 0 0 6 6
use CELL  110
transform -1 0 3756 0 -1 7855
box 0 0 6 6
use CELL  111
transform -1 0 2936 0 1 7849
box 0 0 6 6
use CELL  112
transform -1 0 3560 0 1 1783
box 0 0 6 6
use CELL  113
transform -1 0 3743 0 1 3775
box 0 0 6 6
use CELL  114
transform -1 0 3779 0 1 6821
box 0 0 6 6
use CELL  115
transform -1 0 2946 0 1 1783
box 0 0 6 6
use CELL  116
transform -1 0 3830 0 1 4658
box 0 0 6 6
use CELL  117
transform 1 0 3049 0 -1 1440
box 0 0 6 6
use CELL  118
transform -1 0 3146 0 -1 7395
box 0 0 6 6
use CELL  119
transform -1 0 3543 0 1 2211
box 0 0 6 6
use CELL  120
transform -1 0 3017 0 1 8734
box 0 0 6 6
use CELL  121
transform -1 0 4008 0 1 5920
box 0 0 6 6
use CELL  122
transform -1 0 3894 0 1 4068
box 0 0 6 6
use CELL  123
transform -1 0 3610 0 1 6554
box 0 0 6 6
use CELL  124
transform -1 0 3232 0 1 5009
box 0 0 6 6
use CELL  125
transform 1 0 3834 0 1 6554
box 0 0 6 6
use CELL  126
transform -1 0 2905 0 1 1990
box 0 0 6 6
use CELL  127
transform -1 0 3828 0 1 6554
box 0 0 6 6
use CELL  128
transform -1 0 2923 0 1 7632
box 0 0 6 6
use CELL  129
transform 1 0 3905 0 1 5009
box 0 0 6 6
use CELL  130
transform 1 0 3768 0 -1 7102
box 0 0 6 6
use CELL  131
transform 1 0 2996 0 -1 8321
box 0 0 6 6
use CELL  132
transform 1 0 2869 0 -1 1996
box 0 0 6 6
use CELL  133
transform -1 0 3115 0 1 8510
box 0 0 6 6
use CELL  134
transform -1 0 3750 0 1 3775
box 0 0 6 6
use CELL  135
transform -1 0 3624 0 1 7632
box 0 0 6 6
use CELL  136
transform -1 0 2979 0 1 2667
box 0 0 6 6
use CELL  137
transform -1 0 3889 0 1 6261
box 0 0 6 6
use CELL  138
transform -1 0 3047 0 1 3153
box 0 0 6 6
use CELL  139
transform -1 0 3011 0 1 6554
box 0 0 6 6
use CELL  140
transform 1 0 2999 0 1 1505
box 0 0 6 6
use CELL  141
transform -1 0 3659 0 1 2211
box 0 0 6 6
use CELL  142
transform -1 0 2948 0 1 7849
box 0 0 6 6
use CELL  143
transform -1 0 3851 0 1 5009
box 0 0 6 6
use CELL  144
transform -1 0 2941 0 1 1630
box 0 0 6 6
use CELL  145
transform 1 0 2977 0 -1 8321
box 0 0 6 6
use CELL  146
transform -1 0 2976 0 1 1630
box 0 0 6 6
use CELL  147
transform -1 0 3044 0 1 1630
box 0 0 6 6
use CELL  148
transform -1 0 2989 0 1 3452
box 0 0 6 6
use CELL  149
transform -1 0 3287 0 1 8510
box 0 0 6 6
use CELL  150
transform -1 0 3108 0 1 2924
box 0 0 6 6
use CELL  151
transform 1 0 3606 0 1 1990
box 0 0 6 6
use CELL  152
transform -1 0 3257 0 1 1783
box 0 0 6 6
use CELL  153
transform -1 0 3813 0 1 4068
box 0 0 6 6
use CELL  154
transform -1 0 2939 0 1 2667
box 0 0 6 6
use CELL  155
transform -1 0 2927 0 1 1783
box 0 0 6 6
use CELL  156
transform 1 0 3147 0 1 8653
box 0 0 6 6
use CELL  157
transform -1 0 3930 0 1 4658
box 0 0 6 6
use CELL  158
transform -1 0 2922 0 1 1630
box 0 0 6 6
use CELL  159
transform -1 0 3723 0 1 2924
box 0 0 6 6
use CELL  160
transform -1 0 3865 0 1 5009
box 0 0 6 6
use CELL  161
transform 1 0 3437 0 1 1630
box 0 0 6 6
use CELL  162
transform -1 0 3144 0 1 4658
box 0 0 6 6
use CELL  163
transform 1 0 3179 0 -1 1511
box 0 0 6 6
use CELL  164
transform -1 0 3830 0 1 5617
box 0 0 6 6
use CELL  165
transform -1 0 3668 0 1 8096
box 0 0 6 6
use CELL  166
transform -1 0 3088 0 1 6261
box 0 0 6 6
use CELL  167
transform -1 0 3051 0 1 8096
box 0 0 6 6
use CELL  168
transform 1 0 3071 0 -1 1511
box 0 0 6 6
use CELL  169
transform -1 0 3622 0 1 2667
box 0 0 6 6
use CELL  170
transform -1 0 3632 0 1 6261
box 0 0 6 6
use CELL  171
transform 1 0 3743 0 1 7849
box 0 0 6 6
use CELL  172
transform -1 0 2874 0 1 4658
box 0 0 6 6
use CELL  173
transform -1 0 2983 0 1 6261
box 0 0 6 6
use CELL  174
transform -1 0 2918 0 1 3452
box 0 0 6 6
use CELL  175
transform 1 0 3625 0 -1 2460
box 0 0 6 6
use CELL  176
transform -1 0 2925 0 1 3452
box 0 0 6 6
use CELL  177
transform -1 0 2990 0 -1 7102
box 0 0 6 6
use CELL  178
transform -1 0 3038 0 1 5920
box 0 0 6 6
use CELL  179
transform -1 0 2930 0 1 7632
box 0 0 6 6
use CELL  180
transform 1 0 3010 0 1 7632
box 0 0 6 6
use CELL  181
transform -1 0 2904 0 1 4345
box 0 0 6 6
use CELL  182
transform -1 0 3840 0 1 3153
box 0 0 6 6
use CELL  183
transform -1 0 2916 0 1 3153
box 0 0 6 6
use CELL  184
transform -1 0 2974 0 1 7096
box 0 0 6 6
use CELL  185
transform -1 0 3760 0 1 7096
box 0 0 6 6
use CELL  186
transform 1 0 3388 0 -1 8516
box 0 0 6 6
use CELL  187
transform -1 0 3354 0 1 1630
box 0 0 6 6
use CELL  188
transform -1 0 2925 0 1 2454
box 0 0 6 6
use CELL  189
transform 1 0 3736 0 1 7849
box 0 0 6 6
use CELL  190
transform -1 0 3588 0 1 2454
box 0 0 6 6
use CELL  191
transform -1 0 2926 0 1 6821
box 0 0 6 6
use CELL  192
transform -1 0 3203 0 1 3452
box 0 0 6 6
use CELL  193
transform -1 0 2905 0 1 4068
box 0 0 6 6
use CELL  194
transform -1 0 3777 0 1 5009
box 0 0 6 6
use CELL  195
transform -1 0 3339 0 1 1990
box 0 0 6 6
use CELL  196
transform -1 0 3757 0 1 3775
box 0 0 6 6
use CELL  197
transform -1 0 3761 0 1 3452
box 0 0 6 6
use CELL  198
transform -1 0 3605 0 1 8096
box 0 0 6 6
use CELL  199
transform -1 0 3028 0 1 2211
box 0 0 6 6
use CELL  200
transform 1 0 3765 0 1 3775
box 0 0 6 6
use CELL  201
transform -1 0 2922 0 1 7849
box 0 0 6 6
use CELL  202
transform 1 0 3007 0 1 1434
box 0 0 6 6
use CELL  203
transform -1 0 3570 0 1 1990
box 0 0 6 6
use CELL  204
transform 1 0 2966 0 -1 2673
box 0 0 6 6
use CELL  205
transform -1 0 2948 0 1 2924
box 0 0 6 6
use CELL  206
transform -1 0 3001 0 1 6261
box 0 0 6 6
use CELL  207
transform -1 0 3154 0 1 2454
box 0 0 6 6
use CELL  208
transform -1 0 3729 0 1 4068
box 0 0 6 6
use CELL  209
transform -1 0 3327 0 1 8510
box 0 0 6 6
use CELL  210
transform -1 0 3703 0 -1 2673
box 0 0 6 6
use CELL  211
transform -1 0 3823 0 1 5617
box 0 0 6 6
use CELL  212
transform -1 0 2868 0 1 1990
box 0 0 6 6
use CELL  213
transform 1 0 3833 0 1 3452
box 0 0 6 6
use CELL  214
transform -1 0 3613 0 1 2454
box 0 0 6 6
use CELL  215
transform 1 0 3131 0 1 8653
box 0 0 6 6
use CELL  216
transform 1 0 3800 0 1 4068
box 0 0 6 6
use CELL  217
transform -1 0 2911 0 1 6261
box 0 0 6 6
use CELL  218
transform -1 0 3029 0 1 2924
box 0 0 6 6
use CELL  219
transform -1 0 3000 0 1 8510
box 0 0 6 6
use CELL  220
transform -1 0 3553 0 1 2454
box 0 0 6 6
use CELL  221
transform -1 0 3753 0 1 4658
box 0 0 6 6
use CELL  222
transform -1 0 3656 0 1 6821
box 0 0 6 6
use CELL  223
transform -1 0 3038 0 1 3775
box 0 0 6 6
use CELL  224
transform -1 0 3813 0 1 3153
box 0 0 6 6
use CELL  225
transform -1 0 3110 0 1 3153
box 0 0 6 6
use CELL  226
transform -1 0 3143 0 -1 1511
box 0 0 6 6
use CELL  227
transform -1 0 3810 0 1 7096
box 0 0 6 6
use CELL  228
transform -1 0 2983 0 1 4068
box 0 0 6 6
use CELL  229
transform 1 0 3655 0 1 8096
box 0 0 6 6
use CELL  230
transform 1 0 2905 0 1 2211
box 0 0 6 6
use CELL  231
transform -1 0 2957 0 1 6261
box 0 0 6 6
use CELL  232
transform 1 0 3777 0 -1 7395
box 0 0 6 6
use CELL  233
transform -1 0 2899 0 1 2667
box 0 0 6 6
use CELL  234
transform 1 0 3530 0 -1 8321
box 0 0 6 6
use CELL  235
transform 1 0 2956 0 -1 4074
box 0 0 6 6
use CELL  236
transform -1 0 3682 0 1 7096
box 0 0 6 6
use CELL  237
transform -1 0 3076 0 -1 1789
box 0 0 6 6
use CELL  238
transform -1 0 3769 0 1 7389
box 0 0 6 6
use CELL  239
transform -1 0 3905 0 1 4658
box 0 0 6 6
use CELL  240
transform -1 0 2957 0 1 6554
box 0 0 6 6
use CELL  241
transform -1 0 3091 0 1 1783
box 0 0 6 6
use CELL  242
transform -1 0 3829 0 -1 7102
box 0 0 6 6
use CELL  243
transform 1 0 3817 0 1 4658
box 0 0 6 6
use CELL  244
transform -1 0 4001 0 1 5920
box 0 0 6 6
use CELL  245
transform 1 0 2936 0 1 7632
box 0 0 6 6
use CELL  246
transform -1 0 3137 0 1 4658
box 0 0 6 6
use CELL  247
transform 1 0 3051 0 -1 5926
box 0 0 6 6
use CELL  248
transform -1 0 3025 0 1 1434
box 0 0 6 6
use CELL  249
transform -1 0 3159 0 1 4658
box 0 0 6 6
use CELL  250
transform -1 0 3769 0 1 7849
box 0 0 6 6
use CELL  251
transform -1 0 3149 0 1 4345
box 0 0 6 6
use CELL  252
transform -1 0 3777 0 1 2924
box 0 0 6 6
use CELL  253
transform -1 0 2983 0 1 6554
box 0 0 6 6
use CELL  254
transform -1 0 2967 0 1 7632
box 0 0 6 6
use CELL  255
transform -1 0 3673 0 1 5009
box 0 0 6 6
use CELL  256
transform 1 0 3755 0 -1 3159
box 0 0 6 6
use CELL  257
transform -1 0 3192 0 1 8653
box 0 0 6 6
use CELL  258
transform -1 0 2997 0 1 2454
box 0 0 6 6
use CELL  259
transform -1 0 3013 0 1 1783
box 0 0 6 6
use CELL  260
transform -1 0 3730 0 1 2924
box 0 0 6 6
use CELL  261
transform -1 0 3857 0 1 7096
box 0 0 6 6
use CELL  262
transform -1 0 2963 0 1 4345
box 0 0 6 6
use CELL  263
transform -1 0 3729 0 1 7632
box 0 0 6 6
use CELL  264
transform 1 0 3743 0 1 2924
box 0 0 6 6
use CELL  265
transform -1 0 2955 0 1 8315
box 0 0 6 6
use CELL  266
transform -1 0 3572 0 1 2454
box 0 0 6 6
use CELL  267
transform -1 0 3094 0 1 7096
box 0 0 6 6
use CELL  268
transform -1 0 3912 0 -1 4664
box 0 0 6 6
use CELL  269
transform -1 0 3696 0 1 2924
box 0 0 6 6
use CELL  270
transform -1 0 2913 0 1 5617
box 0 0 6 6
use CELL  271
transform -1 0 3853 0 1 3452
box 0 0 6 6
use CELL  272
transform -1 0 3213 0 1 4345
box 0 0 6 6
use CELL  273
transform -1 0 3550 0 1 8315
box 0 0 6 6
use CELL  274
transform 1 0 2958 0 1 8734
box 0 0 6 6
use CELL  275
transform 1 0 3750 0 1 2924
box 0 0 6 6
use CELL  276
transform -1 0 2918 0 1 2454
box 0 0 6 6
use CELL  277
transform -1 0 3557 0 1 2211
box 0 0 6 6
use CELL  278
transform -1 0 2974 0 1 5318
box 0 0 6 6
use CELL  279
transform -1 0 3096 0 1 2667
box 0 0 6 6
use CELL  280
transform 1 0 2910 0 -1 8102
box 0 0 6 6
use CELL  281
transform -1 0 2929 0 1 7849
box 0 0 6 6
use CELL  282
transform -1 0 3008 0 1 4658
box 0 0 6 6
use CELL  283
transform 1 0 2874 0 -1 8740
box 0 0 6 6
use CELL  284
transform 1 0 3949 0 -1 5926
box 0 0 6 6
use CELL  285
transform -1 0 2929 0 1 8734
box 0 0 6 6
use CELL  286
transform -1 0 2998 0 1 1505
box 0 0 6 6
use CELL  287
transform 1 0 3461 0 1 1783
box 0 0 6 6
use CELL  288
transform -1 0 3560 0 -1 7638
box 0 0 6 6
use CELL  289
transform -1 0 2980 0 1 8734
box 0 0 6 6
use CELL  290
transform -1 0 3842 0 1 6261
box 0 0 6 6
use CELL  291
transform -1 0 3595 0 1 2454
box 0 0 6 6
use CELL  292
transform 1 0 3820 0 1 6821
box 0 0 6 6
use CELL  293
transform 1 0 2950 0 1 8096
box 0 0 6 6
use CELL  294
transform 1 0 2943 0 1 7096
box 0 0 6 6
use CELL  295
transform 1 0 3570 0 1 2211
box 0 0 6 6
use CELL  296
transform -1 0 3641 0 1 5318
box 0 0 6 6
use CELL  297
transform -1 0 3025 0 1 3452
box 0 0 6 6
use CELL  298
transform -1 0 2906 0 1 1783
box 0 0 6 6
use CELL  299
transform -1 0 3027 0 1 7849
box 0 0 6 6
use CELL  300
transform -1 0 3784 0 1 2924
box 0 0 6 6
use CELL  301
transform 1 0 3730 0 1 3153
box 0 0 6 6
use CELL  302
transform -1 0 3234 0 -1 1511
box 0 0 6 6
use CELL  303
transform -1 0 3877 0 1 5009
box 0 0 6 6
use CELL  304
transform -1 0 2977 0 1 8096
box 0 0 6 6
use CELL  305
transform 1 0 3013 0 1 4345
box 0 0 6 6
use CELL  306
transform 1 0 2966 0 1 2454
box 0 0 6 6
use CELL  307
transform -1 0 3677 0 1 6821
box 0 0 6 6
use CELL  308
transform 1 0 2931 0 -1 8102
box 0 0 6 6
use CELL  309
transform -1 0 2981 0 1 2924
box 0 0 6 6
use CELL  310
transform 1 0 3676 0 -1 2460
box 0 0 6 6
use CELL  311
transform -1 0 2958 0 1 3775
box 0 0 6 6
use CELL  312
transform -1 0 3828 0 1 4345
box 0 0 6 6
use CELL  313
transform -1 0 2976 0 1 6261
box 0 0 6 6
use CELL  314
transform -1 0 3030 0 1 8096
box 0 0 6 6
use CELL  315
transform 1 0 2944 0 1 2211
box 0 0 6 6
use CELL  316
transform 1 0 3202 0 -1 8659
box 0 0 6 6
use CELL  317
transform 1 0 3921 0 -1 4074
box 0 0 6 6
use CELL  318
transform -1 0 2880 0 1 6554
box 0 0 6 6
use CELL  319
transform -1 0 3891 0 1 4658
box 0 0 6 6
use CELL  320
transform 1 0 2944 0 1 5318
box 0 0 6 6
use CELL  321
transform 1 0 3746 0 1 2667
box 0 0 6 6
use CELL  322
transform -1 0 2898 0 1 5009
box 0 0 6 6
use CELL  323
transform -1 0 3826 0 1 3775
box 0 0 6 6
use CELL  324
transform -1 0 3764 0 1 6554
box 0 0 6 6
use CELL  325
transform -1 0 3801 0 1 5318
box 0 0 6 6
use CELL  326
transform -1 0 3816 0 1 5617
box 0 0 6 6
use CELL  327
transform -1 0 3032 0 1 5009
box 0 0 6 6
use CELL  328
transform 1 0 3087 0 1 2211
box 0 0 6 6
use CELL  329
transform -1 0 3777 0 1 6261
box 0 0 6 6
use CELL  330
transform 1 0 3682 0 -1 7638
box 0 0 6 6
use CELL  331
transform -1 0 3365 0 1 1783
box 0 0 6 6
use CELL  332
transform -1 0 3662 0 1 3153
box 0 0 6 6
use CELL  333
transform -1 0 3176 0 1 8653
box 0 0 6 6
use CELL  334
transform -1 0 3050 0 1 4068
box 0 0 6 6
use CELL  335
transform -1 0 2981 0 1 7096
box 0 0 6 6
use CELL  336
transform -1 0 3734 0 1 5318
box 0 0 6 6
use CELL  337
transform -1 0 2944 0 1 3775
box 0 0 6 6
use CELL  338
transform -1 0 3645 0 1 2667
box 0 0 6 6
use CELL  339
transform 1 0 3844 0 1 7096
box 0 0 6 6
use CELL  340
transform 1 0 2887 0 1 1783
box 0 0 6 6
use CELL  341
transform -1 0 2982 0 1 1990
box 0 0 6 6
use CELL  342
transform 1 0 3721 0 1 7389
box 0 0 6 6
use CELL  343
transform -1 0 3917 0 1 5009
box 0 0 6 6
use CELL  344
transform -1 0 3708 0 1 7389
box 0 0 6 6
use CELL  345
transform -1 0 2905 0 -1 5015
box 0 0 6 6
use CELL  346
transform -1 0 3655 0 1 7849
box 0 0 6 6
use CELL  347
transform -1 0 3007 0 1 3452
box 0 0 6 6
use CELL  348
transform -1 0 3784 0 1 6261
box 0 0 6 6
use CELL  349
transform -1 0 3294 0 1 8510
box 0 0 6 6
use CELL  350
transform -1 0 2962 0 1 7849
box 0 0 6 6
use CELL  351
transform 1 0 2964 0 1 4345
box 0 0 6 6
use CELL  352
transform 1 0 3207 0 1 1505
box 0 0 6 6
use CELL  353
transform -1 0 3794 0 1 5318
box 0 0 6 6
use CELL  354
transform -1 0 2965 0 1 2211
box 0 0 6 6
use CELL  355
transform -1 0 3809 0 -1 4351
box 0 0 6 6
use CELL  356
transform -1 0 2923 0 1 7389
box 0 0 6 6
use CELL  357
transform 1 0 3401 0 1 5318
box 0 0 6 6
use CELL  358
transform -1 0 3013 0 1 5920
box 0 0 6 6
use CELL  359
transform -1 0 2820 0 1 8510
box 0 0 6 6
use CELL  360
transform -1 0 2988 0 1 7632
box 0 0 6 6
use CELL  361
transform -1 0 3550 0 1 2211
box 0 0 6 6
use CELL  362
transform 1 0 2914 0 -1 5623
box 0 0 6 6
use CELL  363
transform -1 0 3929 0 1 4345
box 0 0 6 6
use CELL  364
transform -1 0 3869 0 1 5318
box 0 0 6 6
use CELL  365
transform -1 0 2965 0 1 3775
box 0 0 6 6
use CELL  366
transform -1 0 2955 0 1 1434
box 0 0 6 6
use CELL  367
transform 1 0 2904 0 1 5920
box 0 0 6 6
use CELL  368
transform -1 0 2936 0 1 2211
box 0 0 6 6
use CELL  369
transform -1 0 3741 0 1 4345
box 0 0 6 6
use CELL  370
transform 1 0 3347 0 1 8510
box 0 0 6 6
use CELL  371
transform -1 0 3162 0 1 2924
box 0 0 6 6
use CELL  372
transform -1 0 3537 0 -1 1996
box 0 0 6 6
use CELL  373
transform -1 0 3037 0 1 1630
box 0 0 6 6
use CELL  374
transform -1 0 3062 0 1 7389
box 0 0 6 6
use CELL  375
transform -1 0 2955 0 1 4068
box 0 0 6 6
use CELL  376
transform -1 0 2886 0 1 1783
box 0 0 6 6
use CELL  377
transform 1 0 3066 0 1 2924
box 0 0 6 6
use CELL  378
transform -1 0 3806 0 1 3153
box 0 0 6 6
use CELL  379
transform 1 0 3928 0 -1 4074
box 0 0 6 6
use CELL  380
transform -1 0 2917 0 1 5920
box 0 0 6 6
use CELL  381
transform 1 0 3395 0 -1 8516
box 0 0 6 6
use CELL  382
transform -1 0 3738 0 1 2667
box 0 0 6 6
use CELL  383
transform -1 0 2918 0 1 6261
box 0 0 6 6
use CELL  384
transform 1 0 2913 0 1 1990
box 0 0 6 6
use CELL  385
transform 1 0 3959 0 -1 4664
box 0 0 6 6
use CELL  386
transform -1 0 2998 0 1 8653
box 0 0 6 6
use CELL  387
transform -1 0 3771 0 1 6554
box 0 0 6 6
use CELL  388
transform 1 0 3721 0 1 6554
box 0 0 6 6
use CELL  389
transform -1 0 3039 0 1 6554
box 0 0 6 6
use CELL  390
transform -1 0 3866 0 1 6821
box 0 0 6 6
use CELL  391
transform -1 0 3005 0 1 5318
box 0 0 6 6
use CELL  392
transform -1 0 3041 0 1 2924
box 0 0 6 6
use CELL  393
transform -1 0 3731 0 -1 2673
box 0 0 6 6
use CELL  394
transform 1 0 2935 0 1 2454
box 0 0 6 6
use CELL  395
transform -1 0 2898 0 1 6821
box 0 0 6 6
use CELL  396
transform -1 0 3095 0 1 6261
box 0 0 6 6
use CELL  397
transform -1 0 2963 0 1 1990
box 0 0 6 6
use CELL  398
transform -1 0 2939 0 1 5617
box 0 0 6 6
use CELL  399
transform 1 0 3487 0 1 8315
box 0 0 6 6
use CELL  400
transform -1 0 3647 0 1 8096
box 0 0 6 6
use CELL  401
transform -1 0 3029 0 1 4658
box 0 0 6 6
use CELL  402
transform -1 0 2887 0 1 8734
box 0 0 6 6
use CELL  403
transform -1 0 2992 0 1 1783
box 0 0 6 6
use CELL  404
transform -1 0 3889 0 1 5617
box 0 0 6 6
use CELL  405
transform -1 0 3887 0 1 4068
box 0 0 6 6
use CELL  406
transform -1 0 2904 0 1 6261
box 0 0 6 6
use CELL  407
transform 1 0 2942 0 1 8315
box 0 0 6 6
use CELL  408
transform -1 0 3020 0 1 5920
box 0 0 6 6
use CELL  409
transform -1 0 2962 0 1 1434
box 0 0 6 6
use CELL  410
transform -1 0 2962 0 1 1630
box 0 0 6 6
use CELL  411
transform -1 0 3114 0 1 1990
box 0 0 6 6
use CELL  412
transform -1 0 2957 0 1 6821
box 0 0 6 6
use CELL  413
transform -1 0 3103 0 1 2454
box 0 0 6 6
use CELL  414
transform -1 0 3028 0 1 5617
box 0 0 6 6
use CELL  415
transform 1 0 3769 0 1 3452
box 0 0 6 6
use CELL  416
transform -1 0 3702 0 1 7632
box 0 0 6 6
use CELL  417
transform -1 0 3748 0 1 5617
box 0 0 6 6
use CELL  418
transform 1 0 3711 0 1 2667
box 0 0 6 6
use CELL  419
transform -1 0 2904 0 1 2211
box 0 0 6 6
use CELL  420
transform -1 0 3610 0 1 2667
box 0 0 6 6
use CELL  421
transform -1 0 3837 0 1 5617
box 0 0 6 6
use CELL  422
transform -1 0 3787 0 1 4068
box 0 0 6 6
use CELL  423
transform 1 0 3177 0 -1 8659
box 0 0 6 6
use CELL  424
transform 1 0 2808 0 1 4345
box 0 0 6 6
use CELL  425
transform -1 0 2974 0 1 8510
box 0 0 6 6
use CELL  426
transform -1 0 2912 0 1 6821
box 0 0 6 6
use CELL  427
transform -1 0 3714 0 1 7849
box 0 0 6 6
use CELL  428
transform -1 0 3707 0 1 6261
box 0 0 6 6
use CELL  429
transform -1 0 2936 0 1 8315
box 0 0 6 6
use CELL  430
transform -1 0 3792 0 1 5920
box 0 0 6 6
use CELL  431
transform -1 0 3241 0 1 1505
box 0 0 6 6
use CELL  432
transform -1 0 3116 0 1 1783
box 0 0 6 6
use CELL  433
transform -1 0 3859 0 1 3775
box 0 0 6 6
use CELL  434
transform -1 0 3956 0 1 4345
box 0 0 6 6
use CELL  435
transform -1 0 3616 0 1 7096
box 0 0 6 6
use CELL  436
transform -1 0 3653 0 1 7389
box 0 0 6 6
use CELL  437
transform -1 0 3654 0 -1 8102
box 0 0 6 6
use CELL  438
transform 1 0 2926 0 1 3775
box 0 0 6 6
use CELL  439
transform 1 0 3702 0 1 2924
box 0 0 6 6
use CELL  440
transform 1 0 2894 0 1 5617
box 0 0 6 6
use CELL  441
transform -1 0 2962 0 1 8510
box 0 0 6 6
use CELL  442
transform -1 0 3641 0 1 7849
box 0 0 6 6
use CELL  443
transform -1 0 2911 0 1 3452
box 0 0 6 6
use CELL  444
transform 1 0 3613 0 1 1990
box 0 0 6 6
use CELL  445
transform -1 0 3515 0 1 7849
box 0 0 6 6
use CELL  446
transform -1 0 3346 0 1 8510
box 0 0 6 6
use CELL  447
transform -1 0 2970 0 1 3452
box 0 0 6 6
use CELL  448
transform -1 0 3113 0 1 5318
box 0 0 6 6
use CELL  449
transform 1 0 2922 0 1 8653
box 0 0 6 6
use CELL  450
transform 1 0 3865 0 1 3452
box 0 0 6 6
use CELL  451
transform 1 0 2954 0 1 7632
box 0 0 6 6
use CELL  452
transform -1 0 3039 0 1 5009
box 0 0 6 6
use CELL  453
transform -1 0 3130 0 1 8653
box 0 0 6 6
use CELL  454
transform -1 0 2922 0 1 8315
box 0 0 6 6
use CELL  455
transform 1 0 3541 0 -1 8102
box 0 0 6 6
use CELL  456
transform 1 0 3494 0 1 1783
box 0 0 6 6
use CELL  457
transform 1 0 4029 0 1 5920
box 0 0 6 6
use CELL  458
transform 1 0 3531 0 1 1783
box 0 0 6 6
use CELL  459
transform -1 0 2950 0 1 6261
box 0 0 6 6
use CELL  460
transform -1 0 2924 0 1 5920
box 0 0 6 6
use CELL  461
transform -1 0 3009 0 1 1990
box 0 0 6 6
use CELL  462
transform -1 0 3019 0 1 4068
box 0 0 6 6
use CELL  463
transform -1 0 3044 0 1 4345
box 0 0 6 6
use CELL  464
transform 1 0 3517 0 1 1783
box 0 0 6 6
use CELL  465
transform -1 0 2893 0 1 5617
box 0 0 6 6
use CELL  466
transform -1 0 3985 0 -1 4664
box 0 0 6 6
use CELL  467
transform 1 0 2965 0 1 5009
box 0 0 6 6
use CELL  468
transform -1 0 3913 0 1 5920
box 0 0 6 6
use CELL  469
transform -1 0 3047 0 1 4658
box 0 0 6 6
use CELL  470
transform 1 0 3710 0 1 7632
box 0 0 6 6
use CELL  471
transform -1 0 2924 0 1 5009
box 0 0 6 6
use CELL  472
transform -1 0 2935 0 1 3153
box 0 0 6 6
use CELL  473
transform 1 0 3592 0 1 1990
box 0 0 6 6
use CELL  474
transform -1 0 2956 0 1 5920
box 0 0 6 6
use CELL  475
transform -1 0 3847 0 1 6554
box 0 0 6 6
use CELL  476
transform -1 0 2963 0 1 8096
box 0 0 6 6
use CELL  477
transform -1 0 2892 0 1 5920
box 0 0 6 6
use CELL  478
transform -1 0 2884 0 1 5009
box 0 0 6 6
use CELL  479
transform -1 0 3819 0 1 6821
box 0 0 6 6
use CELL  480
transform -1 0 3645 0 1 7632
box 0 0 6 6
use CELL  481
transform -1 0 3581 0 1 2454
box 0 0 6 6
use CELL  482
transform -1 0 2937 0 1 4345
box 0 0 6 6
use CELL  483
transform -1 0 2956 0 1 4345
box 0 0 6 6
use CELL  484
transform -1 0 2920 0 1 1783
box 0 0 6 6
use CELL  485
transform 1 0 3718 0 1 2667
box 0 0 6 6
use CELL  486
transform -1 0 2904 0 -1 3458
box 0 0 6 6
use CELL  487
transform -1 0 3192 0 1 1505
box 0 0 6 6
use CELL  488
transform -1 0 3255 0 1 1990
box 0 0 6 6
use CELL  489
transform -1 0 2929 0 -1 1511
box 0 0 6 6
use CELL  490
transform -1 0 2892 0 1 4345
box 0 0 6 6
use CELL  491
transform -1 0 2920 0 -1 4664
box 0 0 6 6
use CELL  492
transform -1 0 2904 0 -1 3159
box 0 0 6 6
use CELL  493
transform -1 0 3723 0 1 7632
box 0 0 6 6
use CELL  494
transform -1 0 3920 0 1 4068
box 0 0 6 6
use CELL  495
transform -1 0 3091 0 1 2454
box 0 0 6 6
use CELL  496
transform 1 0 3545 0 1 1783
box 0 0 6 6
use CELL  497
transform 1 0 2994 0 -1 7855
box 0 0 6 6
use CELL  498
transform 1 0 3132 0 1 4068
box 0 0 6 6
use CELL  499
transform -1 0 3745 0 1 2667
box 0 0 6 6
use CELL  500
transform -1 0 3590 0 1 2211
box 0 0 6 6
use CELL  501
transform -1 0 3767 0 1 7096
box 0 0 6 6
use CELL  502
transform -1 0 3736 0 1 4068
box 0 0 6 6
use CELL  503
transform -1 0 3683 0 1 3153
box 0 0 6 6
use CELL  504
transform -1 0 3679 0 1 5617
box 0 0 6 6
use CELL  505
transform -1 0 2937 0 1 3452
box 0 0 6 6
use CELL  506
transform 1 0 3503 0 1 1783
box 0 0 6 6
use CELL  507
transform -1 0 3641 0 1 2211
box 0 0 6 6
use CELL  508
transform -1 0 3666 0 1 2211
box 0 0 6 6
use CELL  509
transform -1 0 3752 0 1 5009
box 0 0 6 6
use CELL  510
transform -1 0 3640 0 1 8096
box 0 0 6 6
use CELL  511
transform 1 0 3756 0 1 7849
box 0 0 6 6
use CELL  512
transform -1 0 3064 0 1 8653
box 0 0 6 6
use CELL  513
transform -1 0 4022 0 1 5920
box 0 0 6 6
use CELL  514
transform -1 0 3227 0 1 1505
box 0 0 6 6
use CELL  515
transform 1 0 2885 0 -1 5015
box 0 0 6 6
use CELL  516
transform -1 0 3451 0 1 5009
box 0 0 6 6
use CELL  517
transform -1 0 2936 0 1 2924
box 0 0 6 6
use CELL  518
transform 1 0 2886 0 1 2667
box 0 0 6 6
use CELL  519
transform -1 0 3690 0 1 3153
box 0 0 6 6
use CELL  520
transform -1 0 2958 0 1 5617
box 0 0 6 6
use CELL  521
transform -1 0 3674 0 1 6261
box 0 0 6 6
use CELL  522
transform 1 0 3774 0 -1 3159
box 0 0 6 6
use CELL  523
transform -1 0 3714 0 1 3153
box 0 0 6 6
use CELL  524
transform -1 0 3160 0 -1 8659
box 0 0 6 6
use CELL  525
transform -1 0 3855 0 1 5617
box 0 0 6 6
use CELL  526
transform -1 0 2949 0 1 3452
box 0 0 6 6
use CELL  527
transform -1 0 3822 0 1 5318
box 0 0 6 6
use CELL  528
transform 1 0 3872 0 1 7096
box 0 0 6 6
use CELL  529
transform -1 0 2993 0 1 8510
box 0 0 6 6
use CELL  530
transform -1 0 2912 0 1 4068
box 0 0 6 6
use CELL  531
transform 1 0 3620 0 1 8096
box 0 0 6 6
use CELL  532
transform -1 0 2899 0 1 1783
box 0 0 6 6
use CELL  533
transform -1 0 3479 0 1 1783
box 0 0 6 6
use CELL  534
transform -1 0 3840 0 1 3775
box 0 0 6 6
use CELL  535
transform -1 0 3763 0 -1 2930
box 0 0 6 6
use CELL  536
transform -1 0 3075 0 1 1630
box 0 0 6 6
use CELL  537
transform -1 0 3735 0 1 7849
box 0 0 6 6
use CELL  538
transform 1 0 3430 0 1 1630
box 0 0 6 6
use CELL  539
transform 1 0 3592 0 1 8096
box 0 0 6 6
use CELL  540
transform -1 0 4015 0 1 5920
box 0 0 6 6
use CELL  541
transform -1 0 2950 0 1 6554
box 0 0 6 6
use CELL  542
transform -1 0 3701 0 1 3775
box 0 0 6 6
use CELL  543
transform -1 0 3008 0 1 5009
box 0 0 6 6
use CELL  544
transform -1 0 3011 0 1 7389
box 0 0 6 6
use CELL  545
transform -1 0 3791 0 -1 2930
box 0 0 6 6
use CELL  546
transform -1 0 3904 0 1 5009
box 0 0 6 6
use CELL  547
transform -1 0 3780 0 1 5617
box 0 0 6 6
use CELL  548
transform -1 0 3670 0 1 7849
box 0 0 6 6
use CELL  549
transform -1 0 2912 0 1 6554
box 0 0 6 6
use CELL  550
transform 1 0 3666 0 1 5617
box 0 0 6 6
use CELL  551
transform 1 0 2965 0 -1 1440
box 0 0 6 6
use CELL  552
transform -1 0 2929 0 1 2211
box 0 0 6 6
use CELL  553
transform -1 0 3052 0 1 7632
box 0 0 6 6
use CELL  554
transform -1 0 3557 0 1 8315
box 0 0 6 6
use CELL  555
transform -1 0 3943 0 1 4345
box 0 0 6 6
use CELL  556
transform -1 0 3937 0 1 5920
box 0 0 6 6
use CELL  557
transform -1 0 2947 0 1 3153
box 0 0 6 6
use CELL  558
transform -1 0 3051 0 1 1630
box 0 0 6 6
use CELL  559
transform -1 0 3962 0 1 5920
box 0 0 6 6
use CELL  560
transform -1 0 2943 0 1 4068
box 0 0 6 6
use CELL  561
transform -1 0 3059 0 1 5318
box 0 0 6 6
use CELL  562
transform -1 0 3675 0 1 2454
box 0 0 6 6
use CELL  563
transform -1 0 3876 0 1 4345
box 0 0 6 6
use CELL  564
transform -1 0 2917 0 1 7096
box 0 0 6 6
use CELL  565
transform -1 0 3046 0 1 7096
box 0 0 6 6
use CELL  566
transform -1 0 3171 0 1 1990
box 0 0 6 6
use CELL  567
transform -1 0 2901 0 1 4658
box 0 0 6 6
use CELL  568
transform -1 0 3035 0 1 2211
box 0 0 6 6
use CELL  569
transform -1 0 2956 0 1 7096
box 0 0 6 6
use CELL  570
transform -1 0 2996 0 1 8096
box 0 0 6 6
use CELL  571
transform -1 0 2937 0 1 7389
box 0 0 6 6
use CELL  572
transform -1 0 3560 0 1 2454
box 0 0 6 6
use CELL  573
transform 1 0 3857 0 -1 5324
box 0 0 6 6
use CELL  574
transform -1 0 2978 0 1 7389
box 0 0 6 6
use CELL  575
transform 1 0 2856 0 1 5920
box 0 0 6 6
use CELL  576
transform -1 0 3757 0 1 6554
box 0 0 6 6
use CELL  577
transform -1 0 2931 0 -1 5324
box 0 0 6 6
use CELL  578
transform -1 0 3652 0 1 2454
box 0 0 6 6
use CELL  579
transform -1 0 2881 0 1 4658
box 0 0 6 6
use CELL  580
transform -1 0 2886 0 -1 5623
box 0 0 6 6
use CELL  581
transform -1 0 3787 0 1 3153
box 0 0 6 6
use CELL  582
transform 1 0 3606 0 1 8096
box 0 0 6 6
use CELL  583
transform -1 0 3131 0 1 6261
box 0 0 6 6
use CELL  584
transform 1 0 2957 0 1 5920
box 0 0 6 6
use CELL  585
transform -1 0 3164 0 -1 1511
box 0 0 6 6
use CELL  586
transform 1 0 3359 0 -1 3781
box 0 0 6 6
use CELL  587
transform -1 0 2911 0 1 4345
box 0 0 6 6
use CELL  588
transform -1 0 3807 0 1 6554
box 0 0 6 6
use CELL  589
transform -1 0 2976 0 1 6554
box 0 0 6 6
use CELL  590
transform -1 0 2969 0 1 7849
box 0 0 6 6
use CELL  591
transform -1 0 3709 0 1 7632
box 0 0 6 6
use CELL  592
transform -1 0 3866 0 1 3775
box 0 0 6 6
use CELL  593
transform -1 0 3228 0 1 5617
box 0 0 6 6
use CELL  594
transform -1 0 3394 0 1 2454
box 0 0 6 6
use CELL  595
transform -1 0 2976 0 1 6821
box 0 0 6 6
use CELL  596
transform -1 0 2964 0 1 1783
box 0 0 6 6
use CELL  597
transform -1 0 3564 0 1 8315
box 0 0 6 6
use CELL  598
transform -1 0 3366 0 1 1630
box 0 0 6 6
use CELL  599
transform -1 0 3802 0 1 4345
box 0 0 6 6
use CELL  600
transform 1 0 3367 0 1 1630
box 0 0 6 6
use CELL  601
transform -1 0 2990 0 1 2454
box 0 0 6 6
use CELL  602
transform -1 0 3876 0 1 5617
box 0 0 6 6
use CELL  603
transform 1 0 2963 0 1 1630
box 0 0 6 6
use CELL  604
transform -1 0 3858 0 1 5009
box 0 0 6 6
use CELL  605
transform -1 0 3951 0 1 4658
box 0 0 6 6
use CELL  606
transform -1 0 2967 0 1 2924
box 0 0 6 6
use CELL  607
transform -1 0 3126 0 1 2667
box 0 0 6 6
use CELL  608
transform -1 0 3563 0 1 1990
box 0 0 6 6
use CELL  609
transform -1 0 3015 0 1 2667
box 0 0 6 6
use CELL  610
transform -1 0 3882 0 -1 6267
box 0 0 6 6
use CELL  611
transform -1 0 2959 0 1 4658
box 0 0 6 6
use CELL  612
transform -1 0 2956 0 1 3452
box 0 0 6 6
use CELL  613
transform -1 0 3936 0 1 4345
box 0 0 6 6
use CELL  614
transform -1 0 2980 0 1 3153
box 0 0 6 6
use CELL  615
transform -1 0 2964 0 1 7389
box 0 0 6 6
use CELL  616
transform -1 0 2989 0 1 1505
box 0 0 6 6
use CELL  617
transform -1 0 2964 0 1 6821
box 0 0 6 6
use CELL  618
transform 1 0 3010 0 1 3153
box 0 0 6 6
use CELL  619
transform 1 0 3645 0 -1 1996
box 0 0 6 6
use CELL  620
transform -1 0 3782 0 1 3452
box 0 0 6 6
use CELL  621
transform 1 0 2900 0 -1 5623
box 0 0 6 6
use CELL  622
transform -1 0 3845 0 1 6821
box 0 0 6 6
use CELL  623
transform -1 0 2995 0 1 8734
box 0 0 6 6
use CELL  624
transform -1 0 3386 0 1 7389
box 0 0 6 6
use CELL  625
transform 1 0 2808 0 -1 7638
box 0 0 6 6
use CELL  626
transform -1 0 2906 0 1 3775
box 0 0 6 6
use CELL  627
transform -1 0 3748 0 1 7096
box 0 0 6 6
use CELL  628
transform -1 0 3060 0 1 8734
box 0 0 6 6
use CELL  629
transform -1 0 2929 0 1 8510
box 0 0 6 6
use CELL  630
transform -1 0 3901 0 1 4068
box 0 0 6 6
use CELL  631
transform 1 0 2984 0 1 6554
box 0 0 6 6
use CELL  632
transform -1 0 2935 0 1 8653
box 0 0 6 6
use CELL  633
transform 1 0 3627 0 1 8096
box 0 0 6 6
use CELL  634
transform -1 0 2910 0 1 7096
box 0 0 6 6
use CELL  635
transform -1 0 2893 0 1 7849
box 0 0 6 6
use CELL  636
transform -1 0 3667 0 1 2924
box 0 0 6 6
use CELL  637
transform -1 0 3125 0 1 7849
box 0 0 6 6
use CELL  638
transform -1 0 3167 0 1 7849
box 0 0 6 6
use CELL  639
transform -1 0 2951 0 1 3775
box 0 0 6 6
use CELL  640
transform -1 0 3489 0 1 8096
box 0 0 6 6
use CELL  641
transform -1 0 3687 0 -1 2673
box 0 0 6 6
use CELL  642
transform 1 0 3749 0 1 7389
box 0 0 6 6
use CELL  643
transform 1 0 3891 0 1 4345
box 0 0 6 6
use CELL  644
transform -1 0 3727 0 1 5318
box 0 0 6 6
use CELL  645
transform -1 0 2990 0 1 6821
box 0 0 6 6
use CELL  646
transform -1 0 2977 0 1 5617
box 0 0 6 6
use CELL  647
transform -1 0 3663 0 1 2667
box 0 0 6 6
use CELL  648
transform -1 0 3019 0 1 6261
box 0 0 6 6
use CELL  649
transform -1 0 2924 0 1 2924
box 0 0 6 6
use CELL  650
transform 1 0 3435 0 1 1990
box 0 0 6 6
use CELL  651
transform -1 0 2999 0 1 2924
box 0 0 6 6
use CELL  652
transform -1 0 2923 0 1 3153
box 0 0 6 6
use CELL  653
transform -1 0 3114 0 -1 8102
box 0 0 6 6
use CELL  654
transform -1 0 3084 0 -1 2460
box 0 0 6 6
use CELL  655
transform -1 0 2975 0 1 1505
box 0 0 6 6
use CELL  656
transform -1 0 2926 0 1 1990
box 0 0 6 6
use CELL  657
transform -1 0 3025 0 1 8510
box 0 0 6 6
use CELL  658
transform 1 0 3193 0 1 1505
box 0 0 6 6
use CELL  659
transform -1 0 3715 0 -1 7395
box 0 0 6 6
use CELL  660
transform 1 0 3820 0 1 3153
box 0 0 6 6
use CELL  661
transform 1 0 3480 0 -1 1789
box 0 0 6 6
use CELL  662
transform -1 0 3048 0 1 2924
box 0 0 6 6
use CELL  663
transform -1 0 3039 0 1 7096
box 0 0 6 6
use CELL  664
transform -1 0 3206 0 -1 1511
box 0 0 6 6
use CELL  665
transform -1 0 2827 0 -1 3781
box 0 0 6 6
use CELL  666
transform -1 0 3540 0 1 8096
box 0 0 6 6
use CELL  667
transform -1 0 3019 0 1 3775
box 0 0 6 6
use CELL  668
transform 1 0 3033 0 1 8096
box 0 0 6 6
use CELL  669
transform -1 0 2930 0 1 4345
box 0 0 6 6
use CELL  670
transform 1 0 2943 0 1 8096
box 0 0 6 6
use CELL  671
transform -1 0 2874 0 1 6261
box 0 0 6 6
use CELL  672
transform -1 0 2970 0 1 5617
box 0 0 6 6
use CELL  673
transform -1 0 3878 0 1 3452
box 0 0 6 6
use CELL  674
transform -1 0 3339 0 1 8510
box 0 0 6 6
use CELL  675
transform 1 0 3132 0 -1 2673
box 0 0 6 6
use CELL  676
transform -1 0 3864 0 1 7096
box 0 0 6 6
use CELL  677
transform 1 0 2999 0 1 8096
box 0 0 6 6
use CELL  678
transform -1 0 2927 0 1 5617
box 0 0 6 6
use CELL  679
transform -1 0 3871 0 1 7096
box 0 0 6 6
use CELL  680
transform -1 0 3895 0 1 5920
box 0 0 6 6
use CELL  681
transform -1 0 3105 0 1 2211
box 0 0 6 6
use CELL  682
transform 1 0 3715 0 -1 7855
box 0 0 6 6
use CELL  683
transform -1 0 2969 0 1 4068
box 0 0 6 6
use CELL  684
transform -1 0 3605 0 -1 1996
box 0 0 6 6
use CELL  685
transform -1 0 3582 0 1 1990
box 0 0 6 6
use CELL  686
transform -1 0 3793 0 1 6821
box 0 0 6 6
use CELL  687
transform 1 0 3621 0 1 2211
box 0 0 6 6
use CELL  688
transform 1 0 3957 0 -1 4351
box 0 0 6 6
use CELL  689
transform -1 0 3062 0 1 2211
box 0 0 6 6
use CELL  690
transform -1 0 3843 0 1 7096
box 0 0 6 6
use CELL  691
transform 1 0 3543 0 -1 1996
box 0 0 6 6
use CELL  692
transform -1 0 3156 0 1 4345
box 0 0 6 6
use CELL  693
transform 1 0 3814 0 1 3153
box 0 0 6 6
use CELL  694
transform 1 0 3476 0 1 3775
box 0 0 6 6
use CELL  695
transform -1 0 3837 0 1 4658
box 0 0 6 6
use CELL  696
transform -1 0 3002 0 1 8734
box 0 0 6 6
use CELL  697
transform 1 0 3819 0 1 3452
box 0 0 6 6
use CELL  698
transform -1 0 2974 0 1 2924
box 0 0 6 6
use CELL  699
transform -1 0 2920 0 1 3775
box 0 0 6 6
use CELL  700
transform -1 0 3937 0 1 4658
box 0 0 6 6
use CELL  701
transform 1 0 3952 0 -1 4664
box 0 0 6 6
use CELL  702
transform -1 0 3857 0 1 5318
box 0 0 6 6
use CELL  703
transform -1 0 4029 0 1 5920
box 0 0 6 6
use CELL  704
transform 1 0 2937 0 1 2211
box 0 0 6 6
use CELL  705
transform -1 0 2949 0 1 5920
box 0 0 6 6
use CELL  706
transform -1 0 2982 0 1 3452
box 0 0 6 6
use CELL  707
transform -1 0 3030 0 1 1630
box 0 0 6 6
use CELL  708
transform -1 0 2916 0 1 7632
box 0 0 6 6
use CELL  709
transform -1 0 3010 0 -1 2217
box 0 0 6 6
use CELL  710
transform -1 0 2969 0 1 6554
box 0 0 6 6
use CELL  711
transform -1 0 3694 0 1 2667
box 0 0 6 6
use CELL  712
transform -1 0 2898 0 1 1990
box 0 0 6 6
use CELL  713
transform -1 0 3689 0 1 2924
box 0 0 6 6
use CELL  714
transform -1 0 2899 0 -1 6560
box 0 0 6 6
use CELL  715
transform -1 0 3784 0 1 5009
box 0 0 6 6
use CELL  716
transform -1 0 3714 0 1 6261
box 0 0 6 6
use CELL  717
transform -1 0 3764 0 1 3775
box 0 0 6 6
use CELL  718
transform 1 0 3863 0 1 5617
box 0 0 6 6
use CELL  719
transform -1 0 2886 0 1 3775
box 0 0 6 6
use CELL  720
transform -1 0 2893 0 1 8653
box 0 0 6 6
use CELL  721
transform -1 0 3070 0 -1 1440
box 0 0 6 6
use CELL  722
transform -1 0 3149 0 1 5318
box 0 0 6 6
use CELL  723
transform 1 0 3630 0 -1 2673
box 0 0 6 6
use CELL  724
transform 1 0 2972 0 1 5009
box 0 0 6 6
use CELL  725
transform 1 0 3562 0 1 8096
box 0 0 6 6
use CELL  726
transform -1 0 3257 0 1 3452
box 0 0 6 6
use CELL  727
transform -1 0 3450 0 -1 1636
box 0 0 6 6
use CELL  728
transform -1 0 3408 0 -1 8516
box 0 0 6 6
use CELL  729
transform -1 0 3754 0 1 3153
box 0 0 6 6
use CELL  730
transform 1 0 2907 0 1 2667
box 0 0 6 6
use CELL  731
transform 1 0 3722 0 1 7849
box 0 0 6 6
use CELL  732
transform -1 0 2952 0 1 5009
box 0 0 6 6
use CELL  733
transform 1 0 3808 0 1 6554
box 0 0 6 6
use CELL  734
transform -1 0 3783 0 -1 6560
box 0 0 6 6
use CELL  735
transform -1 0 2997 0 1 6821
box 0 0 6 6
use CELL  736
transform -1 0 3713 0 1 3775
box 0 0 6 6
use CELL  737
transform -1 0 3025 0 -1 6827
box 0 0 6 6
use CELL  738
transform 1 0 2983 0 -1 8102
box 0 0 6 6
use CELL  739
transform -1 0 3948 0 1 4068
box 0 0 6 6
use CELL  740
transform -1 0 2906 0 1 2667
box 0 0 6 6
use CELL  741
transform 1 0 2956 0 1 8315
box 0 0 6 6
use CELL  742
transform -1 0 3134 0 1 7389
box 0 0 6 6
use CELL  743
transform -1 0 2946 0 1 5617
box 0 0 6 6
use CELL  744
transform -1 0 2923 0 1 8096
box 0 0 6 6
use CELL  745
transform -1 0 3047 0 1 3775
box 0 0 6 6
use CELL  746
transform 1 0 2892 0 1 7096
box 0 0 6 6
use CELL  747
transform -1 0 3821 0 1 6554
box 0 0 6 6
use CELL  748
transform -1 0 2904 0 1 1630
box 0 0 6 6
use CELL  749
transform 1 0 2991 0 -1 7102
box 0 0 6 6
use CELL  750
transform -1 0 3874 0 1 6554
box 0 0 6 6
use CELL  751
transform -1 0 3654 0 1 5617
box 0 0 6 6
use CELL  752
transform -1 0 3725 0 1 3452
box 0 0 6 6
use CELL  753
transform -1 0 3583 0 1 2211
box 0 0 6 6
use CELL  754
transform -1 0 3876 0 1 5920
box 0 0 6 6
use CELL  755
transform -1 0 3195 0 1 1630
box 0 0 6 6
use CELL  756
transform -1 0 3202 0 1 7096
box 0 0 6 6
use CELL  757
transform -1 0 3770 0 1 5009
box 0 0 6 6
use CELL  758
transform 1 0 3116 0 1 5318
box 0 0 6 6
use CELL  759
transform 1 0 3907 0 -1 4074
box 0 0 6 6
use CELL  760
transform -1 0 2961 0 1 8653
box 0 0 6 6
use CELL  761
transform 1 0 3963 0 1 5920
box 0 0 6 6
use CELL  762
transform -1 0 3898 0 1 4658
box 0 0 6 6
use CELL  763
transform -1 0 3749 0 1 6821
box 0 0 6 6
use CELL  764
transform -1 0 3323 0 1 7632
box 0 0 6 6
use CELL  765
transform -1 0 2936 0 1 1505
box 0 0 6 6
use CELL  766
transform -1 0 3479 0 1 8315
box 0 0 6 6
use CELL  767
transform -1 0 3380 0 1 1630
box 0 0 6 6
use CELL  768
transform -1 0 2995 0 1 2211
box 0 0 6 6
use CELL  769
transform -1 0 3843 0 1 5318
box 0 0 6 6
use CELL  770
transform -1 0 3847 0 1 3775
box 0 0 6 6
use CELL  771
transform -1 0 2955 0 1 2924
box 0 0 6 6
use CELL  772
transform -1 0 3859 0 1 6821
box 0 0 6 6
use CELL  773
transform -1 0 3043 0 1 4068
box 0 0 6 6
use CELL  774
transform -1 0 3972 0 1 4658
box 0 0 6 6
use CELL  775
transform -1 0 3883 0 -1 5623
box 0 0 6 6
use CELL  776
transform -1 0 2892 0 1 6554
box 0 0 6 6
use CELL  777
transform -1 0 2917 0 1 5318
box 0 0 6 6
use CELL  778
transform -1 0 2919 0 1 6554
box 0 0 6 6
use CELL  779
transform -1 0 3798 0 1 6261
box 0 0 6 6
use CELL  780
transform -1 0 3922 0 1 4345
box 0 0 6 6
use CELL  781
transform -1 0 3129 0 1 4068
box 0 0 6 6
use CELL  782
transform -1 0 3836 0 1 5318
box 0 0 6 6
use CELL  783
transform -1 0 3108 0 1 5617
box 0 0 6 6
use CELL  784
transform -1 0 2948 0 -1 2460
box 0 0 6 6
use CELL  785
transform -1 0 2932 0 -1 2460
box 0 0 6 6
use CELL  786
transform -1 0 2930 0 1 7389
box 0 0 6 6
use CELL  787
transform 1 0 3388 0 1 1630
box 0 0 6 6
use CELL  788
transform -1 0 3741 0 1 4658
box 0 0 6 6
use CELL  789
transform -1 0 3873 0 1 4068
box 0 0 6 6
use CELL  790
transform 1 0 3662 0 1 2454
box 0 0 6 6
use CELL  791
transform -1 0 3191 0 1 7849
box 0 0 6 6
use CELL  792
transform -1 0 2970 0 1 1990
box 0 0 6 6
use CELL  793
transform -1 0 3387 0 1 1630
box 0 0 6 6
use CELL  794
transform 1 0 2971 0 -1 8659
box 0 0 6 6
use CELL  795
transform -1 0 3018 0 1 6821
box 0 0 6 6
use CELL  796
transform -1 0 3875 0 1 6261
box 0 0 6 6
use CELL  797
transform 1 0 3669 0 1 2667
box 0 0 6 6
use CELL  798
transform 1 0 3638 0 1 1990
box 0 0 6 6
use CELL  799
transform -1 0 3833 0 1 3153
box 0 0 6 6
use CELL  800
transform -1 0 2995 0 1 8315
box 0 0 6 6
use CELL  801
transform -1 0 3720 0 1 5318
box 0 0 6 6
use CELL  802
transform -1 0 2926 0 1 6554
box 0 0 6 6
use CELL  803
transform -1 0 3868 0 1 6554
box 0 0 6 6
use CELL  804
transform 1 0 2927 0 -1 6827
box 0 0 6 6
use CELL  805
transform -1 0 2981 0 1 5318
box 0 0 6 6
use CELL  806
transform 1 0 3749 0 1 5617
box 0 0 6 6
use CELL  807
transform 1 0 3970 0 1 5920
box 0 0 6 6
use CELL  808
transform -1 0 3030 0 1 1990
box 0 0 6 6
use CELL  809
transform 1 0 3014 0 -1 8321
box 0 0 6 6
use CELL  810
transform -1 0 3679 0 1 2211
box 0 0 6 6
use CELL  811
transform -1 0 3422 0 1 1630
box 0 0 6 6
use CELL  812
transform -1 0 2955 0 1 7389
box 0 0 6 6
use CELL  813
transform -1 0 2995 0 1 5920
box 0 0 6 6
use CELL  814
transform -1 0 3037 0 1 4345
box 0 0 6 6
use CELL  815
transform -1 0 3760 0 1 4068
box 0 0 6 6
use CELL  816
transform -1 0 3816 0 1 4658
box 0 0 6 6
use CELL  817
transform 1 0 3012 0 -1 6560
box 0 0 6 6
use CELL  818
transform 1 0 3689 0 -1 5324
box 0 0 6 6
use CELL  819
transform -1 0 3084 0 1 2924
box 0 0 6 6
use CELL  820
transform -1 0 2954 0 1 8653
box 0 0 6 6
use CELL  821
transform -1 0 3408 0 1 1630
box 0 0 6 6
use CELL  822
transform -1 0 2971 0 1 7389
box 0 0 6 6
use CELL  823
transform -1 0 2953 0 1 2667
box 0 0 6 6
use CELL  824
transform -1 0 2919 0 1 6821
box 0 0 6 6
use CELL  825
transform -1 0 3073 0 1 8653
box 0 0 6 6
use CELL  826
transform -1 0 2911 0 1 2454
box 0 0 6 6
use CELL  827
transform -1 0 3741 0 1 7389
box 0 0 6 6
use CELL  828
transform -1 0 3648 0 1 7849
box 0 0 6 6
use CELL  829
transform -1 0 3036 0 1 8315
box 0 0 6 6
use CELL  830
transform 1 0 3354 0 -1 8516
box 0 0 6 6
use CELL  831
transform -1 0 3524 0 1 8315
box 0 0 6 6
use CELL  832
transform -1 0 3041 0 1 1505
box 0 0 6 6
use CELL  833
transform -1 0 2943 0 1 1505
box 0 0 6 6
use CELL  834
transform 1 0 3935 0 1 4068
box 0 0 6 6
use CELL  835
transform -1 0 2949 0 1 4345
box 0 0 6 6
use CELL  836
transform -1 0 2929 0 1 8315
box 0 0 6 6
use CELL  837
transform -1 0 3530 0 1 1783
box 0 0 6 6
use CELL  838
transform -1 0 2894 0 1 4658
box 0 0 6 6
use CELL  839
transform -1 0 3009 0 1 2454
box 0 0 6 6
use CELL  840
transform -1 0 3849 0 1 6261
box 0 0 6 6
use CELL  841
transform -1 0 3023 0 1 8096
box 0 0 6 6
use CELL  842
transform 1 0 2940 0 -1 1440
box 0 0 6 6
use CELL  843
transform -1 0 2945 0 1 5009
box 0 0 6 6
use CELL  844
transform -1 0 2905 0 1 6821
box 0 0 6 6
use CELL  845
transform -1 0 3822 0 1 7096
box 0 0 6 6
use CELL  846
transform -1 0 3748 0 1 4345
box 0 0 6 6
use CELL  847
transform -1 0 3144 0 1 8653
box 0 0 6 6
use CELL  848
transform -1 0 2924 0 1 7096
box 0 0 6 6
use CELL  849
transform -1 0 3169 0 1 8653
box 0 0 6 6
use CELL  850
transform -1 0 2938 0 1 4658
box 0 0 6 6
use CELL  851
transform -1 0 3680 0 1 5009
box 0 0 6 6
use CELL  852
transform -1 0 2955 0 1 8510
box 0 0 6 6
use CELL  853
transform -1 0 3000 0 1 1630
box 0 0 6 6
use CELL  854
transform -1 0 2881 0 1 6261
box 0 0 6 6
use CELL  855
transform 1 0 3628 0 1 2211
box 0 0 6 6
use CELL  856
transform -1 0 3057 0 1 4068
box 0 0 6 6
use CELL  857
transform -1 0 2913 0 1 3775
box 0 0 6 6
use CELL  858
transform -1 0 3385 0 1 8510
box 0 0 6 6
use CELL  859
transform -1 0 3486 0 1 8315
box 0 0 6 6
use CELL  860
transform 1 0 2970 0 1 7849
box 0 0 6 6
use CELL  861
transform -1 0 2966 0 1 3153
box 0 0 6 6
use CELL  862
transform -1 0 2973 0 1 3153
box 0 0 6 6
use CELL  863
transform -1 0 3660 0 1 2924
box 0 0 6 6
use CELL  864
transform -1 0 3337 0 1 7096
box 0 0 6 6
use CELL  865
transform 1 0 3263 0 1 7632
box 0 0 6 6
use CELL  866
transform -1 0 3047 0 1 7389
box 0 0 6 6
use CELL  867
transform -1 0 2934 0 1 1783
box 0 0 6 6
use CELL  868
transform -1 0 3050 0 1 5920
box 0 0 6 6
use CELL  869
transform -1 0 3567 0 1 1783
box 0 0 6 6
use CELL  870
transform -1 0 2954 0 -1 3159
box 0 0 6 6
use CELL  871
transform -1 0 2947 0 1 8653
box 0 0 6 6
use CELL  872
transform -1 0 3032 0 1 3452
box 0 0 6 6
use CELL  873
transform 1 0 3878 0 1 5009
box 0 0 6 6
use CELL  874
transform 1 0 2983 0 -1 8659
box 0 0 6 6
use CELL  875
transform -1 0 3098 0 1 1783
box 0 0 6 6
use CELL  876
transform -1 0 3560 0 1 3775
box 0 0 6 6
use CELL  877
transform 1 0 3025 0 1 3775
box 0 0 6 6
use CELL  878
transform -1 0 3852 0 1 6821
box 0 0 6 6
use CELL  879
transform -1 0 2898 0 1 4068
box 0 0 6 6
use CELL  880
transform -1 0 2905 0 -1 6560
box 0 0 6 6
use CELL  881
transform -1 0 3062 0 1 4345
box 0 0 6 6
use CELL  882
transform 1 0 3742 0 -1 7395
box 0 0 6 6
use CELL  883
transform -1 0 3729 0 1 3153
box 0 0 6 6
use CELL  884
transform -1 0 3043 0 1 8315
box 0 0 6 6
use CELL  885
transform -1 0 2910 0 1 5318
box 0 0 6 6
use CELL  886
transform -1 0 3220 0 1 1505
box 0 0 6 6
use CELL  887
transform -1 0 2931 0 1 4068
box 0 0 6 6
use CELL  888
transform -1 0 3617 0 1 7632
box 0 0 6 6
use CELL  889
transform -1 0 2974 0 1 8315
box 0 0 6 6
use CELL  890
transform 1 0 2975 0 1 7632
box 0 0 6 6
use CELL  891
transform -1 0 3883 0 1 4345
box 0 0 6 6
use CELL  892
transform 1 0 3241 0 -1 1511
box 0 0 6 6
use CELL  893
transform -1 0 2924 0 1 4068
box 0 0 6 6
use CELL  894
transform 1 0 3021 0 -1 2673
box 0 0 6 6
use CELL  895
transform -1 0 2917 0 1 2924
box 0 0 6 6
use CELL  896
transform -1 0 3433 0 1 5009
box 0 0 6 6
use CELL  897
transform 1 0 2923 0 1 1630
box 0 0 6 6
use CELL  898
transform -1 0 2946 0 1 2667
box 0 0 6 6
use CELL  899
transform 1 0 2958 0 1 5009
box 0 0 6 6
use CELL  900
transform -1 0 3419 0 1 7632
box 0 0 6 6
use CELL  901
transform -1 0 3944 0 1 4658
box 0 0 6 6
use CELL  902
transform -1 0 3029 0 1 8734
box 0 0 6 6
use CELL  903
transform -1 0 3516 0 1 1783
box 0 0 6 6
use CELL  904
transform 1 0 2880 0 1 8653
box 0 0 6 6
use CELL  905
transform -1 0 2989 0 1 1434
box 0 0 6 6
use CELL  906
transform -1 0 3798 0 1 2924
box 0 0 6 6
use CELL  907
transform -1 0 3122 0 1 3153
box 0 0 6 6
use CELL  908
transform -1 0 3890 0 1 4345
box 0 0 6 6
use CELL  909
transform 1 0 2916 0 -1 8740
box 0 0 6 6
use CELL  910
transform -1 0 3770 0 1 2924
box 0 0 6 6
use CELL  911
transform -1 0 3789 0 1 3452
box 0 0 6 6
use CELL  912
transform -1 0 3835 0 1 6261
box 0 0 6 6
use CELL  913
transform -1 0 2970 0 1 8096
box 0 0 6 6
use CELL  914
transform -1 0 3768 0 1 3452
box 0 0 6 6
use CELL  915
transform -1 0 2932 0 1 6261
box 0 0 6 6
use CELL  916
transform -1 0 3122 0 1 8510
box 0 0 6 6
use CELL  917
transform -1 0 3836 0 1 7096
box 0 0 6 6
use CELL  918
transform 1 0 3550 0 -1 1996
box 0 0 6 6
use CELL  919
transform -1 0 2998 0 1 3153
box 0 0 6 6
use CELL  920
transform -1 0 2982 0 1 1505
box 0 0 6 6
use CELL  921
transform -1 0 3838 0 -1 6827
box 0 0 6 6
use CELL  922
transform 1 0 3756 0 -1 7395
box 0 0 6 6
use CELL  923
transform -1 0 3808 0 1 5318
box 0 0 6 6
use CELL  924
transform 1 0 3409 0 1 8510
box 0 0 6 6
use CELL  925
transform -1 0 2962 0 1 5318
box 0 0 6 6
use CELL  926
transform -1 0 3620 0 -1 2217
box 0 0 6 6
use CELL  927
transform -1 0 3815 0 1 5318
box 0 0 6 6
use CELL  928
transform -1 0 3032 0 1 6821
box 0 0 6 6
use CELL  929
transform -1 0 4042 0 -1 5926
box 0 0 6 6
use CELL  930
transform -1 0 3672 0 1 2211
box 0 0 6 6
use CELL  931
transform -1 0 3201 0 -1 8659
box 0 0 6 6
use CELL  932
transform -1 0 3069 0 -1 2217
box 0 0 6 6
use CELL  933
transform -1 0 3734 0 1 7389
box 0 0 6 6
use CELL  934
transform 1 0 3537 0 1 8315
box 0 0 6 6
use CELL  935
transform -1 0 3145 0 1 2667
box 0 0 6 6
use CELL  936
transform -1 0 3979 0 1 4658
box 0 0 6 6
use CELL  937
transform 1 0 2944 0 1 1505
box 0 0 6 6
use CELL  938
transform -1 0 3378 0 1 8510
box 0 0 6 6
use CELL  939
transform -1 0 3035 0 1 5617
box 0 0 6 6
use CELL  940
transform -1 0 3018 0 1 1990
box 0 0 6 6
use CELL  941
transform -1 0 2893 0 1 3775
box 0 0 6 6
use CELL  942
transform -1 0 2983 0 1 6821
box 0 0 6 6
use CELL  943
transform 1 0 2949 0 1 7849
box 0 0 6 6
use CELL  944
transform -1 0 2977 0 1 5920
box 0 0 6 6
use CELL  945
transform -1 0 3007 0 1 8510
box 0 0 6 6
use CELL  946
transform -1 0 2880 0 -1 3458
box 0 0 6 6
use CELL  947
transform 1 0 3423 0 1 1630
box 0 0 6 6
use CELL  948
transform -1 0 3569 0 1 2211
box 0 0 6 6
use CELL  949
transform -1 0 3777 0 1 4658
box 0 0 6 6
use CELL  950
transform 1 0 3395 0 1 1630
box 0 0 6 6
use CELL  951
transform 1 0 3585 0 1 1990
box 0 0 6 6
use CELL  952
transform -1 0 3821 0 1 4345
box 0 0 6 6
use CELL  953
transform -1 0 2943 0 -1 5324
box 0 0 6 6
use CELL  954
transform -1 0 3174 0 1 4068
box 0 0 6 6
use CELL  955
transform -1 0 3762 0 1 5617
box 0 0 6 6
use CELL  956
transform -1 0 2931 0 1 7096
box 0 0 6 6
use CELL  957
transform 1 0 3655 0 1 2454
box 0 0 6 6
use CELL  958
transform -1 0 3068 0 1 6821
box 0 0 6 6
use CELL  959
transform -1 0 3713 0 1 5009
box 0 0 6 6
use CELL  960
transform -1 0 3090 0 1 6554
box 0 0 6 6
use CELL  961
transform -1 0 2952 0 1 4658
box 0 0 6 6
use CELL  962
transform -1 0 2973 0 1 8734
box 0 0 6 6
use CELL  963
transform -1 0 3854 0 1 6554
box 0 0 6 6
use CELL  964
transform -1 0 3341 0 1 6821
box 0 0 6 6
use CELL  965
transform 1 0 3704 0 1 2667
box 0 0 6 6
use CELL  966
transform -1 0 3658 0 1 1990
box 0 0 6 6
use CELL  967
transform -1 0 2966 0 1 4658
box 0 0 6 6
use CELL  968
transform -1 0 3076 0 1 7096
box 0 0 6 6
use CELL  969
transform 1 0 3058 0 1 1434
box 0 0 6 6
use CELL  970
transform -1 0 3832 0 1 3452
box 0 0 6 6
use CELL  971
transform -1 0 2931 0 1 5009
box 0 0 6 6
use CELL  972
transform -1 0 3040 0 1 3153
box 0 0 6 6
use CELL  973
transform 1 0 3555 0 -1 8102
box 0 0 6 6
use CELL  974
transform -1 0 2970 0 1 8653
box 0 0 6 6
use CELL  975
transform -1 0 3799 0 1 3153
box 0 0 6 6
use CELL  976
transform 1 0 3035 0 -1 7855
box 0 0 6 6
use CELL  977
transform -1 0 3034 0 1 7849
box 0 0 6 6
use CELL  978
transform -1 0 3472 0 1 8315
box 0 0 6 6
use CELL  979
transform -1 0 3844 0 1 5009
box 0 0 6 6
use CELL  980
transform 1 0 3409 0 -1 1636
box 0 0 6 6
use CELL  981
transform 1 0 2869 0 -1 5015
box 0 0 6 6
use CELL  982
transform 1 0 3759 0 1 5920
box 0 0 6 6
use CELL  983
transform -1 0 3141 0 1 1990
box 0 0 6 6
use CELL  984
transform -1 0 3850 0 1 5318
box 0 0 6 6
use CELL  985
transform -1 0 3645 0 -1 2460
box 0 0 6 6
use CELL  986
transform -1 0 3614 0 1 6821
box 0 0 6 6
use CELL  987
transform -1 0 3899 0 1 3452
box 0 0 6 6
use CELL  988
transform 1 0 3538 0 1 1783
box 0 0 6 6
use CELL  989
transform -1 0 3812 0 1 6821
box 0 0 6 6
use CELL  990
transform 1 0 2814 0 1 3775
box 0 0 6 6
use CELL  991
transform 1 0 2920 0 -1 4664
box 0 0 6 6
use CELL  992
transform 1 0 3886 0 -1 3458
box 0 0 6 6
use CELL  993
transform -1 0 3009 0 1 7632
box 0 0 6 6
use CELL  994
transform -1 0 2922 0 1 8510
box 0 0 6 6
use CELL  995
transform -1 0 2904 0 1 2454
box 0 0 6 6
use CELL  996
transform -1 0 3674 0 1 2924
box 0 0 6 6
use CELL  997
transform 1 0 2937 0 1 8510
box 0 0 6 6
use CELL  998
transform 1 0 2907 0 1 1783
box 0 0 6 6
use CELL  999
transform 1 0 3731 0 1 2924
box 0 0 6 6
use CELL  1000
transform -1 0 3638 0 -1 2460
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 3068 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 3207 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 3402 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 3248 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 3060 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 3035 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 3250 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 3080 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 3351 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 3336 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 3224 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 3272 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 3287 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 3288 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 3330 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 3324 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 3056 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 3148 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 3593 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 3598 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 3347 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 3383 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 3413 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 3363 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 3295 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 3272 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 3638 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 3546 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 3609 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 3299 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 3556 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 3366 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 3465 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 3468 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 3620 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 3698 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 3494 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 3489 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 3562 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 3526 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 3384 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 3519 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 3449 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 2937 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 2938 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 2932 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 2939 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 3843 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 3982 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 3846 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 3985 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 3849 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 3828 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 3826 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 3865 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 3912 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 3897 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 3432 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 3050 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 3104 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 3086 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 3087 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 3060 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 3016 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 3166 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 3192 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 3248 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 3224 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 3203 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 3918 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 3903 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 3901 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 3847 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 3853 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 3787 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 3670 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 3651 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 3715 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 3810 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 3654 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 3063 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 3293 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 3286 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 3164 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 3294 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 3296 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 3474 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 3159 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 3218 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 3319 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 3408 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 3228 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 3438 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 3120 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 3110 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 3085 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 3239 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 3236 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 3859 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 3658 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 3861 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 3783 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 3789 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 3736 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 3711 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 3675 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 3613 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 3864 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-109
transform 1 0 3852 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-110
transform 1 0 3855 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-111
transform 1 0 3808 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-112
transform 1 0 3770 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-113
transform 1 0 3792 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-114
transform 1 0 3937 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-115
transform 1 0 3804 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-116
transform 1 0 3789 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-117
transform 1 0 3097 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-118
transform 1 0 3117 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-119
transform 1 0 3116 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-120
transform 1 0 3134 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-121
transform 1 0 2993 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-122
transform 1 0 3009 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-123
transform 1 0 3006 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-124
transform 1 0 2999 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-125
transform 1 0 2875 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-126
transform 1 0 3641 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-127
transform 1 0 3644 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-128
transform 1 0 3724 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-129
transform 1 0 3581 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-130
transform 1 0 3572 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-131
transform 1 0 3569 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-132
transform 1 0 3477 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-133
transform 1 0 3448 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-134
transform 1 0 3315 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-135
transform 1 0 3611 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-136
transform 1 0 3528 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-137
transform 1 0 3635 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-138
transform 1 0 3748 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-139
transform 1 0 3749 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-140
transform 1 0 3568 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-141
transform 1 0 3524 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-142
transform 1 0 3385 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-143
transform 1 0 3192 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-144
transform 1 0 3813 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-145
transform 1 0 3807 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-146
transform 1 0 3855 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-147
transform 1 0 3864 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-148
transform 1 0 3879 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-149
transform 1 0 3832 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-150
transform 1 0 3782 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-151
transform 1 0 3804 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-152
transform 1 0 3943 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-153
transform 1 0 3816 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-154
transform 1 0 3795 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-155
transform 1 0 3793 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-156
transform 1 0 3798 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-157
transform 1 0 3660 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-158
transform 1 0 3816 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-159
transform 1 0 3810 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-160
transform 1 0 3858 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-161
transform 1 0 3867 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-162
transform 1 0 3882 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-163
transform 1 0 3835 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-164
transform 1 0 3785 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-165
transform 1 0 3807 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-166
transform 1 0 3742 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-167
transform 1 0 3795 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-168
transform 1 0 3789 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-169
transform 1 0 3837 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-170
transform 1 0 3051 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-171
transform 1 0 3038 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-172
transform 1 0 2939 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-173
transform 1 0 3462 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-174
transform 1 0 3459 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-175
transform 1 0 3409 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-176
transform 1 0 3542 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-177
transform 1 0 3551 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-178
transform 1 0 3652 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-179
transform 1 0 3626 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-180
transform 1 0 3658 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-181
transform 1 0 3695 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-182
transform 1 0 3777 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-183
transform 1 0 3275 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-184
transform 1 0 3115 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-185
transform 1 0 3067 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-186
transform 1 0 3138 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-187
transform 1 0 3088 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-188
transform 1 0 3227 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-189
transform 1 0 3206 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-190
transform 1 0 3240 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-191
transform 1 0 3019 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-192
transform 1 0 3094 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-193
transform 1 0 3129 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-194
transform 1 0 3117 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-195
transform 1 0 3146 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-196
transform 1 0 3236 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-197
transform 1 0 3146 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-198
transform 1 0 3031 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-199
transform 1 0 3025 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-200
transform 1 0 3017 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-201
transform 1 0 3020 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-202
transform 1 0 3011 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-203
transform 1 0 3007 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-204
transform 1 0 3001 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-205
transform 1 0 3007 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-206
transform 1 0 3061 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-207
transform 1 0 3015 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-208
transform 1 0 2966 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-209
transform 1 0 2946 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-210
transform 1 0 3228 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-211
transform 1 0 3339 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-212
transform 1 0 3283 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-213
transform 1 0 3346 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-214
transform 1 0 3429 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-215
transform 1 0 3311 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-216
transform 1 0 3266 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-217
transform 1 0 3414 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-218
transform 1 0 3423 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-219
transform 1 0 3468 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-220
transform 1 0 3337 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-221
transform 1 0 3323 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-222
transform 1 0 3219 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-223
transform 1 0 2971 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-224
transform 1 0 2989 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-225
transform 1 0 2983 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-226
transform 1 0 2972 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-227
transform 1 0 3314 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-228
transform 1 0 2977 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-229
transform 1 0 2995 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-230
transform 1 0 3368 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-231
transform 1 0 3324 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-232
transform 1 0 3274 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-233
transform 1 0 3262 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-234
transform 1 0 3187 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-235
transform 1 0 3315 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-236
transform 1 0 3701 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-237
transform 1 0 3623 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-238
transform 1 0 3222 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-239
transform 1 0 3333 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-240
transform 1 0 3261 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-241
transform 1 0 3559 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-242
transform 1 0 3230 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-243
transform 1 0 3612 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-244
transform 1 0 3384 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-245
transform 1 0 3277 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-246
transform 1 0 3281 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-247
transform 1 0 3171 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-248
transform 1 0 3332 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-249
transform 1 0 3340 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-250
transform 1 0 3245 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-251
transform 1 0 3170 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-252
transform 1 0 3128 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-253
transform 1 0 3342 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-254
transform 1 0 3155 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-255
transform 1 0 3148 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-256
transform 1 0 3122 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-257
transform 1 0 3137 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-258
transform 1 0 3107 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-259
transform 1 0 3819 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-260
transform 1 0 3834 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-261
transform 1 0 3843 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-262
transform 1 0 3802 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-263
transform 1 0 3758 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-264
transform 1 0 3786 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-265
transform 1 0 3946 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-266
transform 1 0 3819 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-267
transform 1 0 3798 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-268
transform 1 0 3777 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-269
transform 1 0 3813 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-270
transform 1 0 3098 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-271
transform 1 0 3147 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-272
transform 1 0 2983 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-273
transform 1 0 2987 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-274
transform 1 0 2990 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-275
transform 1 0 2978 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-276
transform 1 0 2995 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-277
transform 1 0 2989 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-278
transform 1 0 2990 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-279
transform 1 0 2983 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-280
transform 1 0 2989 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-281
transform 1 0 2993 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-282
transform 1 0 2996 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-283
transform 1 0 2996 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-284
transform 1 0 3007 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-285
transform 1 0 3007 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-286
transform 1 0 3416 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-287
transform 1 0 3376 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-288
transform 1 0 3285 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-289
transform 1 0 3522 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-290
transform 1 0 3070 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-291
transform 1 0 3507 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-292
transform 1 0 3525 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-293
transform 1 0 3504 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-294
transform 1 0 3368 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-295
transform 1 0 3374 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-296
transform 1 0 3139 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-297
transform 1 0 3125 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-298
transform 1 0 3131 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-299
transform 1 0 3111 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-300
transform 1 0 3137 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-301
transform 1 0 3056 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-302
transform 1 0 3163 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-303
transform 1 0 3025 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-304
transform 1 0 3092 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-305
transform 1 0 3259 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-306
transform 1 0 3311 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-307
transform 1 0 3183 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-308
transform 1 0 3629 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-309
transform 1 0 3464 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-310
transform 1 0 3459 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-311
transform 1 0 3356 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-312
transform 1 0 3291 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-313
transform 1 0 3586 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-314
transform 1 0 3535 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-315
transform 1 0 3375 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-316
transform 1 0 3525 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-317
transform 1 0 3455 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-318
transform 1 0 3354 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-319
transform 1 0 3149 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-320
transform 1 0 3132 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-321
transform 1 0 3140 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-322
transform 1 0 2893 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-323
transform 1 0 3218 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-324
transform 1 0 2955 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-325
transform 1 0 2965 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-326
transform 1 0 2962 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-327
transform 1 0 3182 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-328
transform 1 0 3198 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-329
transform 1 0 3206 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-330
transform 1 0 3267 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-331
transform 1 0 3315 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-332
transform 1 0 3308 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-333
transform 1 0 3306 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-334
transform 1 0 3290 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-335
transform 1 0 3317 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-336
transform 1 0 3301 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-337
transform 1 0 3390 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-338
transform 1 0 3399 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-339
transform 1 0 3375 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-340
transform 1 0 3290 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-341
transform 1 0 3380 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-342
transform 1 0 3317 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-343
transform 1 0 3333 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-344
transform 1 0 3292 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-345
transform 1 0 3124 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-346
transform 1 0 3095 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-347
transform 1 0 3110 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-348
transform 1 0 3041 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-349
transform 1 0 3705 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-350
transform 1 0 3690 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-351
transform 1 0 3683 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-352
transform 1 0 3692 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-353
transform 1 0 3620 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-354
transform 1 0 3588 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-355
transform 1 0 3598 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-356
transform 1 0 3528 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-357
transform 1 0 3655 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-358
transform 1 0 3449 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-359
transform 1 0 3687 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-360
transform 1 0 3686 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-361
transform 1 0 3695 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-362
transform 1 0 3623 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-363
transform 1 0 3591 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-364
transform 1 0 3601 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-365
transform 1 0 3461 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-366
transform 1 0 3632 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-367
transform 1 0 3647 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-368
transform 1 0 3652 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-369
transform 1 0 3694 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-370
transform 1 0 3737 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-371
transform 1 0 3761 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-372
transform 1 0 3862 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-373
transform 1 0 3795 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-374
transform 1 0 3843 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-375
transform 1 0 3551 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-376
transform 1 0 3635 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-377
transform 1 0 3650 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-378
transform 1 0 3460 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-379
transform 1 0 3327 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-380
transform 1 0 3745 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-381
transform 1 0 3752 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-382
transform 1 0 3748 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-383
transform 1 0 3731 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-384
transform 1 0 3751 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-385
transform 1 0 3864 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-386
transform 1 0 3736 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-387
transform 1 0 3674 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-388
transform 1 0 3695 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-389
transform 1 0 3753 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-390
transform 1 0 3757 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-391
transform 1 0 3748 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-392
transform 1 0 3701 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-393
transform 1 0 3713 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-394
transform 1 0 3280 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-395
transform 1 0 3725 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-396
transform 1 0 3733 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-397
transform 1 0 3765 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-398
transform 1 0 3867 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-399
transform 1 0 3739 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-400
transform 1 0 3719 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-401
transform 1 0 3727 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-402
transform 1 0 3768 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-403
transform 1 0 3792 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-404
transform 1 0 3706 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-405
transform 1 0 3677 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-406
transform 1 0 3713 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-407
transform 1 0 3730 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-408
transform 1 0 3638 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-409
transform 1 0 3605 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-410
transform 1 0 3614 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-411
transform 1 0 3531 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-412
transform 1 0 3421 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-413
transform 1 0 3294 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-414
transform 1 0 3682 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-415
transform 1 0 3665 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-416
transform 1 0 3673 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-417
transform 1 0 3434 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-418
transform 1 0 3654 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-419
transform 1 0 3366 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-420
transform 1 0 3505 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-421
transform 1 0 3586 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-422
transform 1 0 3688 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-423
transform 1 0 3669 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-424
transform 1 0 3696 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-425
transform 1 0 3792 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-426
transform 1 0 3767 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-427
transform 1 0 3369 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-428
transform 1 0 3508 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-429
transform 1 0 3589 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-430
transform 1 0 3691 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-431
transform 1 0 3672 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-432
transform 1 0 3699 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-433
transform 1 0 3795 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-434
transform 1 0 3770 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-435
transform 1 0 3493 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-436
transform 1 0 3574 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-437
transform 1 0 3676 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-438
transform 1 0 3657 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-439
transform 1 0 3684 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-440
transform 1 0 3780 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-441
transform 1 0 3755 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-442
transform 1 0 3771 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-443
transform 1 0 3810 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-444
transform 1 0 3925 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-445
transform 1 0 3780 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-446
transform 1 0 3041 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-447
transform 1 0 3020 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-448
transform 1 0 3047 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-449
transform 1 0 3106 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-450
transform 1 0 3089 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-451
transform 1 0 3092 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-452
transform 1 0 3087 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-453
transform 1 0 3074 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-454
transform 1 0 3032 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-455
transform 1 0 3047 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-456
transform 1 0 3048 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-457
transform 1 0 3033 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-458
transform 1 0 3018 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-459
transform 1 0 3016 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-460
transform 1 0 3078 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-461
transform 1 0 3064 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-462
transform 1 0 3069 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-463
transform 1 0 3272 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-464
transform 1 0 3318 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-465
transform 1 0 3314 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-466
transform 1 0 3079 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-467
transform 1 0 3135 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-468
transform 1 0 3164 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-469
transform 1 0 3122 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-470
transform 1 0 3108 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-471
transform 1 0 3149 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-472
transform 1 0 3383 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-473
transform 1 0 3402 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-474
transform 1 0 3492 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-475
transform 1 0 3599 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-476
transform 1 0 3608 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-477
transform 1 0 3344 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-478
transform 1 0 3102 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-479
transform 1 0 3344 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-480
transform 1 0 3099 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-481
transform 1 0 3191 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-482
transform 1 0 3462 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-483
transform 1 0 3399 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-484
transform 1 0 3161 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-485
transform 1 0 3370 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-486
transform 1 0 3453 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-487
transform 1 0 3482 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-488
transform 1 0 3304 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-489
transform 1 0 3187 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-490
transform 1 0 3150 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-491
transform 1 0 3173 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-492
transform 1 0 3428 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-493
transform 1 0 3366 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-494
transform 1 0 3399 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-495
transform 1 0 3347 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-496
transform 1 0 3186 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-497
transform 1 0 3330 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-498
transform 1 0 3035 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-499
transform 1 0 3265 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-500
transform 1 0 3182 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-501
transform 1 0 3213 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-502
transform 1 0 3278 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-503
transform 1 0 3276 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-504
transform 1 0 3266 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-505
transform 1 0 3232 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-506
transform 1 0 3221 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-507
transform 1 0 3248 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-508
transform 1 0 3218 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-509
transform 1 0 3174 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-510
transform 1 0 3142 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-511
transform 1 0 3040 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-512
transform 1 0 3629 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-513
transform 1 0 3655 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-514
transform 1 0 3554 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-515
transform 1 0 3545 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-516
transform 1 0 3425 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-517
transform 1 0 3240 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-518
transform 1 0 3412 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-519
transform 1 0 3661 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-520
transform 1 0 3041 0 1 8734
box 0 0 3 6
use FEEDTHRU  F-521
transform 1 0 3118 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-522
transform 1 0 3188 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-523
transform 1 0 3044 0 1 8734
box 0 0 3 6
use FEEDTHRU  F-524
transform 1 0 3079 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-525
transform 1 0 3029 0 1 8734
box 0 0 3 6
use FEEDTHRU  F-526
transform 1 0 3314 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-527
transform 1 0 3356 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-528
transform 1 0 3452 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-529
transform 1 0 3678 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-530
transform 1 0 3774 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-531
transform 1 0 3681 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-532
transform 1 0 3027 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-533
transform 1 0 3054 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-534
transform 1 0 3059 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-535
transform 1 0 3050 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-536
transform 1 0 3059 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-537
transform 1 0 3063 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-538
transform 1 0 3228 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-539
transform 1 0 3522 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-540
transform 1 0 3452 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-541
transform 1 0 3342 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-542
transform 1 0 3507 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-543
transform 1 0 3437 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-544
transform 1 0 3345 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-545
transform 1 0 3128 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-546
transform 1 0 3501 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-547
transform 1 0 3431 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-548
transform 1 0 3330 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-549
transform 1 0 3725 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-550
transform 1 0 3731 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-551
transform 1 0 3696 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-552
transform 1 0 3674 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-553
transform 1 0 3728 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-554
transform 1 0 3766 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-555
transform 1 0 3787 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-556
transform 1 0 3786 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-557
transform 1 0 3737 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-558
transform 1 0 3734 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-559
transform 1 0 3699 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-560
transform 1 0 3363 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-561
transform 1 0 3363 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-562
transform 1 0 3083 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-563
transform 1 0 3005 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-564
transform 1 0 3028 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-565
transform 1 0 3075 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-566
transform 1 0 3120 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-567
transform 1 0 3099 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-568
transform 1 0 3079 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-569
transform 1 0 3274 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-570
transform 1 0 3342 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-571
transform 1 0 3368 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-572
transform 1 0 3467 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-573
transform 1 0 3527 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-574
transform 1 0 3616 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-575
transform 1 0 3429 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-576
transform 1 0 3294 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-577
transform 1 0 3307 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-578
transform 1 0 3278 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-579
transform 1 0 3338 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-580
transform 1 0 3077 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-581
transform 1 0 3913 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-582
transform 1 0 3768 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-583
transform 1 0 3752 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-584
transform 1 0 3868 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-585
transform 1 0 3915 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-586
transform 1 0 3900 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-587
transform 1 0 3201 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-588
transform 1 0 3420 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-589
transform 1 0 3102 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-590
transform 1 0 3539 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-591
transform 1 0 3348 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-592
transform 1 0 3120 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-593
transform 1 0 3281 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-594
transform 1 0 3177 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-595
transform 1 0 3437 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-596
transform 1 0 3460 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-597
transform 1 0 3901 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-598
transform 1 0 3904 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-599
transform 1 0 3359 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-600
transform 1 0 3343 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-601
transform 1 0 3095 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-602
transform 1 0 3714 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-603
transform 1 0 3696 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-604
transform 1 0 3663 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-605
transform 1 0 3619 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-606
transform 1 0 3602 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-607
transform 1 0 3570 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-608
transform 1 0 3500 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-609
transform 1 0 3749 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-610
transform 1 0 3762 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-611
transform 1 0 3755 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-612
transform 1 0 3734 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-613
transform 1 0 3784 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-614
transform 1 0 3873 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-615
transform 1 0 3820 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-616
transform 1 0 3764 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-617
transform 1 0 3876 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-618
transform 1 0 3823 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-619
transform 1 0 3578 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-620
transform 1 0 3599 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-621
transform 1 0 3712 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-622
transform 1 0 3689 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-623
transform 1 0 3715 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-624
transform 1 0 3759 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-625
transform 1 0 3858 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-626
transform 1 0 2993 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-627
transform 1 0 3264 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-628
transform 1 0 3282 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-629
transform 1 0 3158 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-630
transform 1 0 3212 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-631
transform 1 0 3236 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-632
transform 1 0 2990 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-633
transform 1 0 3011 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-634
transform 1 0 3563 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-635
transform 1 0 3536 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-636
transform 1 0 3566 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-637
transform 1 0 3883 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-638
transform 1 0 3313 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-639
transform 1 0 3233 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-640
transform 1 0 3135 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-641
transform 1 0 2985 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-642
transform 1 0 3034 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-643
transform 1 0 2988 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-644
transform 1 0 2965 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-645
transform 1 0 3039 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-646
transform 1 0 3003 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-647
transform 1 0 3357 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-648
transform 1 0 2947 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-649
transform 1 0 2952 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-650
transform 1 0 2997 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-651
transform 1 0 2971 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-652
transform 1 0 2978 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-653
transform 1 0 3849 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-654
transform 1 0 3846 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-655
transform 1 0 3796 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-656
transform 1 0 3746 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-657
transform 1 0 3474 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-658
transform 1 0 3541 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-659
transform 1 0 3444 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-660
transform 1 0 3143 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-661
transform 1 0 3167 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-662
transform 1 0 3125 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-663
transform 1 0 3132 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-664
transform 1 0 3076 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-665
transform 1 0 3016 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-666
transform 1 0 3040 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-667
transform 1 0 3029 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-668
transform 1 0 3064 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-669
transform 1 0 3086 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-670
transform 1 0 3035 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-671
transform 1 0 3225 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-672
transform 1 0 3536 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-673
transform 1 0 3198 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-674
transform 1 0 3501 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-675
transform 1 0 3000 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-676
transform 1 0 3013 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-677
transform 1 0 3072 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-678
transform 1 0 2963 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-679
transform 1 0 3798 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-680
transform 1 0 3846 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-681
transform 1 0 3849 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-682
transform 1 0 3762 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-683
transform 1 0 3861 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-684
transform 1 0 3712 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-685
transform 1 0 3683 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-686
transform 1 0 3740 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-687
transform 1 0 3789 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-688
transform 1 0 3840 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-689
transform 1 0 3747 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-690
transform 1 0 3718 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-691
transform 1 0 3692 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-692
transform 1 0 3715 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-693
transform 1 0 3602 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-694
transform 1 0 3581 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-695
transform 1 0 3661 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-696
transform 1 0 3519 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-697
transform 1 0 3463 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-698
transform 1 0 3330 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-699
transform 1 0 3655 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-700
transform 1 0 3005 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-701
transform 1 0 3002 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-702
transform 1 0 3052 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-703
transform 1 0 3582 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-704
transform 1 0 3608 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-705
transform 1 0 3665 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-706
transform 1 0 3647 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-707
transform 1 0 3515 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-708
transform 1 0 3432 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-709
transform 1 0 3659 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-710
transform 1 0 3531 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-711
transform 1 0 3708 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-712
transform 1 0 3531 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-713
transform 1 0 3658 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-714
transform 1 0 3362 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-715
transform 1 0 3621 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-716
transform 1 0 3780 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-717
transform 1 0 3653 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-718
transform 1 0 3495 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-719
transform 1 0 3402 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-720
transform 1 0 3321 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-721
transform 1 0 3598 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-722
transform 1 0 3326 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-723
transform 1 0 3624 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-724
transform 1 0 3387 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-725
transform 1 0 3698 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-726
transform 1 0 3685 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-727
transform 1 0 3545 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-728
transform 1 0 3539 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-729
transform 1 0 3676 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-730
transform 1 0 3692 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-731
transform 1 0 3741 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-732
transform 1 0 3630 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-733
transform 1 0 3467 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-734
transform 1 0 3756 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-735
transform 1 0 3714 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-736
transform 1 0 3043 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-737
transform 1 0 3110 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-738
transform 1 0 3276 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-739
transform 1 0 3377 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-740
transform 1 0 3453 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-741
transform 1 0 3168 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-742
transform 1 0 3529 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-743
transform 1 0 3565 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-744
transform 1 0 3198 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-745
transform 1 0 3215 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-746
transform 1 0 3512 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-747
transform 1 0 3566 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-748
transform 1 0 3207 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-749
transform 1 0 3243 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-750
transform 1 0 3222 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-751
transform 1 0 3457 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-752
transform 1 0 3197 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-753
transform 1 0 3567 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-754
transform 1 0 3204 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-755
transform 1 0 3641 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-756
transform 1 0 3366 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-757
transform 1 0 3596 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-758
transform 1 0 3601 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-759
transform 1 0 3332 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-760
transform 1 0 3341 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-761
transform 1 0 3359 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-762
transform 1 0 3407 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-763
transform 1 0 3357 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-764
transform 1 0 3289 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-765
transform 1 0 3173 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-766
transform 1 0 3378 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-767
transform 1 0 3528 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-768
transform 1 0 3458 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-769
transform 1 0 3264 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-770
transform 1 0 3538 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-771
transform 1 0 3589 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-772
transform 1 0 3237 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-773
transform 1 0 3324 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-774
transform 1 0 3478 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-775
transform 1 0 3514 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-776
transform 1 0 3228 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-777
transform 1 0 3221 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-778
transform 1 0 3632 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-779
transform 1 0 3002 0 1 8734
box 0 0 3 6
use FEEDTHRU  F-780
transform 1 0 3928 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-781
transform 1 0 3783 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-782
transform 1 0 3701 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-783
transform 1 0 3758 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-784
transform 1 0 3921 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-785
transform 1 0 3906 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-786
transform 1 0 3904 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-787
transform 1 0 3850 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-788
transform 1 0 3724 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-789
transform 1 0 3704 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-790
transform 1 0 3761 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-791
transform 1 0 3792 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-792
transform 1 0 3760 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-793
transform 1 0 3775 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-794
transform 1 0 3759 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-795
transform 1 0 3713 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-796
transform 1 0 3656 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-797
transform 1 0 3691 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-798
transform 1 0 3822 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-799
transform 1 0 3735 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-800
transform 1 0 3703 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-801
transform 1 0 3701 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-802
transform 1 0 3588 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-803
transform 1 0 3602 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-804
transform 1 0 3528 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-805
transform 1 0 3579 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-806
transform 1 0 3591 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-807
transform 1 0 3587 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-808
transform 1 0 3586 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-809
transform 1 0 3371 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-810
transform 1 0 3387 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-811
transform 1 0 3366 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-812
transform 1 0 3501 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-813
transform 1 0 3829 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-814
transform 1 0 3718 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-815
transform 1 0 3623 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-816
transform 1 0 3599 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-817
transform 1 0 3623 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-818
transform 1 0 3831 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-819
transform 1 0 3852 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-820
transform 1 0 3828 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-821
transform 1 0 3700 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-822
transform 1 0 3201 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-823
transform 1 0 2963 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-824
transform 1 0 3232 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-825
transform 1 0 3300 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-826
transform 1 0 3293 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-827
transform 1 0 3242 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-828
transform 1 0 3188 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-829
transform 1 0 3144 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-830
transform 1 0 2983 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-831
transform 1 0 2960 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-832
transform 1 0 2985 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-833
transform 1 0 3017 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-834
transform 1 0 3022 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-835
transform 1 0 3013 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-836
transform 1 0 3007 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-837
transform 1 0 3697 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-838
transform 1 0 3726 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-839
transform 1 0 3804 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-840
transform 1 0 3685 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-841
transform 1 0 3668 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-842
transform 1 0 3725 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-843
transform 1 0 3765 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-844
transform 1 0 3781 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-845
transform 1 0 3729 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-846
transform 1 0 3798 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-847
transform 1 0 3688 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-848
transform 1 0 3671 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-849
transform 1 0 3728 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-850
transform 1 0 3700 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-851
transform 1 0 3695 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-852
transform 1 0 3706 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-853
transform 1 0 3287 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-854
transform 1 0 2999 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-855
transform 1 0 3003 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-856
transform 1 0 3804 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-857
transform 1 0 3620 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-858
transform 1 0 3610 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-859
transform 1 0 3656 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-860
transform 1 0 3453 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-861
transform 1 0 2956 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-862
transform 1 0 2932 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-863
transform 1 0 3149 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-864
transform 1 0 3226 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-865
transform 1 0 3512 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-866
transform 1 0 3727 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-867
transform 1 0 3599 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-868
transform 1 0 3594 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-869
transform 1 0 3632 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-870
transform 1 0 3450 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-871
transform 1 0 3657 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-872
transform 1 0 3437 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-873
transform 1 0 3575 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-874
transform 1 0 3572 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-875
transform 1 0 3480 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-876
transform 1 0 3451 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-877
transform 1 0 3196 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-878
transform 1 0 3181 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-879
transform 1 0 3183 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-880
transform 1 0 3162 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-881
transform 1 0 3140 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-882
transform 1 0 3093 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-883
transform 1 0 3732 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-884
transform 1 0 3816 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-885
transform 1 0 3819 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-886
transform 1 0 3697 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-887
transform 1 0 3680 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-888
transform 1 0 3743 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-889
transform 1 0 3470 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-890
transform 1 0 3465 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-891
transform 1 0 3376 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-892
transform 1 0 3310 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-893
transform 1 0 3167 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-894
transform 1 0 3161 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-895
transform 1 0 3173 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-896
transform 1 0 3365 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-897
transform 1 0 3138 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-898
transform 1 0 3137 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-899
transform 1 0 3105 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-900
transform 1 0 3013 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-901
transform 1 0 3611 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-902
transform 1 0 3601 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-903
transform 1 0 3651 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-904
transform 1 0 3680 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-905
transform 1 0 3702 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-906
transform 1 0 3737 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-907
transform 1 0 3719 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-908
transform 1 0 3775 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-909
transform 1 0 3590 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-910
transform 1 0 3604 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-911
transform 1 0 3654 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-912
transform 1 0 3811 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-913
transform 1 0 3858 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-914
transform 1 0 3855 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-915
transform 1 0 3736 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-916
transform 1 0 3786 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-917
transform 1 0 3792 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-918
transform 1 0 3739 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-919
transform 1 0 3714 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-920
transform 1 0 3678 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-921
transform 1 0 3616 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-922
transform 1 0 3557 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-923
transform 1 0 3537 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-924
transform 1 0 3467 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-925
transform 1 0 3773 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-926
transform 1 0 3795 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-927
transform 1 0 3940 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-928
transform 1 0 3807 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-929
transform 1 0 3123 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-930
transform 1 0 3170 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-931
transform 1 0 3033 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-932
transform 1 0 3055 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-933
transform 1 0 3057 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-934
transform 1 0 3077 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-935
transform 1 0 3113 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-936
transform 1 0 3052 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-937
transform 1 0 3084 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-938
transform 1 0 3069 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-939
transform 1 0 3060 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-940
transform 1 0 3063 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-941
transform 1 0 3012 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-942
transform 1 0 3058 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-943
transform 1 0 3090 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-944
transform 1 0 3075 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-945
transform 1 0 3066 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-946
transform 1 0 3084 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-947
transform 1 0 3090 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-948
transform 1 0 3110 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-949
transform 1 0 3128 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-950
transform 1 0 3224 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-951
transform 1 0 3017 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-952
transform 1 0 3143 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-953
transform 1 0 3114 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-954
transform 1 0 3126 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-955
transform 1 0 3091 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-956
transform 1 0 3155 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-957
transform 1 0 3113 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-958
transform 1 0 3117 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-959
transform 1 0 3116 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-960
transform 1 0 3119 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-961
transform 1 0 3133 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-962
transform 1 0 3101 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-963
transform 1 0 3176 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-964
transform 1 0 3258 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-965
transform 1 0 3328 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-966
transform 1 0 3265 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-967
transform 1 0 3286 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-968
transform 1 0 3255 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-969
transform 1 0 3429 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-970
transform 1 0 3353 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-971
transform 1 0 3350 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-972
transform 1 0 3141 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-973
transform 1 0 3317 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-974
transform 1 0 3402 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-975
transform 1 0 3186 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-976
transform 1 0 3271 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-977
transform 1 0 3211 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-978
transform 1 0 3720 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-979
transform 1 0 3671 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-980
transform 1 0 3686 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-981
transform 1 0 3581 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-982
transform 1 0 3531 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-983
transform 1 0 3568 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-984
transform 1 0 3717 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-985
transform 1 0 3717 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-986
transform 1 0 3702 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-987
transform 1 0 3661 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-988
transform 1 0 3479 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-989
transform 1 0 3045 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-990
transform 1 0 3040 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-991
transform 1 0 3042 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-992
transform 1 0 3053 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-993
transform 1 0 3030 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-994
transform 1 0 3244 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-995
transform 1 0 3072 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-996
transform 1 0 3025 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-997
transform 1 0 3054 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-998
transform 1 0 3037 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-999
transform 1 0 3318 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1000
transform 1 0 3310 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1001
transform 1 0 3390 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1002
transform 1 0 3701 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1003
transform 1 0 3641 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1004
transform 1 0 3784 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1005
transform 1 0 2982 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1006
transform 1 0 3031 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1007
transform 1 0 3048 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1008
transform 1 0 3035 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1009
transform 1 0 3677 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1010
transform 1 0 3583 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1011
transform 1 0 3716 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1012
transform 1 0 3388 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1013
transform 1 0 3248 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1014
transform 1 0 3396 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1015
transform 1 0 3186 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1016
transform 1 0 3519 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1017
transform 1 0 3537 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1018
transform 1 0 3198 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1019
transform 1 0 3322 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1020
transform 1 0 3195 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1021
transform 1 0 3152 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-1022
transform 1 0 3357 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1023
transform 1 0 3246 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1024
transform 1 0 3753 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1025
transform 1 0 3686 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1026
transform 1 0 3646 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1027
transform 1 0 3796 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1028
transform 1 0 3801 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1029
transform 1 0 3629 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1030
transform 1 0 3132 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1031
transform 1 0 3138 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1032
transform 1 0 3199 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1033
transform 1 0 3234 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1034
transform 1 0 3331 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1035
transform 1 0 3289 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1036
transform 1 0 3403 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1037
transform 1 0 3261 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1038
transform 1 0 3239 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1039
transform 1 0 3533 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1040
transform 1 0 3590 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1041
transform 1 0 3500 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1042
transform 1 0 3401 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1043
transform 1 0 3345 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1044
transform 1 0 3440 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1045
transform 1 0 3463 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1046
transform 1 0 3395 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1047
transform 1 0 3629 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1048
transform 1 0 3008 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1049
transform 1 0 3008 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1050
transform 1 0 3498 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1051
transform 1 0 3249 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1052
transform 1 0 3062 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1053
transform 1 0 3071 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1054
transform 1 0 3068 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1055
transform 1 0 3074 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1056
transform 1 0 3532 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1057
transform 1 0 3290 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1058
transform 1 0 3305 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1059
transform 1 0 3290 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1060
transform 1 0 3359 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1061
transform 1 0 3303 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1062
transform 1 0 3162 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1063
transform 1 0 3186 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1064
transform 1 0 3037 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1065
transform 1 0 3257 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1066
transform 1 0 3021 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1067
transform 1 0 3032 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1068
transform 1 0 3057 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1069
transform 1 0 3028 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1070
transform 1 0 3069 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1071
transform 1 0 3047 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1072
transform 1 0 3065 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1073
transform 1 0 3079 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1074
transform 1 0 3077 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1075
transform 1 0 3074 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1076
transform 1 0 3069 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1077
transform 1 0 3065 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1078
transform 1 0 3113 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1079
transform 1 0 3098 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1080
transform 1 0 3096 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1081
transform 1 0 3078 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1082
transform 1 0 3042 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1083
transform 1 0 3050 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1084
transform 1 0 3060 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1085
transform 1 0 3034 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1086
transform 1 0 3062 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1087
transform 1 0 3044 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1088
transform 1 0 3047 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1089
transform 1 0 3095 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1090
transform 1 0 3047 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1091
transform 1 0 3057 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1092
transform 1 0 3084 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1093
transform 1 0 3057 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1094
transform 1 0 3083 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1095
transform 1 0 3101 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1096
transform 1 0 3226 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1097
transform 1 0 3260 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1098
transform 1 0 3095 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1099
transform 1 0 3110 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1100
transform 1 0 3104 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1101
transform 1 0 3105 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1102
transform 1 0 3303 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1103
transform 1 0 3436 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1104
transform 1 0 3513 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1105
transform 1 0 3228 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1106
transform 1 0 3125 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-1107
transform 1 0 3046 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-1108
transform 1 0 3036 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1109
transform 1 0 3069 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1110
transform 1 0 3617 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1111
transform 1 0 3593 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1112
transform 1 0 3617 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1113
transform 1 0 3694 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1114
transform 1 0 3677 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1115
transform 1 0 3774 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1116
transform 1 0 3438 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1117
transform 1 0 3495 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1118
transform 1 0 3419 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1119
transform 1 0 3318 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1120
transform 1 0 3454 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1121
transform 1 0 3502 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1122
transform 1 0 3495 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1123
transform 1 0 3506 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1124
transform 1 0 3641 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1125
transform 1 0 3647 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1126
transform 1 0 3044 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1127
transform 1 0 3045 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1128
transform 1 0 3116 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1129
transform 1 0 3449 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1130
transform 1 0 3522 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1131
transform 1 0 3189 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1132
transform 1 0 3165 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1133
transform 1 0 3425 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1134
transform 1 0 3275 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1135
transform 1 0 3197 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1136
transform 1 0 3216 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1137
transform 1 0 3253 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1138
transform 1 0 3050 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1139
transform 1 0 3053 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1140
transform 1 0 3046 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1141
transform 1 0 3698 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1142
transform 1 0 3459 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1143
transform 1 0 3760 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1144
transform 1 0 3751 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1145
transform 1 0 3704 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1146
transform 1 0 3716 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1147
transform 1 0 3610 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1148
transform 1 0 3380 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1149
transform 1 0 3579 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1150
transform 1 0 3576 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1151
transform 1 0 3555 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1152
transform 1 0 3592 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1153
transform 1 0 3644 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1154
transform 1 0 3437 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1155
transform 1 0 3360 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1156
transform 1 0 3650 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1157
transform 1 0 3584 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1158
transform 1 0 3417 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1159
transform 1 0 3578 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1160
transform 1 0 3371 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1161
transform 1 0 3516 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1162
transform 1 0 3587 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1163
transform 1 0 3560 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1164
transform 1 0 3663 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1165
transform 1 0 3646 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1166
transform 1 0 3638 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1167
transform 1 0 3634 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1168
transform 1 0 3650 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1169
transform 1 0 3747 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1170
transform 1 0 3642 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1171
transform 1 0 3611 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1172
transform 1 0 3501 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1173
transform 1 0 3439 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1174
transform 1 0 3306 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1175
transform 1 0 3315 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1176
transform 1 0 3234 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1177
transform 1 0 3111 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1178
transform 1 0 3015 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1179
transform 1 0 3030 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1180
transform 1 0 3020 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1181
transform 1 0 3498 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1182
transform 1 0 3422 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1183
transform 1 0 3321 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1184
transform 1 0 3383 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1185
transform 1 0 3282 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1186
transform 1 0 3155 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-1187
transform 1 0 3323 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1188
transform 1 0 3206 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1189
transform 1 0 3086 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1190
transform 1 0 3240 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1191
transform 1 0 3459 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1192
transform 1 0 3444 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1193
transform 1 0 3313 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1194
transform 1 0 3242 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1195
transform 1 0 3153 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1196
transform 1 0 3420 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1197
transform 1 0 3260 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1198
transform 1 0 3240 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1199
transform 1 0 3208 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1200
transform 1 0 3101 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1201
transform 1 0 3119 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1202
transform 1 0 3129 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1203
transform 1 0 3125 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1204
transform 1 0 3106 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1205
transform 1 0 3126 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1206
transform 1 0 3235 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1207
transform 1 0 3252 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1208
transform 1 0 3297 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1209
transform 1 0 3230 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1210
transform 1 0 3249 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1211
transform 1 0 3530 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1212
transform 1 0 3494 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1213
transform 1 0 3260 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1214
transform 1 0 3209 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1215
transform 1 0 3212 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1216
transform 1 0 3235 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1217
transform 1 0 3276 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1218
transform 1 0 3296 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1219
transform 1 0 3428 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1220
transform 1 0 3422 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1221
transform 1 0 3535 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1222
transform 1 0 3575 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1223
transform 1 0 3582 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1224
transform 1 0 3530 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1225
transform 1 0 3300 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1226
transform 1 0 3247 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1227
transform 1 0 3288 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1228
transform 1 0 3320 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1229
transform 1 0 3636 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1230
transform 1 0 3745 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1231
transform 1 0 3668 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1232
transform 1 0 3626 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1233
transform 1 0 3536 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1234
transform 1 0 3637 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1235
transform 1 0 3696 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1236
transform 1 0 3711 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1237
transform 1 0 3693 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1238
transform 1 0 3009 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1239
transform 1 0 2976 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1240
transform 1 0 2932 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1241
transform 1 0 2973 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1242
transform 1 0 3496 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1243
transform 1 0 3495 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1244
transform 1 0 3483 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1245
transform 1 0 3401 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1246
transform 1 0 3309 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1247
transform 1 0 3173 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-1248
transform 1 0 3499 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1249
transform 1 0 3498 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1250
transform 1 0 3486 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1251
transform 1 0 3404 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1252
transform 1 0 3312 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1253
transform 1 0 3176 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-1254
transform 1 0 3546 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1255
transform 1 0 3510 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1256
transform 1 0 3218 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1257
transform 1 0 3372 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1258
transform 1 0 3035 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1259
transform 1 0 3059 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1260
transform 1 0 3064 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1261
transform 1 0 3360 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1262
transform 1 0 3080 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1263
transform 1 0 3075 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1264
transform 1 0 3053 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1265
transform 1 0 3186 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1266
transform 1 0 3157 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1267
transform 1 0 3211 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1268
transform 1 0 3162 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1269
transform 1 0 3043 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-1270
transform 1 0 3088 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1271
transform 1 0 3172 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1272
transform 1 0 3355 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1273
transform 1 0 3480 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1274
transform 1 0 3590 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1275
transform 1 0 3399 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1276
transform 1 0 3473 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1277
transform 1 0 3320 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1278
transform 1 0 3422 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1279
transform 1 0 3392 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1280
transform 1 0 3393 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1281
transform 1 0 3322 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1282
transform 1 0 3444 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1283
transform 1 0 3441 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1284
transform 1 0 3432 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1285
transform 1 0 3169 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1286
transform 1 0 3155 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1287
transform 1 0 3309 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1288
transform 1 0 3348 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1289
transform 1 0 3179 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1290
transform 1 0 3183 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1291
transform 1 0 3177 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1292
transform 1 0 3189 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1293
transform 1 0 3196 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1294
transform 1 0 3167 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1295
transform 1 0 3144 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1296
transform 1 0 3156 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1297
transform 1 0 3201 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1298
transform 1 0 3356 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1299
transform 1 0 3432 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1300
transform 1 0 3533 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1301
transform 1 0 3524 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1302
transform 1 0 3551 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1303
transform 1 0 3432 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1304
transform 1 0 3358 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1305
transform 1 0 3254 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1306
transform 1 0 3486 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1307
transform 1 0 3125 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1308
transform 1 0 3185 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1309
transform 1 0 3179 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1310
transform 1 0 3441 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1311
transform 1 0 3131 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1312
transform 1 0 3191 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1313
transform 1 0 3185 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1314
transform 1 0 3180 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1315
transform 1 0 3163 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1316
transform 1 0 3103 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1317
transform 1 0 3162 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1318
transform 1 0 3159 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1319
transform 1 0 3051 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1320
transform 1 0 3117 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1321
transform 1 0 3129 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1322
transform 1 0 3137 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1323
transform 1 0 3140 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1324
transform 1 0 3080 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1325
transform 1 0 3105 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1326
transform 1 0 3104 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1327
transform 1 0 3107 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1328
transform 1 0 3082 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1329
transform 1 0 3077 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1330
transform 1 0 3053 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1331
transform 1 0 3081 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1332
transform 1 0 3040 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1333
transform 1 0 3210 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1334
transform 1 0 3194 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1335
transform 1 0 3181 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1336
transform 1 0 3173 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1337
transform 1 0 3188 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1338
transform 1 0 3212 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1339
transform 1 0 3090 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1340
transform 1 0 3083 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1341
transform 1 0 3193 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1342
transform 1 0 3079 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1343
transform 1 0 3605 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1344
transform 1 0 3688 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1345
transform 1 0 3662 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1346
transform 1 0 3670 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1347
transform 1 0 3108 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1348
transform 1 0 3105 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1349
transform 1 0 3120 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1350
transform 1 0 3128 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1351
transform 1 0 3664 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1352
transform 1 0 3644 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1353
transform 1 0 3652 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1354
transform 1 0 3813 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1355
transform 1 0 3771 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1356
transform 1 0 3643 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1357
transform 1 0 3723 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1358
transform 1 0 3705 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1359
transform 1 0 3614 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1360
transform 1 0 3659 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1361
transform 1 0 3644 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1362
transform 1 0 3639 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1363
transform 1 0 3577 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1364
transform 1 0 3520 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1365
transform 1 0 3531 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1366
transform 1 0 3489 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1367
transform 1 0 3407 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1368
transform 1 0 3324 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1369
transform 1 0 3080 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1370
transform 1 0 3058 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1371
transform 1 0 3047 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1372
transform 1 0 3176 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1373
transform 1 0 3200 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1374
transform 1 0 3212 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1375
transform 1 0 3129 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1376
transform 1 0 3149 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1377
transform 1 0 3246 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1378
transform 1 0 3552 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1379
transform 1 0 3576 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1380
transform 1 0 3572 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1381
transform 1 0 3611 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1382
transform 1 0 3419 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1383
transform 1 0 3408 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1384
transform 1 0 3662 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1385
transform 1 0 3640 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1386
transform 1 0 3632 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1387
transform 1 0 3765 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1388
transform 1 0 3660 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1389
transform 1 0 3216 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1390
transform 1 0 3370 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1391
transform 1 0 3221 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1392
transform 1 0 3222 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1393
transform 1 0 3318 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1394
transform 1 0 3245 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1395
transform 1 0 3379 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1396
transform 1 0 3246 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1397
transform 1 0 3315 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1398
transform 1 0 3255 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1399
transform 1 0 3086 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-1400
transform 1 0 3180 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1401
transform 1 0 3227 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1402
transform 1 0 3016 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-1403
transform 1 0 3489 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1404
transform 1 0 3531 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1405
transform 1 0 3510 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1406
transform 1 0 3413 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1407
transform 1 0 3503 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1408
transform 1 0 3245 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1409
transform 1 0 3255 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1410
transform 1 0 3325 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1411
transform 1 0 3309 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1412
transform 1 0 3397 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1413
transform 1 0 3431 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1414
transform 1 0 3423 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1415
transform 1 0 3267 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1416
transform 1 0 3740 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1417
transform 1 0 3764 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1418
transform 1 0 3680 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1419
transform 1 0 3632 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1420
transform 1 0 3742 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1421
transform 1 0 3312 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1422
transform 1 0 3302 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1423
transform 1 0 3310 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1424
transform 1 0 3074 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1425
transform 1 0 3101 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1426
transform 1 0 3083 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1427
transform 1 0 3096 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1428
transform 1 0 3244 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1429
transform 1 0 3403 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1430
transform 1 0 3296 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1431
transform 1 0 3501 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1432
transform 1 0 3288 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1433
transform 1 0 3479 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1434
transform 1 0 3363 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1435
transform 1 0 3389 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1436
transform 1 0 3424 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1437
transform 1 0 3363 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1438
transform 1 0 3432 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1439
transform 1 0 3465 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1440
transform 1 0 3419 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1441
transform 1 0 3498 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1442
transform 1 0 3556 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1443
transform 1 0 3508 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1444
transform 1 0 3160 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-1445
transform 1 0 3266 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1446
transform 1 0 3115 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1447
transform 1 0 3123 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1448
transform 1 0 3147 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1449
transform 1 0 3116 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1450
transform 1 0 3063 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1451
transform 1 0 3121 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1452
transform 1 0 3175 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1453
transform 1 0 3192 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1454
transform 1 0 3159 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1455
transform 1 0 3534 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1456
transform 1 0 3544 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1457
transform 1 0 3502 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1458
transform 1 0 3560 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1459
transform 1 0 3540 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1460
transform 1 0 3470 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1461
transform 1 0 3315 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1462
transform 1 0 3626 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1463
transform 1 0 3189 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1464
transform 1 0 3119 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1465
transform 1 0 3179 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1466
transform 1 0 3183 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1467
transform 1 0 3204 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1468
transform 1 0 3157 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1469
transform 1 0 3161 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1470
transform 1 0 3120 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1471
transform 1 0 3144 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1472
transform 1 0 3095 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1473
transform 1 0 3584 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1474
transform 1 0 3608 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1475
transform 1 0 3691 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1476
transform 1 0 3699 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1477
transform 1 0 3717 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1478
transform 1 0 3752 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1479
transform 1 0 3596 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1480
transform 1 0 3763 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1481
transform 1 0 3778 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1482
transform 1 0 3073 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1483
transform 1 0 3072 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1484
transform 1 0 3071 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1485
transform 1 0 3077 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1486
transform 1 0 3062 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1487
transform 1 0 3076 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1488
transform 1 0 2961 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-1489
transform 1 0 3544 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1490
transform 1 0 3447 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1491
transform 1 0 3414 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1492
transform 1 0 3335 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1493
transform 1 0 3252 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1494
transform 1 0 3242 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1495
transform 1 0 3323 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1496
transform 1 0 3339 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1497
transform 1 0 3347 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1498
transform 1 0 3234 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1499
transform 1 0 3384 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1500
transform 1 0 3762 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1501
transform 1 0 3542 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1502
transform 1 0 3623 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1503
transform 1 0 3560 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1504
transform 1 0 3630 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1505
transform 1 0 3478 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1506
transform 1 0 3448 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1507
transform 1 0 3417 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1508
transform 1 0 3177 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1509
transform 1 0 3131 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1510
transform 1 0 3121 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1511
transform 1 0 3180 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1512
transform 1 0 3128 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1513
transform 1 0 3118 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1514
transform 1 0 3177 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1515
transform 1 0 3156 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1516
transform 1 0 3156 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1517
transform 1 0 3423 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1518
transform 1 0 3416 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1519
transform 1 0 3500 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1520
transform 1 0 2964 0 1 8734
box 0 0 3 6
use FEEDTHRU  F-1521
transform 1 0 2989 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-1522
transform 1 0 3013 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1523
transform 1 0 3094 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1524
transform 1 0 3114 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1525
transform 1 0 3113 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1526
transform 1 0 3131 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1527
transform 1 0 3116 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1528
transform 1 0 3124 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1529
transform 1 0 3161 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1530
transform 1 0 3171 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1531
transform 1 0 3173 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1532
transform 1 0 3192 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1533
transform 1 0 3156 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1534
transform 1 0 3215 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1535
transform 1 0 3208 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1536
transform 1 0 3252 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1537
transform 1 0 3213 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1538
transform 1 0 3231 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1539
transform 1 0 3143 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1540
transform 1 0 3233 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1541
transform 1 0 3072 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1542
transform 1 0 3342 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1543
transform 1 0 3347 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1544
transform 1 0 3187 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1545
transform 1 0 3228 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1546
transform 1 0 3201 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1547
transform 1 0 3408 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1548
transform 1 0 3191 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1549
transform 1 0 3243 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1550
transform 1 0 3432 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1551
transform 1 0 3143 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1552
transform 1 0 3141 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1553
transform 1 0 3131 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1554
transform 1 0 3100 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1555
transform 1 0 3235 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1556
transform 1 0 3249 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1557
transform 1 0 3227 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1558
transform 1 0 3419 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1559
transform 1 0 3197 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1560
transform 1 0 3059 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1561
transform 1 0 3063 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1562
transform 1 0 3061 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1563
transform 1 0 3220 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1564
transform 1 0 3225 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1565
transform 1 0 2887 0 1 8734
box 0 0 3 6
use FEEDTHRU  F-1566
transform 1 0 3735 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1567
transform 1 0 3395 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1568
transform 1 0 3419 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1569
transform 1 0 3258 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1570
transform 1 0 3229 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1571
transform 1 0 3182 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1572
transform 1 0 2983 0 1 8734
box 0 0 3 6
use FEEDTHRU  F-1573
transform 1 0 3025 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-1574
transform 1 0 3055 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1575
transform 1 0 3118 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1576
transform 1 0 3204 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1577
transform 1 0 3236 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1578
transform 1 0 3242 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1579
transform 1 0 3317 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1580
transform 1 0 3322 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1581
transform 1 0 3616 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1582
transform 1 0 3602 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1583
transform 1 0 3622 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1584
transform 1 0 3451 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1585
transform 1 0 3102 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1586
transform 1 0 3101 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1587
transform 1 0 3107 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1588
transform 1 0 3092 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1589
transform 1 0 3582 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1590
transform 1 0 3415 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1591
transform 1 0 3423 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1592
transform 1 0 3507 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1593
transform 1 0 3317 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1594
transform 1 0 3321 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1595
transform 1 0 3279 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1596
transform 1 0 3273 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1597
transform 1 0 3413 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1598
transform 1 0 3299 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1599
transform 1 0 3285 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1600
transform 1 0 3305 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1601
transform 1 0 3227 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1602
transform 1 0 3261 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1603
transform 1 0 3255 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1604
transform 1 0 3049 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1605
transform 1 0 3066 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1606
transform 1 0 3155 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1607
transform 1 0 3668 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1608
transform 1 0 3665 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1609
transform 1 0 3631 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1610
transform 1 0 3768 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1611
transform 1 0 3199 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1612
transform 1 0 3169 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1613
transform 1 0 3204 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1614
transform 1 0 3493 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1615
transform 1 0 3392 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1616
transform 1 0 3407 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1617
transform 1 0 3290 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1618
transform 1 0 3453 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1619
transform 1 0 3524 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1620
transform 1 0 3375 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1621
transform 1 0 3468 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1622
transform 1 0 3423 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1623
transform 1 0 3084 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1624
transform 1 0 3089 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1625
transform 1 0 3089 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1626
transform 1 0 3090 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1627
transform 1 0 3095 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1628
transform 1 0 3095 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1629
transform 1 0 3080 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1630
transform 1 0 3222 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1631
transform 1 0 3209 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1632
transform 1 0 3245 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1633
transform 1 0 3167 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1634
transform 1 0 3243 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1635
transform 1 0 3237 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1636
transform 1 0 3193 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1637
transform 1 0 3127 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1638
transform 1 0 3150 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1639
transform 1 0 3149 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1640
transform 1 0 3225 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1641
transform 1 0 3219 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1642
transform 1 0 3234 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1643
transform 1 0 3720 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1644
transform 1 0 3267 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1645
transform 1 0 3193 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1646
transform 1 0 3152 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1647
transform 1 0 3183 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-1648
transform 1 0 3278 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1649
transform 1 0 3424 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1650
transform 1 0 3498 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1651
transform 1 0 3626 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1652
transform 1 0 3602 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1653
transform 1 0 3563 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1654
transform 1 0 3721 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1655
transform 1 0 3052 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1656
transform 1 0 3063 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1657
transform 1 0 3790 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1658
transform 1 0 3769 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1659
transform 1 0 3548 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1660
transform 1 0 3690 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1661
transform 1 0 3179 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1662
transform 1 0 3181 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1663
transform 1 0 3130 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1664
transform 1 0 3140 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1665
transform 1 0 3195 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1666
transform 1 0 3570 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1667
transform 1 0 3566 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1668
transform 1 0 3393 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1669
transform 1 0 3573 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1670
transform 1 0 3558 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1671
transform 1 0 3563 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1672
transform 1 0 3574 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1673
transform 1 0 3488 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1674
transform 1 0 3540 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1675
transform 1 0 3539 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1676
transform 1 0 3553 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1677
transform 1 0 3587 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1678
transform 1 0 3597 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1679
transform 1 0 3729 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1680
transform 1 0 3620 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1681
transform 1 0 3792 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1682
transform 1 0 3581 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1683
transform 1 0 3813 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1684
transform 1 0 3723 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1685
transform 1 0 3614 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1686
transform 1 0 3564 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1687
transform 1 0 3569 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1688
transform 1 0 3580 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1689
transform 1 0 3521 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1690
transform 1 0 3715 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1691
transform 1 0 3686 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1692
transform 1 0 3586 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1693
transform 1 0 3684 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1694
transform 1 0 3693 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1695
transform 1 0 3233 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1696
transform 1 0 3192 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1697
transform 1 0 3285 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1698
transform 1 0 3285 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1699
transform 1 0 3256 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1700
transform 1 0 3307 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1701
transform 1 0 3435 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1702
transform 1 0 3495 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1703
transform 1 0 3386 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1704
transform 1 0 3673 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1705
transform 1 0 3453 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1706
transform 1 0 3385 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1707
transform 1 0 3377 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1708
transform 1 0 3407 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1709
transform 1 0 3366 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1710
transform 1 0 3402 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1711
transform 1 0 3379 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1712
transform 1 0 3319 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1713
transform 1 0 3306 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1714
transform 1 0 3381 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1715
transform 1 0 3323 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1716
transform 1 0 3240 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1717
transform 1 0 3144 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-1718
transform 1 0 3257 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1719
transform 1 0 3361 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1720
transform 1 0 3435 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1721
transform 1 0 3554 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1722
transform 1 0 3527 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1723
transform 1 0 3536 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1724
transform 1 0 3565 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1725
transform 1 0 3551 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1726
transform 1 0 3552 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1727
transform 1 0 3215 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1728
transform 1 0 3322 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1729
transform 1 0 3396 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1730
transform 1 0 3452 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1731
transform 1 0 3291 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1732
transform 1 0 3251 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1733
transform 1 0 3299 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1734
transform 1 0 3254 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1735
transform 1 0 3273 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1736
transform 1 0 3259 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1737
transform 1 0 3247 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1738
transform 1 0 3309 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1739
transform 1 0 3112 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1740
transform 1 0 3137 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1741
transform 1 0 3147 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1742
transform 1 0 3167 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1743
transform 1 0 3216 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1744
transform 1 0 3470 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1745
transform 1 0 3664 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1746
transform 1 0 3705 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1747
transform 1 0 3609 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1748
transform 1 0 3606 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1749
transform 1 0 3674 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1750
transform 1 0 3689 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1751
transform 1 0 3499 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1752
transform 1 0 3558 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1753
transform 1 0 3237 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1754
transform 1 0 3231 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1755
transform 1 0 3240 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1756
transform 1 0 3175 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1757
transform 1 0 3209 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1758
transform 1 0 3203 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1759
transform 1 0 3505 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1760
transform 1 0 3457 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1761
transform 1 0 3441 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1762
transform 1 0 3423 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1763
transform 1 0 3341 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1764
transform 1 0 3258 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1765
transform 1 0 3198 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1766
transform 1 0 3146 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1767
transform 1 0 3060 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1768
transform 1 0 3104 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1769
transform 1 0 3057 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1770
transform 1 0 2989 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-1771
transform 1 0 3129 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1772
transform 1 0 3692 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1773
transform 1 0 3783 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1774
transform 1 0 3793 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1775
transform 1 0 3772 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1776
transform 1 0 3644 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1777
transform 1 0 3704 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1778
transform 1 0 3720 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1779
transform 1 0 3708 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1780
transform 1 0 3636 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1781
transform 1 0 3572 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1782
transform 1 0 3547 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1783
transform 1 0 3533 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1784
transform 1 0 3528 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1785
transform 1 0 3584 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1786
transform 1 0 3501 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1787
transform 1 0 3555 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1788
transform 1 0 3419 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1789
transform 1 0 3145 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1790
transform 1 0 3428 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1791
transform 1 0 3461 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1792
transform 1 0 3434 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1793
transform 1 0 3452 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1794
transform 1 0 3467 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1795
transform 1 0 3541 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1796
transform 1 0 3527 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1797
transform 1 0 3504 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1798
transform 1 0 3578 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1799
transform 1 0 3465 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1800
transform 1 0 3513 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1801
transform 1 0 3446 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1802
transform 1 0 3465 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1803
transform 1 0 3668 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1804
transform 1 0 3523 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1805
transform 1 0 3548 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1806
transform 1 0 3419 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1807
transform 1 0 3103 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-1808
transform 1 0 3137 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1809
transform 1 0 3119 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1810
transform 1 0 3104 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1811
transform 1 0 3143 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1812
transform 1 0 3120 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1813
transform 1 0 3100 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1814
transform 1 0 3007 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1815
transform 1 0 3494 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1816
transform 1 0 3505 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1817
transform 1 0 3594 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1818
transform 1 0 3621 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1819
transform 1 0 3618 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1820
transform 1 0 3500 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1821
transform 1 0 3575 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1822
transform 1 0 3561 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1823
transform 1 0 3567 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1824
transform 1 0 3590 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1825
transform 1 0 3510 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1826
transform 1 0 3156 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1827
transform 1 0 3160 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1828
transform 1 0 3223 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1829
transform 1 0 3243 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1830
transform 1 0 3522 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1831
transform 1 0 3076 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1832
transform 1 0 3098 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1833
transform 1 0 3111 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1834
transform 1 0 3107 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1835
transform 1 0 3297 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1836
transform 1 0 3082 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1837
transform 1 0 3107 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1838
transform 1 0 3117 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1839
transform 1 0 3113 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1840
transform 1 0 3180 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1841
transform 1 0 3114 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1842
transform 1 0 3203 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1843
transform 1 0 3255 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1844
transform 1 0 3198 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1845
transform 1 0 3272 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1846
transform 1 0 3232 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1847
transform 1 0 3303 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1848
transform 1 0 3297 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1849
transform 1 0 3303 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1850
transform 1 0 3233 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1851
transform 1 0 3261 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1852
transform 1 0 3209 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1853
transform 1 0 3201 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1854
transform 1 0 2820 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1855
transform 1 0 2974 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1856
transform 1 0 2996 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1857
transform 1 0 3012 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1858
transform 1 0 2988 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1859
transform 1 0 2978 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1860
transform 1 0 2981 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1861
transform 1 0 3003 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1862
transform 1 0 3030 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1863
transform 1 0 3025 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1864
transform 1 0 3093 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1865
transform 1 0 3019 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1866
transform 1 0 3113 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1867
transform 1 0 3076 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1868
transform 1 0 3144 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1869
transform 1 0 3128 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1870
transform 1 0 3129 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1871
transform 1 0 3038 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1872
transform 1 0 3092 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1873
transform 1 0 3095 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1874
transform 1 0 3111 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1875
transform 1 0 3075 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1876
transform 1 0 3015 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1877
transform 1 0 3001 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1878
transform 1 0 2994 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1879
transform 1 0 2970 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1880
transform 1 0 2929 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1881
transform 1 0 3417 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1882
transform 1 0 3708 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1883
transform 1 0 3604 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1884
transform 1 0 3623 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1885
transform 1 0 3191 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1886
transform 1 0 3267 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1887
transform 1 0 3273 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1888
transform 1 0 3291 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1889
transform 1 0 3214 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1890
transform 1 0 3251 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1891
transform 1 0 3162 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1892
transform 1 0 3243 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1893
transform 1 0 3179 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1894
transform 1 0 3165 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1895
transform 1 0 3149 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1896
transform 1 0 3118 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1897
transform 1 0 3110 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1898
transform 1 0 3125 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1899
transform 1 0 3149 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1900
transform 1 0 3126 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1901
transform 1 0 3014 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-1902
transform 1 0 3078 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1903
transform 1 0 3141 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1904
transform 1 0 3145 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1905
transform 1 0 3205 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1906
transform 1 0 3462 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1907
transform 1 0 3453 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1908
transform 1 0 3372 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1909
transform 1 0 3361 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1910
transform 1 0 3384 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1911
transform 1 0 3383 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1912
transform 1 0 3452 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1913
transform 1 0 3377 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1914
transform 1 0 3447 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1915
transform 1 0 3351 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1916
transform 1 0 3305 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1917
transform 1 0 3204 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1918
transform 1 0 3113 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-1919
transform 1 0 3126 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-1920
transform 1 0 3173 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1921
transform 1 0 3213 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1922
transform 1 0 3297 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1923
transform 1 0 3214 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-1924
transform 1 0 3295 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-1925
transform 1 0 3309 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1926
transform 1 0 3266 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1927
transform 1 0 3341 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1928
transform 1 0 3257 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1929
transform 1 0 3339 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1930
transform 1 0 3342 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1931
transform 1 0 3333 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1932
transform 1 0 3250 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1933
transform 1 0 3290 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1934
transform 1 0 3252 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1935
transform 1 0 3276 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1936
transform 1 0 3329 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1937
transform 1 0 3164 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1938
transform 1 0 3314 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1939
transform 1 0 3389 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1940
transform 1 0 3206 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1941
transform 1 0 3257 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1942
transform 1 0 3251 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1943
transform 1 0 3339 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1944
transform 1 0 3267 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1945
transform 1 0 3279 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-1946
transform 1 0 3202 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1947
transform 1 0 3239 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1948
transform 1 0 3150 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1949
transform 1 0 3228 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1950
transform 1 0 3161 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1951
transform 1 0 3342 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1952
transform 1 0 3137 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1953
transform 1 0 3245 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1954
transform 1 0 3376 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1955
transform 1 0 3450 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1956
transform 1 0 3536 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1957
transform 1 0 3506 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1958
transform 1 0 3518 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1959
transform 1 0 3571 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1960
transform 1 0 3704 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1961
transform 1 0 3706 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1962
transform 1 0 3738 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1963
transform 1 0 3825 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1964
transform 1 0 3131 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1965
transform 1 0 3076 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-1966
transform 1 0 3096 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-1967
transform 1 0 3117 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-1968
transform 1 0 3622 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-1969
transform 1 0 3031 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-1970
transform 1 0 3061 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1971
transform 1 0 3151 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-1972
transform 1 0 3195 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-1973
transform 1 0 3221 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-1974
transform 1 0 3209 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-1975
transform 1 0 3176 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1976
transform 1 0 3166 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1977
transform 1 0 3209 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1978
transform 1 0 3231 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1979
transform 1 0 3221 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1980
transform 1 0 3282 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1981
transform 1 0 3306 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1982
transform 1 0 3040 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-1983
transform 1 0 3085 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-1984
transform 1 0 3572 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1985
transform 1 0 3588 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-1986
transform 1 0 3549 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-1987
transform 1 0 3440 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-1988
transform 1 0 3320 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-1989
transform 1 0 3328 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-1990
transform 1 0 3230 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-1991
transform 1 0 3336 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-1992
transform 1 0 3338 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-1993
transform 1 0 3336 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-1994
transform 1 0 3332 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-1995
transform 1 0 3407 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-1996
transform 1 0 3269 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-1997
transform 1 0 3348 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-1998
transform 1 0 3366 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-1999
transform 1 0 3351 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2000
transform 1 0 3268 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2001
transform 1 0 3104 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2002
transform 1 0 3350 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2003
transform 1 0 3351 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2004
transform 1 0 3348 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2005
transform 1 0 3338 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2006
transform 1 0 3346 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2007
transform 1 0 3411 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2008
transform 1 0 3519 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2009
transform 1 0 3399 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2010
transform 1 0 3386 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2011
transform 1 0 3317 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2012
transform 1 0 3363 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2013
transform 1 0 3324 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2014
transform 1 0 3350 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2015
transform 1 0 3355 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2016
transform 1 0 3417 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2017
transform 1 0 3414 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2018
transform 1 0 3489 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2019
transform 1 0 3292 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2020
transform 1 0 3302 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2021
transform 1 0 3258 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2022
transform 1 0 3306 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2023
transform 1 0 3239 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2024
transform 1 0 3261 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2025
transform 1 0 3227 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2026
transform 1 0 3298 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2027
transform 1 0 3311 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2028
transform 1 0 3296 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2029
transform 1 0 3341 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2030
transform 1 0 3285 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2031
transform 1 0 3214 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2032
transform 1 0 3106 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2033
transform 1 0 3298 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2034
transform 1 0 3314 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2035
transform 1 0 3264 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2036
transform 1 0 3312 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2037
transform 1 0 2890 0 1 8734
box 0 0 3 6
use FEEDTHRU  F-2038
transform 1 0 3131 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2039
transform 1 0 3090 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2040
transform 1 0 3011 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-2041
transform 1 0 2962 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-2042
transform 1 0 3137 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2043
transform 1 0 3159 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2044
transform 1 0 3180 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2045
transform 1 0 3178 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2046
transform 1 0 3783 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2047
transform 1 0 3627 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2048
transform 1 0 3669 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2049
transform 1 0 3524 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2050
transform 1 0 3240 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2051
transform 1 0 3263 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2052
transform 1 0 3285 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2053
transform 1 0 3269 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2054
transform 1 0 3205 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2055
transform 1 0 3212 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2056
transform 1 0 3227 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2057
transform 1 0 3227 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2058
transform 1 0 3201 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2059
transform 1 0 3169 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2060
transform 1 0 3333 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2061
transform 1 0 3288 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2062
transform 1 0 3332 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2063
transform 1 0 3345 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2064
transform 1 0 3269 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2065
transform 1 0 3315 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2066
transform 1 0 3275 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2067
transform 1 0 3217 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2068
transform 1 0 3224 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2069
transform 1 0 3239 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2070
transform 1 0 3233 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2071
transform 1 0 2998 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-2072
transform 1 0 3062 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-2073
transform 1 0 2977 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-2074
transform 1 0 3029 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-2075
transform 1 0 3075 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2076
transform 1 0 3122 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2077
transform 1 0 3189 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2078
transform 1 0 3200 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2079
transform 1 0 3153 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2080
transform 1 0 3201 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2081
transform 1 0 3210 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2082
transform 1 0 3202 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2083
transform 1 0 3283 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2084
transform 1 0 3315 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2085
transform 1 0 3278 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2086
transform 1 0 3365 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2087
transform 1 0 3281 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2088
transform 1 0 3372 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2089
transform 1 0 3396 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2090
transform 1 0 3387 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2091
transform 1 0 3207 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2092
transform 1 0 3216 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2093
transform 1 0 3208 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2094
transform 1 0 3289 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2095
transform 1 0 3330 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2096
transform 1 0 3314 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2097
transform 1 0 3377 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2098
transform 1 0 3287 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2099
transform 1 0 3224 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2100
transform 1 0 3214 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2101
transform 1 0 3146 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2102
transform 1 0 3149 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2103
transform 1 0 3226 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2104
transform 1 0 3509 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2105
transform 1 0 3414 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2106
transform 1 0 3447 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2107
transform 1 0 3635 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2108
transform 1 0 3129 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2109
transform 1 0 3117 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2110
transform 1 0 3396 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2111
transform 1 0 3401 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2112
transform 1 0 3659 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2113
transform 1 0 3694 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2114
transform 1 0 3627 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2115
transform 1 0 3537 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2116
transform 1 0 3174 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2117
transform 1 0 3071 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2118
transform 1 0 3119 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2119
transform 1 0 3125 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2120
transform 1 0 3147 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2121
transform 1 0 3102 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2122
transform 1 0 3048 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2123
transform 1 0 3041 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2124
transform 1 0 3030 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2125
transform 1 0 3004 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2126
transform 1 0 2953 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2127
transform 1 0 2808 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-2128
transform 1 0 3143 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2129
transform 1 0 3153 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2130
transform 1 0 3590 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2131
transform 1 0 3563 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2132
transform 1 0 3506 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2133
transform 1 0 3559 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2134
transform 1 0 3545 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2135
transform 1 0 3534 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2136
transform 1 0 3548 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2137
transform 1 0 3579 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2138
transform 1 0 3507 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2139
transform 1 0 3524 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2140
transform 1 0 3547 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2141
transform 1 0 3660 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2142
transform 1 0 3503 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2143
transform 1 0 3438 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2144
transform 1 0 3364 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2145
transform 1 0 3233 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2146
transform 1 0 3605 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2147
transform 1 0 3411 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2148
transform 1 0 3353 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2149
transform 1 0 3393 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2150
transform 1 0 3419 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2151
transform 1 0 3589 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2152
transform 1 0 3144 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2153
transform 1 0 3179 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2154
transform 1 0 3155 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2155
transform 1 0 3152 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2156
transform 1 0 3142 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2157
transform 1 0 3173 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2158
transform 1 0 3183 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2159
transform 1 0 3185 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2160
transform 1 0 3423 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2161
transform 1 0 3365 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2162
transform 1 0 3387 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2163
transform 1 0 3395 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2164
transform 1 0 3430 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2165
transform 1 0 3327 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2166
transform 1 0 3410 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2167
transform 1 0 3492 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2168
transform 1 0 3534 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2169
transform 1 0 3523 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2170
transform 1 0 3580 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2171
transform 1 0 3564 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2172
transform 1 0 3605 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2173
transform 1 0 3593 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2174
transform 1 0 3512 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2175
transform 1 0 3654 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2176
transform 1 0 3663 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2177
transform 1 0 3624 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2178
transform 1 0 3529 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2179
transform 1 0 3300 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2180
transform 1 0 3243 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2181
transform 1 0 3232 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2182
transform 1 0 3273 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2183
transform 1 0 3168 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2184
transform 1 0 3083 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-2185
transform 1 0 3748 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2186
transform 1 0 3732 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2187
transform 1 0 3628 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2188
transform 1 0 3647 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2189
transform 1 0 3400 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2190
transform 1 0 3371 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2191
transform 1 0 3382 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2192
transform 1 0 3344 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2193
transform 1 0 3386 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2194
transform 1 0 3584 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2195
transform 1 0 3551 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2196
transform 1 0 3455 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2197
transform 1 0 3588 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2198
transform 1 0 3597 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2199
transform 1 0 3588 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2200
transform 1 0 3493 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2201
transform 1 0 3452 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2202
transform 1 0 3552 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2203
transform 1 0 3552 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2204
transform 1 0 3575 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2205
transform 1 0 3555 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2206
transform 1 0 3554 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2207
transform 1 0 3568 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2208
transform 1 0 3455 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2209
transform 1 0 3446 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2210
transform 1 0 3031 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2211
transform 1 0 3133 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2212
transform 1 0 3171 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2213
transform 1 0 3215 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2214
transform 1 0 3191 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2215
transform 1 0 3194 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2216
transform 1 0 3172 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2217
transform 1 0 3215 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2218
transform 1 0 3243 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2219
transform 1 0 3233 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2220
transform 1 0 3324 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2221
transform 1 0 3240 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2222
transform 1 0 3037 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2223
transform 1 0 3004 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-2224
transform 1 0 3194 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2225
transform 1 0 3319 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2226
transform 1 0 3387 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2227
transform 1 0 3440 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2228
transform 1 0 3121 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-2229
transform 1 0 3335 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2230
transform 1 0 3296 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2231
transform 1 0 3329 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2232
transform 1 0 3302 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2233
transform 1 0 3308 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2234
transform 1 0 3368 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2235
transform 1 0 3001 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-2236
transform 1 0 3016 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2237
transform 1 0 3740 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2238
transform 1 0 3173 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2239
transform 1 0 3197 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2240
transform 1 0 3017 0 1 8734
box 0 0 3 6
use FEEDTHRU  F-2241
transform 1 0 3294 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2242
transform 1 0 3168 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2243
transform 1 0 3278 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2244
transform 1 0 3177 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2245
transform 1 0 3192 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2246
transform 1 0 3381 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2247
transform 1 0 3399 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2248
transform 1 0 3328 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2249
transform 1 0 3356 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2250
transform 1 0 3267 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2251
transform 1 0 3158 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2252
transform 1 0 3477 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2253
transform 1 0 3483 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2254
transform 1 0 3431 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2255
transform 1 0 3429 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2256
transform 1 0 3455 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2257
transform 1 0 3330 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2258
transform 1 0 3210 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2259
transform 1 0 3560 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2260
transform 1 0 3672 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2261
transform 1 0 3139 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2262
transform 1 0 3193 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2263
transform 1 0 3264 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2264
transform 1 0 3505 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2265
transform 1 0 3458 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2266
transform 1 0 3402 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2267
transform 1 0 3328 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2268
transform 1 0 3449 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2269
transform 1 0 3466 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2270
transform 1 0 3461 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2271
transform 1 0 3447 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2272
transform 1 0 3443 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2273
transform 1 0 3349 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2274
transform 1 0 3291 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2275
transform 1 0 3315 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2276
transform 1 0 3221 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2277
transform 1 0 3269 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2278
transform 1 0 3272 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2279
transform 1 0 3267 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2280
transform 1 0 3345 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2281
transform 1 0 3327 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2282
transform 1 0 3327 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2283
transform 1 0 3262 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2284
transform 1 0 3249 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2285
transform 1 0 3261 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2286
transform 1 0 3273 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2287
transform 1 0 3155 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2288
transform 1 0 3209 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2289
transform 1 0 3233 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2290
transform 1 0 3234 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2291
transform 1 0 3202 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2292
transform 1 0 3142 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2293
transform 1 0 3177 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2294
transform 1 0 3114 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2295
transform 1 0 3082 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2296
transform 1 0 3279 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2297
transform 1 0 3248 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2298
transform 1 0 3227 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2299
transform 1 0 3173 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2300
transform 1 0 3297 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2301
transform 1 0 3542 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2302
transform 1 0 3536 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2303
transform 1 0 3856 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2304
transform 1 0 3301 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2305
transform 1 0 3234 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2306
transform 1 0 3219 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2307
transform 1 0 3185 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2308
transform 1 0 3574 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2309
transform 1 0 3399 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2310
transform 1 0 3411 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2311
transform 1 0 3436 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2312
transform 1 0 3431 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2313
transform 1 0 3410 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2314
transform 1 0 3525 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2315
transform 1 0 3474 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2316
transform 1 0 3471 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2317
transform 1 0 3425 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2318
transform 1 0 3414 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2319
transform 1 0 3263 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2320
transform 1 0 3284 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2321
transform 1 0 3279 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2322
transform 1 0 3257 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2323
transform 1 0 3203 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2324
transform 1 0 3333 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2325
transform 1 0 3309 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2326
transform 1 0 3492 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2327
transform 1 0 3472 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2328
transform 1 0 3538 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2329
transform 1 0 3606 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2330
transform 1 0 3626 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2331
transform 1 0 3569 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2332
transform 1 0 3506 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2333
transform 1 0 3648 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2334
transform 1 0 3645 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2335
transform 1 0 3642 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2336
transform 1 0 3522 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2337
transform 1 0 3447 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2338
transform 1 0 3513 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2339
transform 1 0 3519 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2340
transform 1 0 3484 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2341
transform 1 0 3550 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2342
transform 1 0 3624 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2343
transform 1 0 3790 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2344
transform 1 0 3581 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2345
transform 1 0 3518 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2346
transform 1 0 3660 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2347
transform 1 0 3687 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2348
transform 1 0 3666 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2349
transform 1 0 3562 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2350
transform 1 0 3578 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2351
transform 1 0 3543 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2352
transform 1 0 3651 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2353
transform 1 0 3542 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2354
transform 1 0 3516 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2355
transform 1 0 3521 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2356
transform 1 0 3529 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2357
transform 1 0 3500 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2358
transform 1 0 3500 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2359
transform 1 0 3539 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2360
transform 1 0 3064 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-2361
transform 1 0 3137 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2362
transform 1 0 3223 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2363
transform 1 0 3252 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2364
transform 1 0 3353 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2365
transform 1 0 3341 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2366
transform 1 0 3287 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2367
transform 1 0 3343 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2368
transform 1 0 3341 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2369
transform 1 0 3131 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2370
transform 1 0 3217 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2371
transform 1 0 3717 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2372
transform 1 0 3164 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-2373
transform 1 0 3270 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2374
transform 1 0 3453 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2375
transform 1 0 3450 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2376
transform 1 0 3459 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2377
transform 1 0 3285 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2378
transform 1 0 3241 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2379
transform 1 0 3199 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2380
transform 1 0 3139 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2381
transform 1 0 3174 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2382
transform 1 0 3512 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2383
transform 1 0 3507 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2384
transform 1 0 3421 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2385
transform 1 0 3216 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2386
transform 1 0 3320 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2387
transform 1 0 3280 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2388
transform 1 0 3369 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2389
transform 1 0 3354 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2390
transform 1 0 3366 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2391
transform 1 0 3239 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2392
transform 1 0 3293 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2393
transform 1 0 3326 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2394
transform 1 0 3321 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2395
transform 1 0 3271 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2396
transform 1 0 3196 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2397
transform 1 0 3240 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2398
transform 1 0 3183 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2399
transform 1 0 3143 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2400
transform 1 0 3600 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2401
transform 1 0 3503 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2402
transform 1 0 3492 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2403
transform 1 0 3442 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2404
transform 1 0 3370 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2405
transform 1 0 3420 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2406
transform 1 0 3369 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2407
transform 1 0 3320 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2408
transform 1 0 3327 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2409
transform 1 0 3097 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2410
transform 1 0 3055 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-2411
transform 1 0 2980 0 1 8734
box 0 0 3 6
use FEEDTHRU  F-2412
transform 1 0 3303 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2413
transform 1 0 3315 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2414
transform 1 0 3141 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2415
transform 1 0 3198 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2416
transform 1 0 3599 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2417
transform 1 0 3624 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2418
transform 1 0 3633 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2419
transform 1 0 3239 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2420
transform 1 0 3285 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2421
transform 1 0 3318 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2422
transform 1 0 3262 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2423
transform 1 0 3337 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2424
transform 1 0 3515 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2425
transform 1 0 3294 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2426
transform 1 0 3374 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2427
transform 1 0 3420 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2428
transform 1 0 3489 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2429
transform 1 0 3714 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2430
transform 1 0 3531 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2431
transform 1 0 3749 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2432
transform 1 0 3799 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2433
transform 1 0 3534 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2434
transform 1 0 3593 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2435
transform 1 0 3568 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2436
transform 1 0 3852 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2437
transform 1 0 3669 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2438
transform 1 0 3711 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2439
transform 1 0 3554 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2440
transform 1 0 3522 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2441
transform 1 0 3213 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2442
transform 1 0 3227 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2443
transform 1 0 3357 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2444
transform 1 0 3219 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2445
transform 1 0 3203 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2446
transform 1 0 3160 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2447
transform 1 0 3316 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2448
transform 1 0 3405 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2449
transform 1 0 3251 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2450
transform 1 0 3266 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2451
transform 1 0 3253 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2452
transform 1 0 3580 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2453
transform 1 0 3767 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2454
transform 1 0 3537 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2455
transform 1 0 3476 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2456
transform 1 0 3481 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2457
transform 1 0 3570 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2458
transform 1 0 3585 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2459
transform 1 0 3570 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2460
transform 1 0 3443 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2461
transform 1 0 3506 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2462
transform 1 0 3545 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2463
transform 1 0 3528 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2464
transform 1 0 3571 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2465
transform 1 0 3376 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2466
transform 1 0 3426 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2467
transform 1 0 3375 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2468
transform 1 0 3476 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2469
transform 1 0 3440 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2470
transform 1 0 3434 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2471
transform 1 0 3434 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2472
transform 1 0 3428 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2473
transform 1 0 3454 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2474
transform 1 0 3449 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2475
transform 1 0 3435 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2476
transform 1 0 3461 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2477
transform 1 0 3573 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2478
transform 1 0 3426 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2479
transform 1 0 3189 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2480
transform 1 0 3004 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-2481
transform 1 0 3068 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-2482
transform 1 0 3132 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2483
transform 1 0 3179 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2484
transform 1 0 3275 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2485
transform 1 0 3260 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2486
transform 1 0 3299 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2487
transform 1 0 3302 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2488
transform 1 0 3427 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2489
transform 1 0 3684 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2490
transform 1 0 3666 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2491
transform 1 0 3681 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2492
transform 1 0 3681 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2493
transform 1 0 3177 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2494
transform 1 0 3473 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2495
transform 1 0 3348 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2496
transform 1 0 3282 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2497
transform 1 0 3487 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2498
transform 1 0 3553 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2499
transform 1 0 3627 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2500
transform 1 0 3179 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2501
transform 1 0 3195 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2502
transform 1 0 3203 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2503
transform 1 0 3339 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2504
transform 1 0 3174 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2505
transform 1 0 3277 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2506
transform 1 0 3348 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2507
transform 1 0 3250 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2508
transform 1 0 3215 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2509
transform 1 0 3321 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2510
transform 1 0 3327 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2511
transform 1 0 3185 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2512
transform 1 0 3239 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2513
transform 1 0 3290 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2514
transform 1 0 3297 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2515
transform 1 0 3229 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2516
transform 1 0 3276 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2517
transform 1 0 3243 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2518
transform 1 0 3209 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2519
transform 1 0 3288 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2520
transform 1 0 3238 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2521
transform 1 0 3313 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2522
transform 1 0 3294 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2523
transform 1 0 3244 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2524
transform 1 0 3319 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2525
transform 1 0 3390 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2526
transform 1 0 3389 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2527
transform 1 0 3359 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2528
transform 1 0 3293 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2529
transform 1 0 3441 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2530
transform 1 0 3438 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2531
transform 1 0 3429 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2532
transform 1 0 3340 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2533
transform 1 0 3190 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2534
transform 1 0 3188 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2535
transform 1 0 3203 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2536
transform 1 0 3295 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2537
transform 1 0 3357 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2538
transform 1 0 3327 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2539
transform 1 0 3293 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2540
transform 1 0 3216 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2541
transform 1 0 3313 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2542
transform 1 0 3385 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2543
transform 1 0 3456 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2544
transform 1 0 3461 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2545
transform 1 0 3440 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2546
transform 1 0 3593 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2547
transform 1 0 3528 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2548
transform 1 0 3504 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2549
transform 1 0 3477 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2550
transform 1 0 3369 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2551
transform 1 0 3303 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2552
transform 1 0 3269 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2553
transform 1 0 3235 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2554
transform 1 0 3245 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2555
transform 1 0 3149 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2556
transform 1 0 3405 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2557
transform 1 0 3425 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2558
transform 1 0 3622 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2559
transform 1 0 3605 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2560
transform 1 0 3573 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2561
transform 1 0 3424 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2562
transform 1 0 3666 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2563
transform 1 0 3582 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2564
transform 1 0 3599 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2565
transform 1 0 3539 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2566
transform 1 0 3467 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2567
transform 1 0 3612 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2568
transform 1 0 3627 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2569
transform 1 0 3612 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2570
transform 1 0 3511 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2571
transform 1 0 3530 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2572
transform 1 0 3450 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2573
transform 1 0 3639 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2574
transform 1 0 3412 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2575
transform 1 0 3484 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2576
transform 1 0 3570 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2577
transform 1 0 3587 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2578
transform 1 0 3269 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2579
transform 1 0 3341 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2580
transform 1 0 3459 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2581
transform 1 0 3323 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2582
transform 1 0 3339 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2583
transform 1 0 3244 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2584
transform 1 0 3336 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2585
transform 1 0 3345 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2586
transform 1 0 3449 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2587
transform 1 0 3615 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2588
transform 1 0 3432 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2589
transform 1 0 3506 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2590
transform 1 0 3249 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2591
transform 1 0 3251 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2592
transform 1 0 3405 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2593
transform 1 0 3234 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2594
transform 1 0 3344 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2595
transform 1 0 3304 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2596
transform 1 0 3255 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2597
transform 1 0 3239 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2598
transform 1 0 3229 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2599
transform 1 0 3218 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2600
transform 1 0 3245 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2601
transform 1 0 3272 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2602
transform 1 0 3210 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2603
transform 1 0 3181 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2604
transform 1 0 3094 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2605
transform 1 0 3037 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-2606
transform 1 0 3642 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2607
transform 1 0 3657 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2608
transform 1 0 3654 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2609
transform 1 0 3541 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2610
transform 1 0 3560 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2611
transform 1 0 3489 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2612
transform 1 0 3563 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2613
transform 1 0 3223 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2614
transform 1 0 3195 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2615
transform 1 0 3391 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2616
transform 1 0 3465 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2617
transform 1 0 3524 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2618
transform 1 0 3479 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2619
transform 1 0 3476 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2620
transform 1 0 3511 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2621
transform 1 0 3500 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2622
transform 1 0 3486 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2623
transform 1 0 3485 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2624
transform 1 0 3657 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2625
transform 1 0 3474 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2626
transform 1 0 3554 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2627
transform 1 0 3535 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2628
transform 1 0 3648 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2629
transform 1 0 3651 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2630
transform 1 0 3636 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2631
transform 1 0 3488 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2632
transform 1 0 3557 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2633
transform 1 0 3614 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2634
transform 1 0 3594 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2635
transform 1 0 3508 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2636
transform 1 0 3436 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2637
transform 1 0 3483 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2638
transform 1 0 3450 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2639
transform 1 0 3371 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2640
transform 1 0 3558 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2641
transform 1 0 3282 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2642
transform 1 0 3678 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2643
transform 1 0 3557 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2644
transform 1 0 3690 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2645
transform 1 0 3518 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2646
transform 1 0 3525 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2647
transform 1 0 3480 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2648
transform 1 0 3684 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2649
transform 1 0 3512 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2650
transform 1 0 3492 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2651
transform 1 0 3506 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2652
transform 1 0 3777 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2653
transform 1 0 3482 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2654
transform 1 0 3485 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2655
transform 1 0 3632 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2656
transform 1 0 3474 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2657
transform 1 0 3400 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2658
transform 1 0 3251 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2659
transform 1 0 3566 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2660
transform 1 0 3365 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2661
transform 1 0 3311 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2662
transform 1 0 3263 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2663
transform 1 0 3393 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2664
transform 1 0 3426 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2665
transform 1 0 3405 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2666
transform 1 0 3275 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2667
transform 1 0 3317 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2668
transform 1 0 3362 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2669
transform 1 0 3378 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2670
transform 1 0 3053 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-2671
transform 1 0 3144 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2672
transform 1 0 3470 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2673
transform 1 0 3539 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2674
transform 1 0 3525 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2675
transform 1 0 3407 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2676
transform 1 0 3464 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2677
transform 1 0 3488 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2678
transform 1 0 3471 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2679
transform 1 0 3494 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2680
transform 1 0 3663 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2681
transform 1 0 3462 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2682
transform 1 0 3548 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2683
transform 1 0 3523 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2684
transform 1 0 3630 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2685
transform 1 0 2986 0 1 8734
box 0 0 3 6
use FEEDTHRU  F-2686
transform 1 0 3386 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2687
transform 1 0 3374 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2688
transform 1 0 3360 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2689
transform 1 0 3360 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2690
transform 1 0 3357 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2691
transform 1 0 3256 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2692
transform 1 0 3308 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2693
transform 1 0 3180 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2694
transform 1 0 3369 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2695
transform 1 0 3215 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2696
transform 1 0 3207 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2697
transform 1 0 3191 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2698
transform 1 0 3178 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2699
transform 1 0 3170 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2700
transform 1 0 3185 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2701
transform 1 0 3209 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2702
transform 1 0 3156 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2703
transform 1 0 3130 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2704
transform 1 0 3106 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-2705
transform 1 0 3185 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2706
transform 1 0 3259 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2707
transform 1 0 3312 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2708
transform 1 0 3416 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2709
transform 1 0 3398 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2710
transform 1 0 3464 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2711
transform 1 0 3394 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2712
transform 1 0 3383 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2713
transform 1 0 3381 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2714
transform 1 0 3389 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2715
transform 1 0 3525 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2716
transform 1 0 3085 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-2717
transform 1 0 3155 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2718
transform 1 0 3253 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2719
transform 1 0 3294 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2720
transform 1 0 3392 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2721
transform 1 0 3371 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2722
transform 1 0 3350 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2723
transform 1 0 3388 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2724
transform 1 0 3377 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2725
transform 1 0 3375 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2726
transform 1 0 3383 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2727
transform 1 0 3507 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2728
transform 1 0 3336 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2729
transform 1 0 3425 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2730
transform 1 0 3418 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2731
transform 1 0 2998 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-2732
transform 1 0 3509 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2733
transform 1 0 3572 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2734
transform 1 0 3629 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2735
transform 1 0 3609 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2736
transform 1 0 3541 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2737
transform 1 0 3475 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2738
transform 1 0 3007 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-2739
transform 1 0 3043 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2740
transform 1 0 3157 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2741
transform 1 0 3183 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2742
transform 1 0 3239 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2743
transform 1 0 3013 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-2744
transform 1 0 3049 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2745
transform 1 0 3163 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2746
transform 1 0 3189 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2747
transform 1 0 3245 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2748
transform 1 0 3221 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2749
transform 1 0 3200 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2750
transform 1 0 3211 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2751
transform 1 0 3221 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2752
transform 1 0 3237 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2753
transform 1 0 3409 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2754
transform 1 0 3337 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2755
transform 1 0 3387 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2756
transform 1 0 3321 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2757
transform 1 0 3338 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2758
transform 1 0 3255 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2759
transform 1 0 3326 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2760
transform 1 0 3344 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2761
transform 1 0 3284 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2762
transform 1 0 3350 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2763
transform 1 0 3264 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2764
transform 1 0 3362 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2765
transform 1 0 3338 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2766
transform 1 0 3346 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2767
transform 1 0 3324 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2768
transform 1 0 3265 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2769
transform 1 0 3540 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2770
transform 1 0 3251 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2771
transform 1 0 3441 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2772
transform 1 0 3314 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2773
transform 1 0 3267 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2774
transform 1 0 3481 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2775
transform 1 0 3352 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2776
transform 1 0 3402 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2777
transform 1 0 3339 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2778
transform 1 0 3311 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2779
transform 1 0 3305 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2780
transform 1 0 3297 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2781
transform 1 0 3281 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2782
transform 1 0 3265 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2783
transform 1 0 3266 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2784
transform 1 0 3269 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2785
transform 1 0 3308 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2786
transform 1 0 3246 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2787
transform 1 0 3211 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2788
transform 1 0 3103 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2789
transform 1 0 3052 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-2790
transform 1 0 3353 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2791
transform 1 0 3281 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2792
transform 1 0 3348 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2793
transform 1 0 3350 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2794
transform 1 0 3287 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2795
transform 1 0 3248 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2796
transform 1 0 3378 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2797
transform 1 0 3393 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2798
transform 1 0 3384 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2799
transform 1 0 3354 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2800
transform 1 0 3277 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2801
transform 1 0 3398 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2802
transform 1 0 3353 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2803
transform 1 0 3356 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2804
transform 1 0 3376 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2805
transform 1 0 3312 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2806
transform 1 0 3231 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2807
transform 1 0 3197 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2808
transform 1 0 3150 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2809
transform 1 0 3065 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-2810
transform 1 0 3001 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-2811
transform 1 0 3420 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2812
transform 1 0 3349 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2813
transform 1 0 3274 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2814
transform 1 0 3330 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2815
transform 1 0 3261 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2816
transform 1 0 3221 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2817
transform 1 0 3174 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2818
transform 1 0 3271 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2819
transform 1 0 3287 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2820
transform 1 0 3303 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2821
transform 1 0 3348 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2822
transform 1 0 3435 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2823
transform 1 0 3384 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2824
transform 1 0 3390 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2825
transform 1 0 3381 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2826
transform 1 0 3274 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2827
transform 1 0 3228 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2828
transform 1 0 3429 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2829
transform 1 0 3275 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2830
transform 1 0 3273 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2831
transform 1 0 3263 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2832
transform 1 0 3100 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-2833
transform 1 0 3280 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2834
transform 1 0 3366 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2835
transform 1 0 3478 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2836
transform 1 0 3467 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2837
transform 1 0 3472 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2838
transform 1 0 3344 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2839
transform 1 0 3305 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2840
transform 1 0 3320 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2841
transform 1 0 3399 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2842
transform 1 0 3245 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2843
transform 1 0 3204 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2844
transform 1 0 3744 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2845
transform 1 0 3633 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2846
transform 1 0 3464 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2847
transform 1 0 3595 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2848
transform 1 0 3546 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2849
transform 1 0 3573 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2850
transform 1 0 3552 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2851
transform 1 0 3389 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2852
transform 1 0 3360 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2853
transform 1 0 3458 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2854
transform 1 0 3433 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2855
transform 1 0 3534 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2856
transform 1 0 3561 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2857
transform 1 0 3540 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2858
transform 1 0 3411 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2859
transform 1 0 3420 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2860
transform 1 0 3357 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2861
transform 1 0 3432 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2862
transform 1 0 3382 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2863
transform 1 0 3454 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2864
transform 1 0 3546 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2865
transform 1 0 3557 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2866
transform 1 0 3414 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2867
transform 1 0 3364 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2868
transform 1 0 3430 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2869
transform 1 0 3522 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2870
transform 1 0 3533 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2871
transform 1 0 3458 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2872
transform 1 0 3395 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2873
transform 1 0 3546 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2874
transform 1 0 3567 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2875
transform 1 0 3540 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2876
transform 1 0 3407 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2877
transform 1 0 3412 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2878
transform 1 0 3398 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2879
transform 1 0 3672 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2880
transform 1 0 3553 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2881
transform 1 0 3584 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2882
transform 1 0 3486 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2883
transform 1 0 3696 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2884
transform 1 0 3345 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2885
transform 1 0 3264 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2886
transform 1 0 3263 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2887
transform 1 0 3210 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2888
transform 1 0 3119 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-2889
transform 1 0 3034 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-2890
transform 1 0 3480 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2891
transform 1 0 3489 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2892
transform 1 0 3452 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2893
transform 1 0 3383 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2894
transform 1 0 3431 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2895
transform 1 0 3450 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2896
transform 1 0 3367 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2897
transform 1 0 3301 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2898
transform 1 0 3363 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2899
transform 1 0 3267 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-2900
transform 1 0 3233 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-2901
transform 1 0 3183 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-2902
transform 1 0 3089 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-2903
transform 1 0 3486 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2904
transform 1 0 3540 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2905
transform 1 0 3669 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2906
transform 1 0 3491 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2907
transform 1 0 3477 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2908
transform 1 0 3479 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2909
transform 1 0 3484 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2910
transform 1 0 3473 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2911
transform 1 0 3458 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2912
transform 1 0 3521 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2913
transform 1 0 3471 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2914
transform 1 0 3397 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2915
transform 1 0 3248 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-2916
transform 1 0 3417 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2917
transform 1 0 3257 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2918
transform 1 0 3323 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2919
transform 1 0 3395 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2920
transform 1 0 3215 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2921
transform 1 0 3263 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2922
transform 1 0 3207 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2923
transform 1 0 3257 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2924
transform 1 0 3564 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2925
transform 1 0 3579 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2926
transform 1 0 3558 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2927
transform 1 0 3531 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2928
transform 1 0 3330 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2929
transform 1 0 3446 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2930
transform 1 0 3542 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2931
transform 1 0 3218 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2932
transform 1 0 3215 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2933
transform 1 0 3055 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-2934
transform 1 0 3143 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-2935
transform 1 0 3504 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2936
transform 1 0 3509 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2937
transform 1 0 3431 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2938
transform 1 0 3395 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2939
transform 1 0 3353 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2940
transform 1 0 3507 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2941
transform 1 0 3528 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2942
transform 1 0 3486 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2943
transform 1 0 3400 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2944
transform 1 0 3428 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2945
transform 1 0 3294 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2946
transform 1 0 3527 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-2947
transform 1 0 3571 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2948
transform 1 0 3494 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2949
transform 1 0 3425 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2950
transform 1 0 3440 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2951
transform 1 0 3709 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2952
transform 1 0 3698 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2953
transform 1 0 3441 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2954
transform 1 0 3455 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2955
transform 1 0 3633 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2956
transform 1 0 3408 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2957
transform 1 0 3518 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2958
transform 1 0 3487 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2959
transform 1 0 3600 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2960
transform 1 0 3603 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-2961
transform 1 0 3651 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2962
transform 1 0 3425 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2963
transform 1 0 3488 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2964
transform 1 0 3569 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2965
transform 1 0 3558 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-2966
transform 1 0 3466 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-2967
transform 1 0 3400 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-2968
transform 1 0 3450 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-2969
transform 1 0 3437 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2970
transform 1 0 3621 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2971
transform 1 0 3390 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2972
transform 1 0 3500 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-2973
transform 1 0 3463 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-2974
transform 1 0 3582 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-2975
transform 1 0 3407 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2976
transform 1 0 3609 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2977
transform 1 0 3372 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-2978
transform 1 0 3291 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-2979
transform 1 0 3293 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-2980
transform 1 0 3471 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-2981
transform 1 0 3293 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-2982
transform 1 0 3301 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2983
transform 1 0 3314 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2984
transform 1 0 3270 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-2985
transform 1 0 3332 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2986
transform 1 0 3281 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2987
transform 1 0 3296 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2988
transform 1 0 3289 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2989
transform 1 0 3473 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-2990
transform 1 0 3524 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-2991
transform 1 0 3611 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-2992
transform 1 0 3284 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-2993
transform 1 0 3233 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-2994
transform 1 0 3236 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2995
transform 1 0 3471 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-2996
transform 1 0 3202 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2997
transform 1 0 3283 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-2998
transform 1 0 3290 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-2999
transform 1 0 3543 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-3000
transform 1 0 3359 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-3001
transform 1 0 3357 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-3002
transform 1 0 3347 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-3003
transform 1 0 3352 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-3004
transform 1 0 3300 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-3005
transform 1 0 3537 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-3006
transform 1 0 3401 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-3007
transform 1 0 3485 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-3008
transform 1 0 3480 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-3009
transform 1 0 3391 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-3010
transform 1 0 3325 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-3011
transform 1 0 3381 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-3012
transform 1 0 3279 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-3013
transform 1 0 3245 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-3014
transform 1 0 3195 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-3015
transform 1 0 3101 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-3016
transform 1 0 3491 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-3017
transform 1 0 3486 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-3018
transform 1 0 3397 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-3019
transform 1 0 3331 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-3020
transform 1 0 3778 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-3021
transform 1 0 3722 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-3022
transform 1 0 3482 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-3023
transform 1 0 3705 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-3024
transform 1 0 3451 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-3025
transform 1 0 3482 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-3026
transform 1 0 3366 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-3027
transform 1 0 3603 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-3028
transform 1 0 3419 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-3029
transform 1 0 3417 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-3030
transform 1 0 3584 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-3031
transform 1 0 3418 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-3032
transform 1 0 3718 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-3033
transform 1 0 3401 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-3034
transform 1 0 3470 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-3035
transform 1 0 3456 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-3036
transform 1 0 3388 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-3037
transform 1 0 3269 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-3038
transform 1 0 3576 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-3039
transform 1 0 3329 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-3040
transform 1 0 3380 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-3041
transform 1 0 3318 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-3042
transform 1 0 3114 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-3043
transform 1 0 3167 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-3044
transform 1 0 3026 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-3045
transform 1 0 3120 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-3046
transform 1 0 3316 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-3047
transform 1 0 3384 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-3048
transform 1 0 3807 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-3049
transform 1 0 3585 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-3050
transform 1 0 3342 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-3051
transform 1 0 3615 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-3052
transform 1 0 3600 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-3053
transform 1 0 3431 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-3054
transform 1 0 3476 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-3055
transform 1 0 3516 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-3056
transform 1 0 3498 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-3057
transform 1 0 3367 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-3058
transform 1 0 3254 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-3059
transform 1 0 3241 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-3060
transform 1 0 3247 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-3061
transform 1 0 3314 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-3062
transform 1 0 3342 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-3063
transform 1 0 3408 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-3064
transform 1 0 3358 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-3065
transform 1 0 3424 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-3066
transform 1 0 3516 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-3067
transform 1 0 3521 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-3068
transform 1 0 3275 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-3069
transform 1 0 3309 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-3070
transform 1 0 3282 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-3071
transform 1 0 3338 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-3072
transform 1 0 3293 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-3073
transform 1 0 3308 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-3074
transform 1 0 3295 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-3075
transform 1 0 3421 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-3076
transform 1 0 3552 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-3077
transform 1 0 3237 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-3078
transform 1 0 3203 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-3079
transform 1 0 3156 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-3080
transform 1 0 3059 0 1 1505
box 0 0 3 6
use FEEDTHRU  F-3081
transform 1 0 2995 0 1 1434
box 0 0 3 6
use FEEDTHRU  F-3082
transform 1 0 3306 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-3083
transform 1 0 3362 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-3084
transform 1 0 3311 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-3085
transform 1 0 3326 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-3086
transform 1 0 3325 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-3087
transform 1 0 3317 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-3088
transform 1 0 3327 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-3089
transform 1 0 3329 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-3090
transform 1 0 3513 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-3091
transform 1 0 3276 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-3092
transform 1 0 3407 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-3093
transform 1 0 3361 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-3094
transform 1 0 3492 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-3095
transform 1 0 3510 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-3096
transform 1 0 3501 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-3097
transform 1 0 3329 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-3098
transform 1 0 3371 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-3099
transform 1 0 3455 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-3100
transform 1 0 3462 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-3101
transform 1 0 3373 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-3102
transform 1 0 3307 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-3103
transform 1 0 3480 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-3104
transform 1 0 3299 0 1 1783
box 0 0 3 6
use FEEDTHRU  F-3105
transform 1 0 3312 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-3106
transform 1 0 3555 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-3107
transform 1 0 3371 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-3108
transform 1 0 3369 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-3109
transform 1 0 3365 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-3110
transform 1 0 3370 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-3111
transform 1 0 3368 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-3112
transform 1 0 3479 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-3113
transform 1 0 3389 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-3114
transform 1 0 3347 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-3115
transform 1 0 3519 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-3116
transform 1 0 3534 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-3117
transform 1 0 3516 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-3118
transform 1 0 3385 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-3119
transform 1 0 3073 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-3120
transform 1 0 3273 0 1 1630
box 0 0 3 6
use FEEDTHRU  F-3121
transform 1 0 3414 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-3122
transform 1 0 3464 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-3123
transform 1 0 3389 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-3124
transform 1 0 3404 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-3125
transform 1 0 3406 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-3126
transform 1 0 3310 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-3127
transform 1 0 3441 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-3128
transform 1 0 3456 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-3129
transform 1 0 3091 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-3130
transform 1 0 3161 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-3131
transform 1 0 3298 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-3132
transform 1 0 3372 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-3133
transform 1 0 3422 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-3134
transform 1 0 3347 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-3135
transform 1 0 3362 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-3136
transform 1 0 3364 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-3137
transform 1 0 3359 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-3138
transform 1 0 3429 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-3139
transform 1 0 3340 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-3140
transform 1 0 3426 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-3141
transform 1 0 3343 0 1 2667
box 0 0 3 6
use FEEDTHRU  F-3142
transform 1 0 3280 0 1 2454
box 0 0 3 6
use FEEDTHRU  F-3143
transform 1 0 3336 0 1 2211
box 0 0 3 6
use FEEDTHRU  F-3144
transform 1 0 3225 0 1 1990
box 0 0 3 6
use FEEDTHRU  F-3145
transform 1 0 3319 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-3146
transform 1 0 3311 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-3147
transform 1 0 3467 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-3148
transform 1 0 3245 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-3149
transform 1 0 3527 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-3150
transform 1 0 3434 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-3151
transform 1 0 3410 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-3152
transform 1 0 3360 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-3153
transform 1 0 3292 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-3154
transform 1 0 3143 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-3155
transform 1 0 3073 0 1 8653
box 0 0 3 6
use FEEDTHRU  F-3156
transform 1 0 3005 0 1 8734
box 0 0 3 6
use FEEDTHRU  F-3157
transform 1 0 3475 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-3158
transform 1 0 3286 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-3159
transform 1 0 3354 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-3160
transform 1 0 3404 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-3161
transform 1 0 3401 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-3162
transform 1 0 3411 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-3163
transform 1 0 3413 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-3164
transform 1 0 3597 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-3165
transform 1 0 3354 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-3166
transform 1 0 3488 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-3167
transform 1 0 3333 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-3168
transform 1 0 3335 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-3169
transform 1 0 3519 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-3170
transform 1 0 3270 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-3171
transform 1 0 3413 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-3172
transform 1 0 3373 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-3173
transform 1 0 3504 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-3174
transform 1 0 3522 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-3175
transform 1 0 3329 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-3176
transform 1 0 3337 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-3177
transform 1 0 3465 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-3178
transform 1 0 3334 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-3179
transform 1 0 3492 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-3180
transform 1 0 3477 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-3181
transform 1 0 3305 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-3182
transform 1 0 3347 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-3183
transform 1 0 3443 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-3184
transform 1 0 3438 0 1 2924
box 0 0 3 6
use FEEDTHRU  F-3185
transform 1 0 3091 0 1 8510
box 0 0 3 6
use FEEDTHRU  F-3186
transform 1 0 3241 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-3187
transform 1 0 3300 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-3188
transform 1 0 3356 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-3189
transform 1 0 3287 0 1 7632
box 0 0 3 6
use FEEDTHRU  F-3190
transform 1 0 3302 0 1 7389
box 0 0 3 6
use FEEDTHRU  F-3191
transform 1 0 3307 0 1 7096
box 0 0 3 6
use FEEDTHRU  F-3192
transform 1 0 3299 0 1 6821
box 0 0 3 6
use FEEDTHRU  F-3193
transform 1 0 3309 0 1 6554
box 0 0 3 6
use FEEDTHRU  F-3194
transform 1 0 3311 0 1 6261
box 0 0 3 6
use FEEDTHRU  F-3195
transform 1 0 3495 0 1 5920
box 0 0 3 6
use FEEDTHRU  F-3196
transform 1 0 3246 0 1 5617
box 0 0 3 6
use FEEDTHRU  F-3197
transform 1 0 3392 0 1 5318
box 0 0 3 6
use FEEDTHRU  F-3198
transform 1 0 3352 0 1 5009
box 0 0 3 6
use FEEDTHRU  F-3199
transform 1 0 3483 0 1 4658
box 0 0 3 6
use FEEDTHRU  F-3200
transform 1 0 3498 0 1 4345
box 0 0 3 6
use FEEDTHRU  F-3201
transform 1 0 3483 0 1 4068
box 0 0 3 6
use FEEDTHRU  F-3202
transform 1 0 3311 0 1 3775
box 0 0 3 6
use FEEDTHRU  F-3203
transform 1 0 3353 0 1 3452
box 0 0 3 6
use FEEDTHRU  F-3204
transform 1 0 3449 0 1 3153
box 0 0 3 6
use FEEDTHRU  F-3205
transform 1 0 3330 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-3206
transform 1 0 3386 0 1 7849
box 0 0 3 6
use FEEDTHRU  F-3207
transform 1 0 3336 0 1 8096
box 0 0 3 6
use FEEDTHRU  F-3208
transform 1 0 3271 0 1 8315
box 0 0 3 6
use FEEDTHRU  F-3209
transform 1 0 3122 0 1 8510
box 0 0 3 6
<< metal1 >>
rect 2941 1415 2964 1416
rect 2944 1417 3036 1418
rect 2947 1419 2954 1420
rect 2957 1419 2979 1420
rect 2960 1421 3000 1422
rect 2966 1423 3006 1424
rect 2984 1425 3003 1426
rect 2987 1427 2997 1428
rect 3011 1427 3015 1428
rect 3017 1427 3021 1428
rect 3026 1427 3033 1428
rect 3044 1427 3051 1428
rect 3047 1429 3060 1430
rect 3056 1431 3069 1432
rect 2809 1441 3243 1442
rect 2938 1443 2991 1444
rect 2944 1445 3115 1446
rect 2947 1447 2968 1448
rect 2953 1449 2981 1450
rect 2973 1451 3085 1452
rect 2978 1453 3031 1454
rect 2984 1455 3018 1456
rect 2987 1457 3103 1458
rect 2987 1459 3055 1460
rect 2993 1461 3175 1462
rect 2996 1463 3061 1464
rect 2999 1465 3064 1466
rect 3000 1467 3015 1468
rect 2950 1469 3016 1470
rect 3002 1471 3067 1472
rect 3005 1473 3070 1474
rect 3011 1475 3019 1476
rect 2963 1477 3013 1478
rect 2952 1479 2965 1480
rect 3023 1479 3088 1480
rect 3026 1481 3094 1482
rect 2931 1483 3028 1484
rect 3035 1483 3121 1484
rect 3036 1485 3130 1486
rect 3039 1487 3091 1488
rect 3044 1489 3112 1490
rect 3047 1491 3127 1492
rect 3056 1493 3145 1494
rect 3150 1493 3237 1494
rect 3153 1495 3184 1496
rect 3156 1497 3212 1498
rect 3165 1499 3226 1500
rect 3177 1501 3230 1502
rect 3190 1503 3198 1504
rect 3204 1503 3252 1504
rect 2920 1512 2987 1513
rect 2920 1514 2994 1515
rect 2936 1516 3125 1517
rect 2938 1518 3257 1519
rect 2934 1520 2940 1521
rect 2933 1522 2949 1523
rect 2917 1524 2949 1525
rect 2941 1526 3254 1527
rect 2955 1528 3002 1529
rect 2809 1530 2955 1531
rect 2957 1530 3064 1531
rect 2924 1532 3065 1533
rect 2960 1534 3077 1535
rect 2964 1536 2974 1537
rect 2970 1538 3008 1539
rect 2971 1540 3332 1541
rect 2990 1542 3059 1543
rect 3015 1544 3080 1545
rect 2967 1546 3017 1547
rect 3018 1546 3043 1547
rect 3025 1548 3031 1549
rect 3035 1548 3344 1549
rect 3046 1550 3161 1551
rect 3069 1552 3134 1553
rect 3072 1554 3094 1555
rect 2984 1556 3095 1557
rect 2917 1558 2984 1559
rect 3084 1558 3170 1559
rect 3087 1560 3182 1561
rect 3102 1562 3197 1563
rect 3111 1564 3278 1565
rect 3114 1566 3206 1567
rect 2931 1568 3116 1569
rect 2930 1570 3216 1571
rect 3120 1572 3212 1573
rect 3027 1574 3122 1575
rect 3126 1574 3230 1575
rect 3032 1576 3128 1577
rect 3129 1576 3347 1577
rect 2977 1578 3131 1579
rect 3141 1578 3203 1579
rect 3142 1580 3362 1581
rect 3144 1582 3400 1583
rect 3054 1584 3146 1585
rect 3150 1584 3356 1585
rect 3066 1586 3152 1587
rect 3153 1586 3359 1587
rect 2998 1588 3155 1589
rect 3156 1588 3284 1589
rect 3060 1590 3158 1591
rect 2902 1592 3062 1593
rect 3162 1592 3218 1593
rect 3165 1594 3272 1595
rect 3174 1596 3311 1597
rect 3175 1598 3379 1599
rect 3177 1600 3314 1601
rect 3178 1602 3194 1603
rect 3183 1604 3248 1605
rect 3090 1606 3185 1607
rect 3012 1608 3092 1609
rect 2974 1610 3014 1611
rect 3187 1610 3376 1611
rect 3222 1612 3326 1613
rect 3225 1614 3317 1615
rect 3236 1616 3329 1617
rect 3241 1618 3386 1619
rect 3259 1620 3418 1621
rect 3274 1622 3407 1623
rect 3295 1624 3435 1625
rect 3319 1626 3383 1627
rect 3322 1628 3404 1629
rect 2894 1637 3451 1638
rect 2917 1639 2942 1640
rect 2933 1641 2978 1642
rect 2932 1643 3146 1644
rect 2944 1645 2972 1646
rect 2930 1647 2972 1648
rect 2954 1649 3006 1650
rect 2948 1651 2954 1652
rect 2974 1651 3054 1652
rect 2881 1653 2975 1654
rect 2983 1653 3033 1654
rect 2990 1655 3139 1656
rect 3010 1657 3208 1658
rect 3011 1659 3161 1660
rect 3035 1661 3502 1662
rect 2986 1663 3036 1664
rect 2987 1665 3080 1666
rect 2929 1667 3081 1668
rect 3039 1669 3226 1670
rect 2922 1671 3039 1672
rect 3041 1671 3071 1672
rect 3007 1673 3072 1674
rect 3046 1675 3179 1676
rect 3049 1677 3145 1678
rect 2902 1679 3051 1680
rect 3058 1679 3106 1680
rect 3013 1681 3060 1682
rect 3001 1683 3015 1684
rect 3061 1683 3148 1684
rect 3016 1685 3063 1686
rect 3064 1685 3118 1686
rect 3083 1687 3449 1688
rect 3124 1689 3172 1690
rect 3076 1691 3124 1692
rect 2915 1693 3078 1694
rect 3130 1693 3214 1694
rect 3151 1695 3199 1696
rect 3089 1697 3151 1698
rect 3175 1697 3223 1698
rect 3127 1699 3175 1700
rect 3184 1699 3235 1700
rect 3190 1701 3353 1702
rect 3142 1703 3352 1704
rect 3094 1705 3142 1706
rect 3093 1707 3122 1708
rect 3193 1707 3359 1708
rect 3202 1709 3358 1710
rect 3154 1711 3202 1712
rect 3205 1711 3307 1712
rect 3157 1713 3205 1714
rect 3211 1713 3265 1714
rect 2998 1715 3211 1716
rect 3229 1715 3350 1716
rect 3181 1717 3229 1718
rect 3133 1719 3181 1720
rect 3091 1721 3133 1722
rect 3187 1721 3349 1722
rect 3025 1723 3187 1724
rect 2925 1725 3027 1726
rect 3231 1725 3361 1726
rect 3247 1727 3466 1728
rect 3196 1729 3247 1730
rect 3253 1729 3337 1730
rect 3256 1731 3340 1732
rect 3271 1733 3407 1734
rect 3270 1735 3372 1736
rect 3274 1737 3515 1738
rect 3283 1739 3385 1740
rect 3295 1741 3376 1742
rect 3217 1743 3295 1744
rect 3028 1745 3217 1746
rect 3300 1745 3418 1746
rect 3310 1747 3403 1748
rect 3313 1749 3406 1750
rect 3312 1751 3526 1752
rect 3316 1753 3472 1754
rect 3315 1755 3390 1756
rect 3319 1757 3421 1758
rect 3255 1759 3319 1760
rect 3322 1759 3424 1760
rect 3325 1761 3409 1762
rect 3241 1763 3325 1764
rect 3073 1765 3241 1766
rect 3331 1765 3433 1766
rect 3343 1767 3454 1768
rect 3259 1769 3343 1770
rect 3346 1769 3439 1770
rect 3355 1771 3457 1772
rect 3354 1773 3364 1774
rect 3372 1773 3411 1774
rect 3328 1775 3412 1776
rect 3378 1777 3460 1778
rect 3277 1779 3379 1780
rect 3276 1781 3393 1782
rect 3468 1781 3478 1782
rect 3552 1781 3573 1782
rect 2863 1790 2975 1791
rect 2866 1792 2871 1793
rect 2884 1792 2889 1793
rect 2894 1792 2933 1793
rect 2901 1794 3068 1795
rect 2904 1796 3051 1797
rect 2914 1798 3078 1799
rect 2918 1800 3124 1801
rect 2922 1802 3044 1803
rect 2925 1804 3042 1805
rect 2928 1806 3065 1807
rect 2953 1808 2999 1809
rect 2959 1810 3197 1811
rect 2962 1812 2988 1813
rect 2968 1814 3169 1815
rect 2971 1816 2996 1817
rect 2983 1818 3063 1819
rect 2990 1820 3133 1821
rect 2989 1822 3036 1823
rect 3007 1824 3039 1825
rect 3014 1826 3074 1827
rect 3026 1828 3056 1829
rect 3032 1830 3050 1831
rect 3005 1832 3032 1833
rect 3004 1834 3179 1835
rect 3034 1836 3172 1837
rect 3053 1838 3086 1839
rect 2941 1840 3053 1841
rect 2940 1842 3012 1843
rect 2977 1844 3011 1845
rect 2977 1846 3131 1847
rect 3059 1848 3092 1849
rect 3061 1850 3578 1851
rect 3080 1852 3101 1853
rect 3079 1854 3512 1855
rect 3089 1856 3214 1857
rect 3096 1858 3335 1859
rect 2917 1860 3098 1861
rect 3111 1860 3275 1861
rect 3136 1862 3226 1863
rect 2911 1864 3227 1865
rect 2910 1866 3071 1867
rect 3138 1866 3161 1867
rect 3141 1868 3164 1869
rect 2897 1870 3143 1871
rect 3144 1870 3185 1871
rect 2903 1872 3146 1873
rect 3166 1872 3217 1873
rect 3169 1874 3181 1875
rect 3174 1876 3215 1877
rect 3186 1878 3221 1879
rect 3190 1880 3202 1881
rect 3112 1882 3203 1883
rect 3204 1882 3239 1883
rect 3210 1884 3245 1885
rect 3222 1886 3263 1887
rect 3231 1888 3299 1889
rect 3198 1890 3233 1891
rect 3147 1892 3200 1893
rect 3117 1894 3149 1895
rect 2921 1896 3119 1897
rect 3234 1896 3269 1897
rect 3235 1898 3475 1899
rect 3240 1900 3287 1901
rect 3207 1902 3242 1903
rect 3109 1904 3209 1905
rect 3246 1904 3281 1905
rect 3150 1906 3248 1907
rect 3255 1906 3352 1907
rect 3264 1908 3545 1909
rect 3016 1910 3266 1911
rect 3270 1910 3305 1911
rect 3276 1912 3311 1913
rect 3294 1914 3329 1915
rect 3300 1916 3526 1917
rect 3114 1918 3302 1919
rect 3083 1920 3116 1921
rect 3306 1920 3353 1921
rect 3322 1922 3340 1923
rect 3312 1924 3341 1925
rect 3324 1926 3383 1927
rect 3336 1928 3416 1929
rect 3348 1930 3401 1931
rect 3354 1932 3431 1933
rect 3370 1934 3482 1935
rect 3384 1936 3566 1937
rect 3402 1938 3485 1939
rect 3318 1940 3404 1941
rect 3405 1940 3488 1941
rect 3408 1942 3491 1943
rect 3411 1944 3494 1945
rect 3412 1946 3548 1947
rect 3420 1948 3497 1949
rect 3375 1950 3422 1951
rect 2896 1952 3377 1953
rect 3423 1952 3500 1953
rect 3342 1954 3425 1955
rect 3315 1956 3344 1957
rect 3438 1956 3509 1957
rect 3448 1958 3647 1959
rect 3450 1960 3521 1961
rect 3372 1962 3452 1963
rect 3453 1962 3524 1963
rect 3378 1964 3455 1965
rect 3456 1964 3527 1965
rect 3459 1966 3530 1967
rect 3468 1968 3539 1969
rect 3471 1970 3542 1971
rect 3552 1970 3637 1971
rect 3418 1972 3552 1973
rect 3558 1972 3584 1973
rect 3228 1974 3559 1975
rect 2980 1976 3230 1977
rect 2980 1978 3106 1979
rect 3562 1978 3575 1979
rect 3572 1980 3634 1981
rect 3501 1982 3572 1983
rect 3432 1984 3503 1985
rect 3357 1986 3434 1987
rect 3358 1988 3604 1989
rect 2866 1997 3011 1998
rect 2896 1999 3176 2000
rect 2903 2001 2959 2002
rect 2870 2003 2958 2004
rect 2902 2005 3071 2006
rect 2909 2007 3035 2008
rect 2915 2009 3053 2010
rect 2921 2011 3065 2012
rect 2924 2013 3197 2014
rect 2934 2015 3056 2016
rect 2940 2017 3040 2018
rect 2961 2019 3248 2020
rect 2960 2021 3158 2022
rect 2963 2023 3074 2024
rect 2966 2025 2990 2026
rect 2968 2027 3284 2028
rect 2972 2029 2999 2030
rect 2977 2031 3200 2032
rect 2984 2033 3146 2034
rect 2995 2035 3003 2036
rect 3005 2035 3131 2036
rect 3016 2037 3068 2038
rect 3017 2039 3080 2040
rect 3020 2041 3242 2042
rect 3023 2043 3113 2044
rect 3025 2045 3239 2046
rect 3028 2047 3152 2048
rect 3033 2049 3290 2050
rect 3036 2051 3050 2052
rect 3043 2053 3055 2054
rect 3031 2055 3043 2056
rect 3030 2057 3296 2058
rect 3051 2059 3062 2060
rect 3070 2059 3086 2060
rect 3076 2061 3092 2062
rect 3100 2061 3122 2062
rect 3109 2063 3191 2064
rect 3118 2065 3131 2066
rect 3097 2067 3119 2068
rect 3124 2067 3149 2068
rect 3142 2069 3200 2070
rect 2931 2071 3143 2072
rect 3160 2071 3182 2072
rect 3166 2073 3434 2074
rect 3169 2075 3350 2076
rect 3169 2077 3455 2078
rect 3178 2079 3194 2080
rect 3115 2081 3179 2082
rect 3184 2081 3242 2082
rect 3163 2083 3185 2084
rect 3139 2085 3164 2086
rect 3187 2085 3404 2086
rect 3202 2087 3212 2088
rect 2900 2089 3203 2090
rect 3208 2089 3218 2090
rect 3226 2089 3338 2090
rect 3232 2091 3314 2092
rect 3235 2093 3317 2094
rect 3220 2095 3236 2096
rect 3244 2095 3278 2096
rect 3244 2097 3302 2098
rect 3250 2099 3275 2100
rect 3250 2101 3254 2102
rect 3253 2103 3299 2104
rect 3214 2105 3299 2106
rect 3256 2107 3431 2108
rect 3262 2109 3332 2110
rect 3265 2111 3347 2112
rect 3268 2113 3365 2114
rect 3286 2115 3320 2116
rect 3307 2117 3383 2118
rect 3280 2119 3383 2120
rect 3310 2121 3640 2122
rect 3322 2123 3389 2124
rect 3340 2125 3404 2126
rect 3229 2127 3341 2128
rect 3229 2129 3524 2130
rect 3343 2131 3410 2132
rect 3103 2133 3344 2134
rect 3352 2133 3536 2134
rect 3358 2135 3434 2136
rect 3328 2137 3359 2138
rect 3367 2137 3401 2138
rect 3376 2139 3428 2140
rect 3376 2141 3527 2142
rect 3379 2143 3530 2144
rect 3385 2145 3521 2146
rect 3400 2147 3413 2148
rect 3418 2147 3546 2148
rect 3418 2149 3549 2150
rect 3424 2151 3443 2152
rect 3439 2153 3497 2154
rect 3448 2155 3524 2156
rect 3415 2157 3449 2158
rect 3415 2159 3578 2160
rect 3445 2161 3579 2162
rect 3481 2163 3671 2164
rect 3484 2165 3497 2166
rect 3451 2167 3485 2168
rect 3451 2169 3619 2170
rect 3490 2171 3533 2172
rect 3421 2173 3491 2174
rect 3370 2175 3422 2176
rect 3304 2177 3371 2178
rect 3493 2177 3536 2178
rect 3493 2179 3640 2180
rect 3499 2181 3566 2182
rect 3487 2183 3500 2184
rect 3502 2183 3527 2184
rect 3508 2185 3530 2186
rect 3514 2187 3654 2188
rect 3520 2189 3665 2190
rect 3538 2191 3559 2192
rect 3325 2193 3539 2194
rect 3555 2193 3613 2194
rect 3561 2195 3568 2196
rect 3541 2197 3562 2198
rect 3265 2199 3542 2200
rect 3571 2199 3604 2200
rect 3574 2201 3607 2202
rect 3583 2203 3610 2204
rect 3591 2205 3655 2206
rect 3633 2207 3649 2208
rect 3636 2209 3652 2210
rect 2902 2218 3131 2219
rect 2915 2220 3040 2221
rect 2924 2222 3074 2223
rect 2923 2224 3047 2225
rect 2927 2226 3228 2227
rect 2927 2228 3119 2229
rect 2934 2230 3249 2231
rect 2933 2232 2958 2233
rect 2961 2232 2985 2233
rect 2964 2234 3203 2235
rect 2966 2236 3041 2237
rect 2972 2238 2980 2239
rect 2985 2238 3284 2239
rect 2988 2240 3113 2241
rect 2993 2242 3093 2243
rect 2992 2244 3037 2245
rect 2920 2246 3038 2247
rect 3004 2248 3312 2249
rect 3007 2250 3101 2251
rect 3020 2252 3096 2253
rect 3017 2254 3020 2255
rect 3002 2256 3017 2257
rect 3023 2256 3317 2257
rect 3030 2258 3278 2259
rect 3031 2260 3055 2261
rect 3042 2262 3050 2263
rect 3043 2264 3052 2265
rect 2906 2266 3053 2267
rect 2906 2268 3200 2269
rect 2967 2270 3201 2271
rect 3060 2272 3347 2273
rect 3061 2274 3071 2275
rect 3067 2276 3251 2277
rect 3067 2278 3077 2279
rect 3076 2280 3122 2281
rect 2995 2282 3123 2283
rect 3079 2284 3314 2285
rect 3098 2286 3549 2287
rect 3103 2288 3194 2289
rect 2902 2290 3105 2291
rect 3116 2290 3125 2291
rect 3128 2290 3152 2291
rect 3140 2292 3176 2293
rect 3142 2294 3147 2295
rect 3143 2296 3179 2297
rect 3157 2298 3162 2299
rect 3169 2298 3531 2299
rect 3173 2300 3368 2301
rect 3176 2302 3306 2303
rect 3179 2304 3182 2305
rect 3182 2306 3185 2307
rect 3187 2306 3273 2307
rect 3197 2308 3242 2309
rect 3203 2310 3212 2311
rect 3163 2312 3213 2313
rect 3209 2314 3218 2315
rect 3215 2316 3299 2317
rect 3229 2318 3527 2319
rect 3233 2320 3245 2321
rect 3239 2322 3290 2323
rect 3245 2324 3296 2325
rect 3251 2326 3350 2327
rect 3256 2328 3288 2329
rect 3088 2330 3258 2331
rect 3089 2332 3236 2333
rect 3236 2334 3254 2335
rect 3263 2334 3320 2335
rect 3265 2336 3540 2337
rect 3275 2338 3332 2339
rect 3281 2340 3338 2341
rect 3284 2342 3341 2343
rect 3290 2344 3580 2345
rect 3296 2346 3359 2347
rect 3302 2348 3365 2349
rect 3307 2350 3321 2351
rect 3325 2350 3480 2351
rect 3326 2352 3383 2353
rect 3332 2354 3568 2355
rect 3338 2356 3389 2357
rect 3343 2358 3556 2359
rect 3350 2360 3577 2361
rect 3353 2362 3404 2363
rect 3359 2364 3410 2365
rect 3365 2366 3416 2367
rect 3370 2368 3556 2369
rect 3371 2370 3422 2371
rect 3379 2372 3542 2373
rect 3383 2374 3434 2375
rect 3385 2376 3528 2377
rect 3392 2378 3546 2379
rect 3400 2380 3586 2381
rect 3401 2382 3452 2383
rect 3057 2384 3453 2385
rect 3437 2386 3485 2387
rect 3439 2388 3587 2389
rect 3442 2390 3459 2391
rect 3445 2392 3543 2393
rect 3448 2394 3546 2395
rect 3418 2396 3450 2397
rect 3455 2396 3584 2397
rect 3473 2398 3494 2399
rect 3476 2400 3582 2401
rect 3481 2402 3678 2403
rect 3485 2404 3521 2405
rect 3490 2406 3644 2407
rect 3503 2408 3562 2409
rect 3509 2410 3568 2411
rect 3514 2412 3662 2413
rect 3521 2414 3533 2415
rect 3523 2416 3665 2417
rect 3524 2418 3536 2419
rect 3376 2420 3537 2421
rect 3377 2422 3428 2423
rect 3533 2422 3630 2423
rect 3558 2424 3618 2425
rect 3314 2426 3559 2427
rect 3564 2426 3615 2427
rect 3571 2428 3675 2429
rect 3488 2430 3674 2431
rect 3573 2432 3664 2433
rect 3603 2434 3621 2435
rect 3602 2436 3655 2437
rect 3606 2438 3624 2439
rect 3591 2440 3606 2441
rect 3609 2440 3626 2441
rect 3608 2442 3652 2443
rect 3425 2444 3651 2445
rect 3612 2446 3658 2447
rect 3611 2448 3627 2449
rect 3636 2448 3671 2449
rect 3308 2450 3637 2451
rect 3648 2450 3654 2451
rect 3413 2452 3648 2453
rect 2894 2461 3107 2462
rect 2899 2463 2934 2464
rect 2901 2465 3279 2466
rect 2904 2467 3110 2468
rect 2906 2469 3231 2470
rect 2913 2471 3059 2472
rect 2916 2473 3074 2474
rect 2918 2475 3077 2476
rect 2934 2477 3047 2478
rect 2943 2479 3243 2480
rect 2951 2481 2989 2482
rect 2955 2483 3029 2484
rect 2992 2485 3117 2486
rect 2995 2487 3324 2488
rect 3010 2489 3294 2490
rect 3013 2491 3180 2492
rect 3016 2493 3077 2494
rect 3019 2495 3035 2496
rect 3022 2497 3255 2498
rect 3037 2499 3071 2500
rect 3043 2501 3080 2502
rect 3052 2503 3119 2504
rect 3061 2505 3065 2506
rect 2974 2507 3062 2508
rect 3095 2507 3131 2508
rect 3094 2509 3393 2510
rect 3101 2511 3228 2512
rect 3104 2513 3165 2514
rect 3049 2515 3104 2516
rect 3128 2515 3195 2516
rect 3092 2517 3128 2518
rect 3146 2517 3207 2518
rect 3152 2519 3237 2520
rect 3091 2521 3237 2522
rect 3158 2523 3213 2524
rect 3161 2525 3225 2526
rect 3170 2527 3201 2528
rect 3140 2529 3201 2530
rect 3140 2531 3363 2532
rect 3188 2533 3306 2534
rect 3212 2535 3273 2536
rect 3197 2537 3273 2538
rect 3182 2539 3198 2540
rect 3233 2539 3577 2540
rect 2964 2541 3234 2542
rect 3248 2541 3261 2542
rect 3266 2541 3288 2542
rect 3281 2543 3345 2544
rect 2927 2545 3282 2546
rect 3284 2545 3348 2546
rect 3203 2547 3285 2548
rect 3143 2549 3204 2550
rect 3143 2551 3252 2552
rect 3296 2551 3556 2552
rect 3215 2553 3297 2554
rect 3302 2553 3369 2554
rect 3086 2555 3303 2556
rect 3067 2557 3086 2558
rect 3308 2557 3375 2558
rect 3257 2559 3309 2560
rect 3314 2559 3387 2560
rect 3239 2561 3315 2562
rect 3320 2561 3381 2562
rect 3245 2563 3321 2564
rect 3031 2565 3246 2566
rect 3326 2565 3393 2566
rect 2985 2567 3327 2568
rect 2961 2569 2987 2570
rect 3332 2569 3399 2570
rect 3290 2571 3333 2572
rect 3209 2573 3291 2574
rect 3004 2575 3210 2576
rect 3004 2577 3041 2578
rect 3338 2577 3411 2578
rect 3263 2579 3339 2580
rect 3350 2579 3693 2580
rect 3275 2581 3351 2582
rect 2915 2583 3276 2584
rect 3353 2583 3483 2584
rect 3356 2585 3552 2586
rect 3365 2587 3432 2588
rect 3371 2589 3444 2590
rect 3176 2591 3372 2592
rect 3122 2593 3177 2594
rect 2979 2595 3122 2596
rect 3401 2595 3468 2596
rect 3416 2597 3420 2598
rect 3422 2597 3662 2598
rect 3425 2599 3668 2600
rect 3359 2601 3426 2602
rect 3452 2601 3594 2602
rect 3458 2603 3507 2604
rect 3479 2605 3516 2606
rect 3449 2607 3480 2608
rect 3485 2607 3552 2608
rect 3413 2609 3486 2610
rect 3488 2609 3555 2610
rect 3497 2611 3612 2612
rect 3500 2613 3609 2614
rect 3509 2615 3558 2616
rect 3437 2617 3510 2618
rect 3521 2617 3579 2618
rect 3524 2619 3582 2620
rect 3527 2621 3564 2622
rect 3533 2623 3657 2624
rect 3545 2625 3568 2626
rect 3503 2627 3546 2628
rect 3455 2629 3504 2630
rect 3383 2631 3456 2632
rect 3530 2631 3567 2632
rect 3569 2631 3587 2632
rect 3536 2633 3588 2634
rect 3573 2635 3638 2636
rect 3377 2637 3573 2638
rect 3311 2639 3378 2640
rect 3575 2639 3744 2640
rect 3584 2641 3591 2642
rect 3539 2643 3591 2644
rect 3473 2645 3540 2646
rect 3599 2645 3651 2646
rect 3605 2647 3656 2648
rect 3329 2649 3606 2650
rect 3617 2649 3680 2650
rect 3404 2651 3618 2652
rect 3620 2651 3665 2652
rect 3623 2653 3648 2654
rect 3542 2655 3625 2656
rect 3476 2657 3543 2658
rect 3653 2657 3696 2658
rect 3602 2659 3653 2660
rect 3602 2661 3641 2662
rect 3670 2661 3690 2662
rect 3677 2663 3734 2664
rect 3614 2665 3677 2666
rect 2890 2674 3201 2675
rect 2897 2676 3110 2677
rect 2905 2678 3134 2679
rect 2915 2680 3007 2681
rect 2931 2682 3071 2683
rect 2934 2684 3282 2685
rect 2908 2686 3281 2687
rect 2937 2688 2968 2689
rect 2941 2690 3207 2691
rect 2944 2692 3269 2693
rect 2943 2694 2949 2695
rect 2946 2696 3210 2697
rect 2965 2698 3434 2699
rect 2974 2700 3198 2701
rect 2976 2702 3195 2703
rect 2986 2704 3019 2705
rect 2997 2706 3213 2707
rect 3004 2708 3359 2709
rect 3028 2710 3056 2711
rect 3027 2712 3159 2713
rect 3034 2714 3050 2715
rect 3036 2716 3065 2717
rect 3046 2718 3303 2719
rect 3061 2720 3089 2721
rect 3073 2722 3246 2723
rect 3076 2724 3113 2725
rect 3079 2726 3098 2727
rect 3079 2728 3110 2729
rect 3082 2730 3315 2731
rect 3085 2732 3092 2733
rect 3058 2734 3086 2735
rect 3094 2734 3137 2735
rect 3103 2736 3149 2737
rect 3103 2738 3461 2739
rect 3106 2740 3122 2741
rect 3106 2742 3267 2743
rect 3115 2744 3128 2745
rect 3124 2746 3309 2747
rect 3140 2748 3618 2749
rect 3151 2750 3189 2751
rect 3022 2752 3188 2753
rect 3164 2754 3182 2755
rect 3170 2756 3206 2757
rect 3176 2758 3194 2759
rect 3199 2758 3567 2759
rect 3217 2760 3255 2761
rect 3224 2762 3245 2763
rect 2979 2764 3224 2765
rect 3230 2764 3299 2765
rect 3229 2766 3516 2767
rect 3233 2768 3302 2769
rect 3236 2770 3251 2771
rect 3203 2772 3236 2773
rect 3238 2772 3591 2773
rect 3242 2774 3287 2775
rect 3256 2776 3327 2777
rect 3262 2778 3405 2779
rect 3275 2780 3326 2781
rect 3260 2782 3275 2783
rect 3259 2784 3330 2785
rect 2969 2786 3329 2787
rect 3284 2788 3317 2789
rect 3293 2790 3335 2791
rect 3292 2792 3588 2793
rect 3296 2794 3311 2795
rect 3323 2794 3395 2795
rect 3272 2796 3323 2797
rect 3332 2796 3621 2797
rect 3290 2798 3332 2799
rect 2915 2800 3290 2801
rect 3344 2800 3428 2801
rect 3356 2802 3688 2803
rect 3278 2804 3356 2805
rect 3368 2804 3452 2805
rect 3367 2806 3662 2807
rect 3374 2808 3464 2809
rect 3362 2810 3374 2811
rect 3380 2810 3404 2811
rect 2950 2812 3380 2813
rect 3386 2812 3458 2813
rect 3160 2814 3386 2815
rect 3398 2814 3488 2815
rect 3397 2816 3606 2817
rect 3410 2818 3663 2819
rect 3409 2820 3755 2821
rect 3425 2822 3518 2823
rect 3431 2824 3524 2825
rect 3347 2826 3431 2827
rect 3439 2826 3673 2827
rect 3443 2828 3494 2829
rect 2972 2830 3443 2831
rect 3455 2830 3548 2831
rect 3371 2832 3455 2833
rect 3467 2832 3560 2833
rect 3377 2834 3467 2835
rect 3475 2834 3625 2835
rect 3479 2836 3692 2837
rect 3482 2838 3659 2839
rect 3392 2840 3482 2841
rect 3320 2842 3392 2843
rect 3415 2842 3659 2843
rect 3490 2844 3564 2845
rect 3496 2846 3504 2847
rect 3499 2848 3558 2849
rect 3506 2850 3641 2851
rect 3505 2852 3632 2853
rect 3509 2854 3596 2855
rect 3422 2856 3509 2857
rect 3350 2858 3422 2859
rect 2922 2860 3350 2861
rect 3526 2860 3685 2861
rect 3529 2862 3573 2863
rect 3485 2864 3572 2865
rect 3532 2866 3570 2867
rect 3535 2868 3546 2869
rect 3539 2870 3608 2871
rect 3542 2872 3611 2873
rect 3541 2874 3683 2875
rect 3551 2876 3626 2877
rect 3554 2878 3629 2879
rect 3565 2880 3582 2881
rect 3575 2882 3769 2883
rect 3578 2884 3641 2885
rect 3589 2886 3600 2887
rect 3592 2888 3603 2889
rect 3652 2888 3682 2889
rect 3655 2890 3719 2891
rect 3338 2892 3656 2893
rect 3039 2894 3338 2895
rect 3676 2894 3713 2895
rect 3679 2896 3716 2897
rect 3584 2898 3679 2899
rect 3583 2900 3668 2901
rect 3689 2900 3759 2901
rect 3695 2902 3739 2903
rect 3708 2904 3727 2905
rect 3637 2906 3710 2907
rect 3637 2908 3699 2909
rect 3664 2910 3698 2911
rect 3361 2912 3666 2913
rect 3729 2912 3737 2913
rect 3601 2914 3736 2915
rect 3675 2916 3729 2917
rect 3733 2916 3787 2917
rect 3740 2918 3748 2919
rect 3700 2920 3748 2921
rect 3741 2922 3773 2923
rect 2914 2931 3086 2932
rect 2931 2933 3287 2934
rect 2950 2935 3364 2936
rect 2953 2937 3359 2938
rect 2962 2939 3074 2940
rect 2934 2941 3073 2942
rect 2921 2943 2934 2944
rect 2961 2943 2995 2944
rect 2971 2945 3428 2946
rect 2976 2947 3194 2948
rect 2993 2949 3469 2950
rect 3006 2951 3030 2952
rect 3014 2953 3245 2954
rect 3018 2955 3024 2956
rect 3027 2955 3188 2956
rect 3043 2957 3422 2958
rect 3045 2959 3163 2960
rect 3055 2961 3061 2962
rect 3069 2961 3104 2962
rect 3079 2963 3304 2964
rect 2979 2965 3079 2966
rect 2978 2967 3380 2968
rect 3097 2969 3100 2970
rect 3096 2971 3113 2972
rect 3091 2973 3112 2974
rect 3106 2975 3260 2976
rect 3109 2977 3124 2978
rect 3115 2979 3145 2980
rect 3126 2981 3149 2982
rect 3118 2983 3148 2984
rect 3117 2985 3476 2986
rect 3130 2987 3139 2988
rect 3121 2989 3130 2990
rect 3120 2991 3379 2992
rect 3133 2993 3142 2994
rect 3151 2993 3175 2994
rect 3157 2995 3239 2996
rect 3160 2997 3374 2998
rect 3181 2999 3187 3000
rect 3180 3001 3443 3002
rect 3210 3003 3224 3004
rect 3222 3005 3230 3006
rect 3228 3007 3251 3008
rect 2899 3009 3250 3010
rect 3237 3011 3766 3012
rect 3240 3013 3263 3014
rect 3246 3015 3257 3016
rect 3255 3017 3275 3018
rect 3261 3019 3659 3020
rect 3268 3021 3274 3022
rect 3267 3023 3311 3024
rect 3038 3025 3310 3026
rect 3280 3027 3286 3028
rect 3279 3029 3317 3030
rect 3292 3031 3358 3032
rect 3291 3033 3299 3034
rect 2975 3035 3298 3036
rect 3294 3037 3302 3038
rect 3312 3037 3431 3038
rect 3315 3039 3332 3040
rect 3318 3041 3335 3042
rect 3325 3043 3370 3044
rect 2943 3045 3325 3046
rect 3333 3045 3338 3046
rect 3349 3045 3352 3046
rect 3372 3045 3686 3046
rect 3403 3047 3661 3048
rect 3397 3049 3403 3050
rect 2912 3051 3397 3052
rect 2911 3053 3085 3054
rect 3409 3053 3421 3054
rect 3367 3055 3409 3056
rect 2965 3057 3367 3058
rect 2964 3059 3206 3060
rect 3415 3059 3427 3060
rect 3439 3059 3445 3060
rect 3361 3061 3439 3062
rect 3454 3061 3484 3062
rect 2946 3063 3454 3064
rect 3466 3063 3472 3064
rect 3460 3065 3466 3066
rect 3499 3065 3757 3066
rect 3505 3067 3511 3068
rect 3493 3069 3505 3070
rect 3487 3071 3493 3072
rect 3481 3073 3487 3074
rect 3082 3075 3481 3076
rect 3508 3075 3514 3076
rect 3496 3077 3508 3078
rect 3490 3079 3496 3080
rect 3535 3079 3729 3080
rect 3523 3081 3535 3082
rect 3517 3083 3523 3084
rect 3433 3085 3517 3086
rect 3432 3087 3452 3088
rect 3450 3089 3670 3090
rect 3541 3091 3688 3092
rect 3526 3093 3541 3094
rect 3543 3093 3692 3094
rect 3585 3095 3704 3096
rect 3589 3097 3622 3098
rect 3571 3099 3589 3100
rect 3559 3101 3571 3102
rect 3547 3103 3559 3104
rect 3529 3105 3547 3106
rect 3528 3107 3728 3108
rect 3595 3109 3616 3110
rect 3610 3111 3631 3112
rect 3612 3113 3797 3114
rect 3625 3115 3792 3116
rect 3592 3117 3625 3118
rect 3628 3117 3794 3118
rect 3607 3119 3628 3120
rect 3565 3121 3607 3122
rect 3637 3121 3747 3122
rect 3640 3123 3646 3124
rect 3657 3123 3750 3124
rect 3669 3125 3780 3126
rect 3601 3127 3779 3128
rect 3583 3129 3601 3130
rect 3532 3131 3583 3132
rect 3678 3131 3719 3132
rect 3681 3133 3704 3134
rect 3700 3135 3719 3136
rect 3694 3137 3701 3138
rect 3706 3137 3795 3138
rect 3709 3139 3722 3140
rect 3738 3139 3763 3140
rect 3712 3141 3738 3142
rect 3741 3141 3766 3142
rect 3715 3143 3741 3144
rect 3697 3145 3716 3146
rect 3675 3147 3698 3148
rect 3772 3147 3790 3148
rect 3743 3149 3772 3150
rect 3788 3149 3809 3150
rect 3797 3151 3802 3152
rect 3824 3151 3832 3152
rect 2906 3160 3070 3161
rect 2909 3162 3130 3163
rect 2913 3164 3142 3165
rect 2916 3166 3076 3167
rect 2933 3168 2950 3169
rect 2935 3170 3259 3171
rect 2945 3172 3030 3173
rect 2944 3174 3322 3175
rect 2951 3176 3364 3177
rect 2958 3178 3370 3179
rect 2961 3180 3313 3181
rect 2968 3182 2981 3183
rect 2968 3184 3310 3185
rect 2977 3186 3502 3187
rect 2984 3188 3157 3189
rect 2987 3190 3145 3191
rect 2993 3192 3003 3193
rect 3014 3192 3106 3193
rect 3014 3194 3024 3195
rect 3020 3196 3307 3197
rect 3023 3198 3415 3199
rect 3030 3200 3469 3201
rect 3033 3202 3049 3203
rect 3042 3204 3169 3205
rect 3045 3206 3472 3207
rect 3051 3208 3061 3209
rect 3057 3210 3728 3211
rect 3063 3212 3073 3213
rect 3078 3212 3340 3213
rect 3084 3214 3103 3215
rect 3087 3216 3106 3217
rect 3093 3218 3097 3219
rect 2911 3220 3097 3221
rect 3099 3220 3115 3221
rect 3108 3222 3118 3223
rect 3111 3224 3130 3225
rect 3123 3226 3166 3227
rect 3123 3228 3151 3229
rect 3138 3230 3142 3231
rect 3174 3230 3430 3231
rect 3162 3232 3175 3233
rect 3066 3234 3163 3235
rect 3201 3234 3277 3235
rect 3207 3236 3325 3237
rect 3213 3238 3238 3239
rect 3147 3240 3238 3241
rect 3222 3242 3634 3243
rect 3243 3244 3295 3245
rect 3255 3246 3301 3247
rect 3264 3248 3286 3249
rect 3267 3250 3343 3251
rect 3270 3252 3274 3253
rect 3273 3254 3289 3255
rect 3282 3256 3355 3257
rect 3288 3258 3352 3259
rect 3294 3260 3328 3261
rect 3297 3262 3337 3263
rect 3303 3264 3331 3265
rect 3312 3266 3367 3267
rect 3279 3268 3367 3269
rect 3318 3270 3382 3271
rect 3120 3272 3319 3273
rect 3120 3274 3127 3275
rect 3324 3274 3397 3275
rect 3252 3276 3397 3277
rect 3348 3278 3445 3279
rect 3354 3280 3451 3281
rect 3360 3282 3391 3283
rect 3372 3284 3757 3285
rect 3372 3286 3457 3287
rect 3375 3288 3713 3289
rect 3378 3290 3661 3291
rect 3315 3292 3379 3293
rect 2961 3294 3316 3295
rect 3390 3294 3481 3295
rect 3393 3296 3424 3297
rect 3402 3298 3689 3299
rect 3402 3300 3487 3301
rect 3408 3302 3658 3303
rect 3333 3304 3409 3305
rect 3426 3304 3682 3305
rect 3027 3306 3427 3307
rect 3435 3306 3529 3307
rect 3441 3308 3463 3309
rect 3459 3310 3535 3311
rect 3240 3312 3535 3313
rect 3240 3314 3292 3315
rect 2921 3316 3292 3317
rect 2920 3318 3484 3319
rect 3471 3320 3541 3321
rect 3477 3322 3798 3323
rect 3483 3324 3707 3325
rect 3489 3326 3571 3327
rect 3492 3328 3724 3329
rect 3504 3330 3710 3331
rect 3246 3332 3505 3333
rect 3210 3334 3247 3335
rect 3210 3336 3235 3337
rect 3234 3338 3786 3339
rect 3507 3340 3643 3341
rect 3507 3342 3547 3343
rect 3513 3344 3686 3345
rect 3216 3346 3514 3347
rect 3516 3346 3649 3347
rect 3522 3348 3785 3349
rect 3525 3350 3613 3351
rect 3420 3352 3613 3353
rect 3228 3354 3421 3355
rect 3228 3356 3250 3357
rect 3540 3356 3601 3357
rect 3552 3358 3586 3359
rect 3564 3360 3898 3361
rect 3570 3362 3628 3363
rect 3573 3364 3631 3365
rect 3465 3366 3631 3367
rect 3465 3368 3781 3369
rect 3576 3370 3828 3371
rect 3582 3372 3688 3373
rect 3582 3374 3792 3375
rect 3594 3376 3607 3377
rect 3621 3376 3694 3377
rect 3645 3378 3661 3379
rect 3438 3380 3646 3381
rect 3666 3380 3670 3381
rect 3669 3382 3747 3383
rect 3192 3384 3748 3385
rect 3186 3386 3193 3387
rect 3180 3388 3187 3389
rect 2964 3390 3181 3391
rect 2965 3392 3205 3393
rect 3681 3392 3766 3393
rect 3690 3394 3767 3395
rect 3697 3396 3733 3397
rect 3624 3398 3697 3399
rect 3543 3400 3625 3401
rect 3700 3400 3736 3401
rect 3495 3402 3700 3403
rect 3261 3404 3496 3405
rect 3705 3404 3722 3405
rect 3715 3406 3845 3407
rect 3678 3408 3715 3409
rect 3737 3408 3791 3409
rect 3703 3410 3739 3411
rect 3195 3412 3703 3413
rect 3743 3412 3797 3413
rect 3357 3414 3745 3415
rect 3357 3416 3454 3417
rect 3384 3418 3454 3419
rect 3384 3420 3433 3421
rect 3432 3422 3511 3423
rect 3750 3422 3842 3423
rect 3752 3424 3795 3425
rect 3718 3426 3754 3427
rect 3717 3428 3852 3429
rect 3740 3430 3794 3431
rect 3741 3432 3867 3433
rect 3762 3434 3864 3435
rect 3768 3436 3818 3437
rect 3788 3438 3855 3439
rect 3588 3440 3788 3441
rect 3804 3440 3888 3441
rect 3811 3442 3877 3443
rect 3815 3444 3858 3445
rect 3771 3446 3815 3447
rect 3831 3446 3839 3447
rect 3558 3448 3831 3449
rect 3558 3450 3616 3451
rect 3860 3450 3881 3451
rect 2815 3459 2823 3460
rect 2878 3459 3220 3460
rect 2884 3461 3217 3462
rect 2899 3463 3085 3464
rect 2908 3465 3103 3466
rect 2913 3467 3070 3468
rect 2916 3469 3064 3470
rect 2915 3471 3076 3472
rect 2918 3473 3283 3474
rect 2920 3475 3292 3476
rect 2935 3477 3265 3478
rect 2939 3479 3205 3480
rect 2942 3481 3130 3482
rect 2949 3483 2955 3484
rect 2958 3483 2973 3484
rect 2961 3485 3268 3486
rect 2965 3487 3331 3488
rect 2968 3489 3337 3490
rect 2978 3491 3316 3492
rect 2980 3493 3325 3494
rect 2987 3495 3163 3496
rect 2990 3497 3358 3498
rect 2993 3499 3316 3500
rect 3008 3501 3015 3502
rect 3014 3503 3028 3504
rect 3033 3503 3076 3504
rect 3039 3505 3094 3506
rect 3042 3507 3169 3508
rect 3048 3509 3097 3510
rect 3051 3511 3061 3512
rect 3051 3513 3106 3514
rect 3054 3515 3253 3516
rect 3057 3517 3139 3518
rect 3066 3519 3115 3520
rect 3072 3521 3121 3522
rect 3081 3523 3142 3524
rect 3087 3525 3208 3526
rect 3114 3527 3157 3528
rect 3120 3529 3181 3530
rect 3036 3531 3181 3532
rect 3126 3533 3166 3534
rect 3126 3535 3187 3536
rect 3132 3537 3193 3538
rect 2960 3539 3193 3540
rect 3144 3541 3235 3542
rect 2947 3543 3235 3544
rect 3147 3545 3238 3546
rect 3156 3547 3211 3548
rect 3159 3549 3214 3550
rect 3168 3551 3247 3552
rect 2891 3553 3247 3554
rect 3186 3555 3241 3556
rect 3189 3557 3244 3558
rect 3198 3559 3427 3560
rect 3198 3561 3421 3562
rect 3020 3563 3421 3564
rect 3201 3565 3451 3566
rect 3204 3567 3259 3568
rect 3222 3569 3271 3570
rect 3225 3571 3274 3572
rect 3240 3573 3295 3574
rect 3249 3575 3289 3576
rect 3252 3577 3301 3578
rect 3255 3579 3433 3580
rect 3258 3581 3343 3582
rect 3264 3583 3313 3584
rect 3270 3585 3409 3586
rect 3276 3587 3767 3588
rect 3276 3589 3319 3590
rect 3023 3591 3319 3592
rect 3279 3593 3340 3594
rect 3282 3595 3367 3596
rect 3174 3597 3367 3598
rect 3174 3599 3229 3600
rect 3228 3601 3307 3602
rect 3288 3603 3379 3604
rect 3291 3605 3382 3606
rect 3294 3607 3361 3608
rect 3300 3609 3415 3610
rect 3306 3611 3349 3612
rect 3312 3613 3355 3614
rect 3321 3615 3424 3616
rect 3324 3617 3364 3618
rect 3330 3619 3373 3620
rect 3348 3621 3391 3622
rect 3354 3623 3397 3624
rect 3369 3625 3376 3626
rect 3378 3625 3454 3626
rect 3384 3627 3454 3628
rect 3150 3629 3385 3630
rect 2956 3631 3151 3632
rect 3390 3631 3724 3632
rect 3396 3633 3460 3634
rect 3402 3635 3721 3636
rect 3408 3637 3778 3638
rect 3414 3639 3505 3640
rect 3417 3641 3502 3642
rect 3426 3643 3490 3644
rect 3429 3645 3749 3646
rect 3432 3647 3478 3648
rect 3435 3649 3895 3650
rect 3444 3651 3508 3652
rect 3456 3653 3553 3654
rect 3465 3655 3788 3656
rect 3468 3657 3541 3658
rect 3471 3659 3781 3660
rect 3474 3661 3526 3662
rect 3483 3663 3724 3664
rect 3489 3665 3559 3666
rect 3045 3667 3559 3668
rect 3495 3669 3532 3670
rect 3501 3671 3577 3672
rect 3507 3673 3571 3674
rect 3510 3675 3574 3676
rect 3513 3677 3568 3678
rect 3513 3679 3595 3680
rect 3441 3681 3595 3682
rect 3519 3683 3583 3684
rect 3525 3685 3764 3686
rect 3534 3687 3592 3688
rect 3537 3689 3858 3690
rect 3543 3691 3898 3692
rect 3549 3693 3822 3694
rect 3561 3695 3625 3696
rect 3573 3697 3613 3698
rect 3579 3699 3757 3700
rect 3585 3701 3760 3702
rect 3597 3703 3754 3704
rect 3600 3705 3836 3706
rect 3615 3707 3661 3708
rect 3621 3709 3700 3710
rect 3387 3711 3700 3712
rect 3624 3713 3703 3714
rect 3627 3715 3670 3716
rect 3630 3717 3745 3718
rect 3645 3719 3756 3720
rect 3645 3721 3706 3722
rect 3651 3723 3753 3724
rect 3666 3725 3858 3726
rect 3648 3727 3667 3728
rect 3642 3729 3649 3730
rect 3672 3729 3688 3730
rect 3675 3731 3691 3732
rect 3684 3733 3694 3734
rect 3687 3735 3697 3736
rect 3633 3737 3697 3738
rect 3633 3739 3682 3740
rect 3702 3739 3715 3740
rect 3705 3741 3718 3742
rect 3720 3741 3739 3742
rect 3654 3743 3739 3744
rect 3726 3745 3733 3746
rect 3741 3745 3843 3746
rect 3660 3747 3742 3748
rect 3750 3747 3874 3748
rect 3770 3749 3852 3750
rect 3778 3751 3832 3752
rect 3784 3753 3791 3754
rect 3787 3755 3794 3756
rect 3790 3757 3797 3758
rect 3796 3759 3864 3760
rect 3799 3761 3869 3762
rect 3808 3763 3815 3764
rect 3735 3765 3815 3766
rect 3811 3767 3818 3768
rect 3729 3769 3818 3770
rect 3838 3769 3849 3770
rect 3848 3771 3855 3772
rect 3860 3771 3888 3772
rect 3564 3773 3862 3774
rect 2881 3782 3220 3783
rect 2893 3784 3247 3785
rect 2904 3786 3362 3787
rect 2908 3788 3431 3789
rect 2915 3790 2927 3791
rect 2942 3790 3239 3791
rect 2946 3792 2958 3793
rect 2949 3794 3347 3795
rect 2960 3796 3199 3797
rect 2963 3798 3009 3799
rect 2918 3800 3009 3801
rect 2953 3802 2965 3803
rect 2953 3804 3190 3805
rect 2967 3806 3413 3807
rect 2972 3808 2991 3809
rect 2971 3810 3280 3811
rect 2884 3812 3281 3813
rect 2978 3814 2997 3815
rect 2978 3816 3164 3817
rect 2981 3818 3133 3819
rect 3014 3820 3383 3821
rect 3017 3822 3437 3823
rect 2950 3824 3018 3825
rect 3036 3824 3322 3825
rect 3039 3826 3131 3827
rect 3038 3828 3316 3829
rect 3042 3830 3473 3831
rect 3045 3832 3325 3833
rect 3048 3834 3059 3835
rect 3048 3836 3311 3837
rect 3060 3838 3065 3839
rect 3066 3838 3071 3839
rect 3081 3838 3107 3839
rect 3084 3840 3365 3841
rect 3112 3842 3139 3843
rect 3114 3844 3119 3845
rect 3120 3844 3191 3845
rect 3124 3846 3649 3847
rect 3126 3848 3488 3849
rect 3139 3850 3367 3851
rect 3144 3852 3233 3853
rect 3156 3854 3275 3855
rect 2922 3856 3158 3857
rect 3168 3856 3245 3857
rect 3174 3858 3299 3859
rect 3072 3860 3176 3861
rect 3180 3860 3185 3861
rect 3186 3860 3329 3861
rect 3204 3862 3335 3863
rect 3208 3864 3568 3865
rect 3222 3866 3317 3867
rect 3223 3868 3625 3869
rect 3225 3870 3338 3871
rect 3150 3872 3227 3873
rect 3228 3872 3263 3873
rect 3234 3874 3305 3875
rect 3240 3876 3368 3877
rect 3087 3878 3242 3879
rect 3075 3880 3089 3881
rect 3054 3882 3077 3883
rect 3055 3884 3440 3885
rect 3256 3886 3481 3887
rect 3258 3888 3341 3889
rect 3264 3890 3395 3891
rect 3276 3892 3407 3893
rect 3282 3894 3374 3895
rect 3159 3896 3284 3897
rect 3286 3896 3301 3897
rect 3288 3898 3756 3899
rect 3291 3900 3377 3901
rect 3252 3902 3293 3903
rect 3294 3902 3443 3903
rect 3306 3904 3479 3905
rect 3312 3906 3485 3907
rect 3318 3908 3323 3909
rect 3369 3908 3506 3909
rect 3378 3910 3449 3911
rect 3249 3912 3380 3913
rect 3250 3914 3532 3915
rect 3384 3916 3404 3917
rect 3387 3918 3401 3919
rect 3390 3920 3554 3921
rect 3396 3922 3548 3923
rect 3408 3924 3763 3925
rect 2939 3926 3410 3927
rect 2929 3928 2939 3929
rect 3417 3928 3425 3929
rect 3418 3930 3586 3931
rect 3420 3932 3467 3933
rect 3444 3934 3572 3935
rect 3033 3936 3446 3937
rect 3032 3938 3148 3939
rect 3450 3938 3524 3939
rect 3456 3940 3590 3941
rect 3468 3942 3614 3943
rect 3469 3944 3622 3945
rect 3474 3946 3944 3947
rect 3489 3948 3638 3949
rect 3453 3950 3491 3951
rect 3454 3952 3709 3953
rect 3496 3954 3655 3955
rect 3501 3956 3620 3957
rect 3330 3958 3503 3959
rect 2897 3960 3332 3961
rect 2896 3962 3217 3963
rect 3507 3962 3650 3963
rect 3354 3964 3509 3965
rect 3510 3964 3897 3965
rect 3414 3966 3512 3967
rect 3267 3968 3416 3969
rect 3192 3970 3269 3971
rect 3513 3970 3656 3971
rect 3525 3972 3883 3973
rect 3526 3974 3732 3975
rect 3529 3976 3595 3977
rect 3532 3978 3661 3979
rect 3519 3980 3662 3981
rect 3348 3982 3521 3983
rect 3270 3984 3350 3985
rect 3537 3984 3916 3985
rect 3538 3986 3735 3987
rect 3541 3988 3559 3989
rect 3543 3990 3919 3991
rect 3549 3992 3771 3993
rect 3555 3994 3592 3995
rect 3559 3996 3843 3997
rect 3561 3998 3632 3999
rect 3573 4000 3578 4001
rect 3579 4000 3712 4001
rect 3580 4002 3753 4003
rect 3597 4004 3765 4005
rect 3600 4006 3626 4007
rect 3432 4008 3602 4009
rect 3051 4010 3434 4011
rect 3607 4010 3676 4011
rect 3627 4012 3869 4013
rect 3633 4014 3744 4015
rect 3643 4016 3862 4017
rect 3645 4018 3774 4019
rect 3651 4020 3822 4021
rect 3426 4022 3653 4023
rect 3666 4022 3742 4023
rect 3667 4024 3947 4025
rect 3670 4026 3886 4027
rect 3684 4028 3692 4029
rect 3694 4030 3858 4031
rect 3705 4032 3753 4033
rect 3615 4034 3707 4035
rect 3720 4034 3777 4035
rect 3721 4036 3767 4037
rect 3726 4038 3818 4039
rect 3696 4040 3728 4041
rect 3729 4040 3768 4041
rect 3737 4042 3788 4043
rect 3748 4044 3760 4045
rect 3460 4046 3759 4047
rect 3702 4048 3750 4049
rect 3761 4048 3890 4049
rect 3778 4050 3815 4051
rect 3723 4052 3780 4053
rect 3784 4052 3863 4053
rect 3790 4054 3839 4055
rect 3796 4056 3845 4057
rect 3808 4058 3857 4059
rect 3718 4060 3809 4061
rect 3811 4060 3860 4061
rect 3672 4062 3812 4063
rect 3820 4062 3832 4063
rect 3848 4062 3903 4063
rect 3799 4064 3848 4065
rect 3851 4064 3906 4065
rect 3865 4066 3879 4067
rect 3925 4066 3930 4067
rect 2809 4075 3176 4076
rect 2887 4077 3281 4078
rect 2907 4079 3059 4080
rect 2918 4081 3434 4082
rect 2922 4083 3431 4084
rect 2926 4085 3458 4086
rect 2925 4087 3395 4088
rect 2928 4089 3392 4090
rect 2935 4091 3317 4092
rect 2941 4093 3299 4094
rect 2944 4095 3386 4096
rect 2947 4097 3287 4098
rect 2954 4099 3347 4100
rect 2961 4101 3191 4102
rect 2971 4103 3431 4104
rect 2981 4105 3488 4106
rect 2984 4107 2991 4108
rect 2996 4107 3740 4108
rect 2996 4109 3173 4110
rect 3026 4111 3033 4112
rect 3038 4111 3473 4112
rect 3041 4113 3437 4114
rect 3042 4115 3383 4116
rect 3045 4117 3065 4118
rect 2899 4119 3046 4120
rect 3048 4119 3293 4120
rect 2896 4121 3293 4122
rect 3052 4123 3404 4124
rect 2903 4125 3052 4126
rect 3057 4125 3311 4126
rect 3076 4127 3082 4128
rect 3070 4129 3076 4130
rect 3088 4129 3094 4130
rect 3112 4129 3133 4130
rect 3111 4131 3148 4132
rect 3124 4133 3518 4134
rect 3151 4135 3488 4136
rect 3154 4137 3287 4138
rect 3160 4139 3164 4140
rect 3178 4139 3185 4140
rect 2958 4141 3185 4142
rect 3190 4141 3524 4142
rect 3196 4143 3212 4144
rect 3202 4145 3410 4146
rect 3214 4147 3233 4148
rect 3220 4149 3227 4150
rect 3014 4151 3227 4152
rect 3229 4151 3440 4152
rect 3232 4153 3239 4154
rect 3238 4155 3245 4156
rect 3208 4157 3245 4158
rect 3208 4159 3425 4160
rect 3250 4161 3728 4162
rect 3256 4163 3317 4164
rect 3256 4165 3263 4166
rect 3262 4167 3275 4168
rect 3265 4169 3284 4170
rect 3268 4171 3275 4172
rect 2950 4173 3269 4174
rect 3280 4173 3323 4174
rect 3298 4175 3305 4176
rect 2910 4177 3305 4178
rect 3310 4177 3335 4178
rect 3223 4179 3335 4180
rect 3322 4181 3329 4182
rect 2951 4183 3329 4184
rect 3325 4185 3332 4186
rect 3337 4185 3353 4186
rect 2906 4187 3338 4188
rect 3340 4187 3344 4188
rect 3355 4187 3368 4188
rect 3349 4189 3368 4190
rect 2938 4191 3350 4192
rect 3373 4191 3398 4192
rect 3379 4193 3395 4194
rect 3403 4193 3497 4194
rect 3406 4195 3428 4196
rect 3412 4197 3422 4198
rect 3415 4199 3425 4200
rect 3169 4201 3416 4202
rect 3433 4201 3467 4202
rect 3439 4203 3443 4204
rect 3442 4205 3446 4206
rect 3448 4205 3735 4206
rect 3451 4207 3461 4208
rect 3241 4209 3461 4210
rect 3454 4211 3464 4212
rect 3466 4211 3470 4212
rect 3475 4211 3527 4212
rect 3478 4213 3494 4214
rect 3481 4215 3491 4216
rect 3484 4217 3500 4218
rect 3505 4217 3527 4218
rect 3505 4219 3530 4220
rect 3508 4221 3530 4222
rect 3508 4223 3798 4224
rect 3520 4225 3536 4226
rect 3400 4227 3521 4228
rect 3376 4229 3401 4230
rect 3532 4229 3710 4230
rect 3511 4231 3533 4232
rect 3502 4233 3512 4234
rect 2975 4235 3503 4236
rect 3538 4235 3783 4236
rect 3032 4237 3539 4238
rect 3541 4237 3563 4238
rect 3547 4239 3569 4240
rect 3547 4241 3802 4242
rect 3418 4243 3801 4244
rect 3553 4245 3575 4246
rect 3553 4247 3578 4248
rect 3571 4249 3587 4250
rect 3577 4251 3581 4252
rect 3559 4253 3581 4254
rect 3559 4255 3817 4256
rect 3589 4257 3599 4258
rect 3601 4257 3617 4258
rect 3604 4259 3653 4260
rect 3607 4261 3611 4262
rect 3613 4261 3629 4262
rect 3619 4263 3623 4264
rect 3625 4263 3635 4264
rect 3631 4265 3756 4266
rect 3637 4267 3653 4268
rect 3643 4269 3659 4270
rect 3646 4271 3650 4272
rect 3655 4271 3665 4272
rect 3667 4271 3686 4272
rect 3682 4273 3942 4274
rect 3694 4275 3713 4276
rect 3694 4277 3872 4278
rect 3706 4279 3725 4280
rect 3691 4281 3707 4282
rect 3721 4281 3809 4282
rect 3721 4283 3916 4284
rect 3731 4285 3827 4286
rect 3743 4287 3923 4288
rect 3749 4289 3759 4290
rect 3749 4291 3952 4292
rect 3767 4293 3789 4294
rect 3773 4295 3795 4296
rect 3776 4297 3875 4298
rect 3761 4299 3777 4300
rect 3752 4301 3762 4302
rect 3779 4301 3909 4302
rect 3764 4303 3780 4304
rect 3782 4303 3928 4304
rect 3785 4305 3793 4306
rect 3770 4307 3792 4308
rect 3688 4309 3771 4310
rect 3661 4311 3689 4312
rect 3785 4311 3932 4312
rect 3814 4313 3890 4314
rect 3670 4315 3889 4316
rect 3670 4317 3900 4318
rect 3820 4319 3836 4320
rect 3523 4321 3820 4322
rect 3838 4321 3872 4322
rect 3844 4323 3869 4324
rect 3847 4325 3851 4326
rect 3847 4327 3919 4328
rect 3853 4329 3866 4330
rect 3856 4331 3866 4332
rect 3737 4333 3857 4334
rect 3859 4333 3869 4334
rect 3862 4335 3879 4336
rect 3882 4335 3925 4336
rect 3898 4337 3937 4338
rect 3905 4339 3908 4340
rect 3902 4341 3905 4342
rect 3901 4343 3918 4344
rect 2882 4352 2992 4353
rect 2890 4354 3263 4355
rect 2896 4356 3323 4357
rect 2899 4358 2922 4359
rect 2906 4360 3365 4361
rect 2909 4362 3341 4363
rect 2925 4364 2973 4365
rect 2924 4366 3407 4367
rect 2928 4368 3386 4369
rect 2932 4370 3293 4371
rect 2933 4372 3311 4373
rect 2947 4374 3350 4375
rect 2954 4376 3239 4377
rect 2957 4378 3428 4379
rect 2961 4380 3332 4381
rect 2961 4382 3494 4383
rect 2964 4384 3182 4385
rect 2973 4386 2985 4387
rect 2975 4388 3212 4389
rect 2979 4390 2997 4391
rect 2994 4392 3266 4393
rect 2876 4394 3266 4395
rect 2997 4396 3009 4397
rect 2872 4398 3010 4399
rect 3003 4400 3227 4401
rect 3017 4402 3503 4403
rect 3018 4404 3027 4405
rect 3024 4406 3257 4407
rect 3032 4408 3422 4409
rect 3035 4410 3584 4411
rect 2943 4412 3037 4413
rect 3045 4412 3049 4413
rect 3051 4412 3055 4413
rect 3057 4412 3503 4413
rect 3057 4414 3326 4415
rect 3075 4416 3079 4417
rect 3090 4416 3094 4417
rect 3096 4416 3112 4417
rect 3105 4418 3109 4419
rect 3117 4418 3121 4419
rect 3126 4418 3133 4419
rect 3132 4420 3161 4421
rect 3135 4422 3815 4423
rect 3138 4424 3935 4425
rect 3139 4426 3197 4427
rect 2892 4428 3197 4429
rect 3142 4430 3200 4431
rect 3144 4432 3218 4433
rect 3129 4434 3146 4435
rect 3151 4434 3817 4435
rect 3154 4436 3482 4437
rect 3166 4438 3191 4439
rect 3178 4440 3191 4441
rect 3157 4442 3179 4443
rect 3157 4444 3311 4445
rect 3184 4446 3206 4447
rect 3214 4446 3254 4447
rect 3220 4448 3236 4449
rect 3223 4450 3245 4451
rect 3229 4452 3410 4453
rect 3202 4454 3230 4455
rect 3232 4454 3242 4455
rect 3247 4454 3317 4455
rect 3262 4456 3335 4457
rect 3274 4458 3293 4459
rect 3274 4460 3281 4461
rect 3268 4462 3281 4463
rect 3147 4464 3269 4465
rect 3295 4464 3431 4465
rect 3304 4466 3317 4467
rect 3298 4468 3305 4469
rect 3322 4468 3404 4469
rect 3334 4470 3344 4471
rect 3337 4472 3347 4473
rect 3355 4472 3371 4473
rect 3358 4474 3362 4475
rect 3081 4476 3362 4477
rect 3081 4478 3353 4479
rect 3352 4480 3368 4481
rect 3364 4482 3434 4483
rect 3367 4484 3467 4485
rect 2947 4486 3467 4487
rect 3382 4488 3392 4489
rect 3385 4490 3395 4491
rect 3388 4492 3398 4493
rect 3391 4494 3401 4495
rect 3042 4496 3401 4497
rect 3412 4496 3521 4497
rect 3415 4498 3419 4499
rect 3424 4498 3470 4499
rect 3424 4500 3509 4501
rect 3430 4502 3440 4503
rect 3433 4504 3443 4505
rect 3442 4506 3458 4507
rect 3445 4508 3461 4509
rect 3451 4510 3455 4511
rect 3460 4510 3762 4511
rect 3463 4512 3740 4513
rect 3472 4514 3476 4515
rect 3478 4514 3506 4515
rect 3481 4516 3752 4517
rect 3484 4518 3500 4519
rect 3487 4520 3744 4521
rect 3487 4522 3530 4523
rect 3490 4524 3533 4525
rect 3493 4526 3512 4527
rect 3499 4528 3518 4529
rect 3505 4530 3524 4531
rect 3508 4532 3527 4533
rect 3511 4534 3548 4535
rect 3517 4536 3536 4537
rect 3520 4538 3539 4539
rect 3523 4540 3805 4541
rect 3529 4542 3771 4543
rect 3532 4544 3710 4545
rect 3535 4546 3563 4547
rect 3541 4548 3569 4549
rect 3547 4550 3575 4551
rect 3553 4552 3822 4553
rect 3553 4554 3886 4555
rect 3556 4556 3578 4557
rect 3559 4558 3798 4559
rect 3559 4560 3872 4561
rect 3565 4562 3581 4563
rect 3571 4564 3587 4565
rect 3589 4564 3599 4565
rect 3595 4566 3623 4567
rect 3601 4568 3605 4569
rect 3613 4568 3629 4569
rect 3616 4570 3918 4571
rect 3625 4572 3665 4573
rect 3631 4574 3936 4575
rect 3634 4576 3833 4577
rect 3643 4578 3647 4579
rect 3649 4578 3653 4579
rect 3655 4578 3659 4579
rect 3667 4578 3689 4579
rect 3673 4580 3962 4581
rect 3682 4582 3954 4583
rect 3682 4584 3939 4585
rect 3685 4586 3942 4587
rect 3685 4588 3695 4589
rect 3691 4590 3887 4591
rect 3697 4592 3713 4593
rect 3703 4594 3719 4595
rect 3706 4596 3774 4597
rect 3610 4598 3707 4599
rect 3709 4598 3925 4599
rect 3721 4600 3827 4601
rect 3715 4602 3826 4603
rect 3733 4604 3750 4605
rect 3754 4604 3759 4605
rect 3757 4606 3879 4607
rect 3760 4608 3777 4609
rect 3577 4610 3776 4611
rect 3766 4612 3783 4613
rect 3769 4614 3921 4615
rect 3779 4616 3875 4617
rect 3791 4618 3890 4619
rect 3790 4620 3928 4621
rect 3785 4622 3929 4623
rect 3784 4624 3795 4625
rect 3793 4626 3824 4627
rect 3805 4628 3975 4629
rect 3808 4630 3943 4631
rect 3811 4632 3829 4633
rect 3835 4632 3845 4633
rect 3856 4632 3860 4633
rect 3853 4634 3857 4635
rect 3670 4636 3854 4637
rect 3865 4636 3881 4637
rect 3868 4638 3884 4639
rect 3874 4640 3949 4641
rect 3661 4642 3950 4643
rect 3877 4644 3946 4645
rect 3898 4646 3914 4647
rect 3901 4648 3917 4649
rect 3850 4650 3901 4651
rect 3847 4652 3851 4653
rect 3904 4652 3920 4653
rect 3724 4654 3904 4655
rect 3907 4654 3923 4655
rect 3763 4656 3908 4657
rect 3951 4656 3978 4657
rect 2876 4665 3010 4666
rect 2869 4667 2877 4668
rect 2872 4669 3010 4670
rect 2885 4671 2995 4672
rect 2892 4673 3347 4674
rect 2896 4675 3197 4676
rect 2899 4677 3317 4678
rect 2903 4679 2919 4680
rect 2906 4681 3279 4682
rect 2912 4683 3261 4684
rect 2926 4685 3049 4686
rect 2936 4687 3236 4688
rect 2936 4689 3082 4690
rect 2940 4691 2951 4692
rect 2943 4693 3332 4694
rect 2947 4695 3167 4696
rect 2959 4697 3386 4698
rect 2961 4699 3542 4700
rect 2964 4701 3644 4702
rect 2973 4703 3046 4704
rect 2991 4705 3013 4706
rect 2979 4707 2992 4708
rect 3003 4707 3222 4708
rect 3018 4709 3022 4710
rect 3024 4709 3300 4710
rect 3044 4711 3165 4712
rect 3047 4713 3055 4714
rect 3057 4713 3150 4714
rect 3065 4715 3362 4716
rect 3071 4717 3509 4718
rect 3078 4719 3081 4720
rect 3077 4721 3146 4722
rect 2903 4723 3147 4724
rect 3083 4725 3109 4726
rect 3090 4727 3108 4728
rect 3122 4727 3182 4728
rect 2933 4729 3183 4730
rect 3135 4731 3218 4732
rect 3120 4733 3135 4734
rect 3119 4735 3179 4736
rect 3139 4737 3521 4738
rect 3126 4739 3141 4740
rect 3096 4741 3126 4742
rect 3154 4741 3491 4742
rect 3158 4743 3206 4744
rect 3170 4745 3434 4746
rect 3176 4747 3242 4748
rect 3188 4749 3230 4750
rect 3190 4751 3198 4752
rect 3194 4753 3266 4754
rect 3036 4755 3267 4756
rect 3037 4757 3345 4758
rect 3203 4759 3281 4760
rect 3209 4761 3254 4762
rect 3215 4763 3293 4764
rect 3027 4765 3294 4766
rect 3027 4767 3287 4768
rect 3223 4769 3459 4770
rect 3230 4771 3503 4772
rect 3233 4773 3305 4774
rect 2957 4775 3306 4776
rect 3245 4777 3341 4778
rect 3247 4779 3381 4780
rect 3251 4781 3335 4782
rect 3257 4783 3359 4784
rect 3268 4785 3773 4786
rect 3269 4787 3353 4788
rect 3274 4789 3751 4790
rect 3275 4791 3383 4792
rect 3281 4793 3371 4794
rect 3132 4795 3372 4796
rect 2886 4797 3132 4798
rect 3295 4797 3309 4798
rect 3302 4799 3392 4800
rect 3310 4801 3399 4802
rect 3311 4803 3443 4804
rect 3314 4805 3446 4806
rect 3317 4807 3407 4808
rect 3320 4809 3410 4810
rect 3322 4811 3600 4812
rect 3199 4813 3324 4814
rect 3335 4813 3467 4814
rect 3338 4815 3470 4816
rect 3341 4817 3431 4818
rect 3347 4819 3413 4820
rect 3353 4821 3485 4822
rect 3356 4823 3419 4824
rect 3362 4825 3494 4826
rect 3374 4827 3506 4828
rect 3377 4829 3773 4830
rect 3386 4831 3518 4832
rect 3388 4833 3740 4834
rect 3142 4835 3390 4836
rect 3404 4835 3672 4836
rect 3416 4837 3425 4838
rect 3422 4839 3554 4840
rect 3428 4841 3473 4842
rect 3431 4843 3482 4844
rect 3434 4845 3536 4846
rect 3446 4847 3455 4848
rect 3452 4849 3897 4850
rect 3460 4851 3700 4852
rect 3464 4853 3584 4854
rect 3476 4855 3940 4856
rect 3482 4857 3572 4858
rect 3494 4859 3590 4860
rect 3506 4861 3596 4862
rect 3523 4863 3776 4864
rect 3524 4865 3632 4866
rect 3532 4867 3660 4868
rect 3536 4869 3650 4870
rect 3542 4871 3656 4872
rect 3529 4873 3657 4874
rect 3530 4875 3626 4876
rect 3547 4877 3597 4878
rect 3548 4879 3662 4880
rect 3554 4881 3674 4882
rect 3556 4883 3594 4884
rect 3367 4885 3558 4886
rect 3368 4887 3500 4888
rect 3500 4889 3560 4890
rect 3262 4891 3561 4892
rect 3263 4893 3329 4894
rect 3329 4895 3401 4896
rect 3401 4897 3488 4898
rect 3488 4899 3602 4900
rect 3563 4901 3668 4902
rect 3364 4903 3669 4904
rect 3565 4905 3783 4906
rect 3569 4907 3854 4908
rect 3577 4909 3894 4910
rect 3587 4911 3686 4912
rect 3605 4913 3710 4914
rect 3478 4915 3709 4916
rect 3611 4917 3776 4918
rect 3623 4919 3961 4920
rect 3629 4921 3734 4922
rect 3632 4923 3770 4924
rect 3511 4925 3769 4926
rect 3512 4927 3614 4928
rect 3638 4927 3698 4928
rect 3644 4929 3901 4930
rect 3581 4931 3900 4932
rect 3662 4933 3704 4934
rect 3665 4935 3707 4936
rect 3678 4937 3847 4938
rect 3682 4939 3933 4940
rect 3691 4941 3840 4942
rect 3693 4943 3984 4944
rect 3696 4945 3755 4946
rect 3702 4947 3929 4948
rect 3715 4949 3833 4950
rect 3714 4951 3761 4952
rect 3717 4953 3904 4954
rect 3726 4955 3767 4956
rect 3419 4957 3766 4958
rect 3738 4959 3788 4960
rect 3741 4961 3791 4962
rect 3744 4963 3864 4964
rect 3757 4965 3829 4966
rect 3759 4967 3923 4968
rect 3763 4969 3836 4970
rect 3762 4971 3794 4972
rect 3779 4973 3887 4974
rect 3797 4975 3894 4976
rect 3800 4977 3903 4978
rect 3803 4979 3845 4980
rect 3805 4981 3910 4982
rect 3808 4983 3971 4984
rect 3809 4985 3857 4986
rect 3812 4987 3860 4988
rect 3821 4989 3875 4990
rect 3824 4991 3878 4992
rect 3833 4993 3881 4994
rect 3836 4995 3884 4996
rect 3729 4997 3883 4998
rect 3850 4999 3897 5000
rect 3866 5001 3914 5002
rect 3784 5003 3913 5004
rect 3747 5005 3786 5006
rect 3869 5005 3917 5006
rect 3889 5007 3920 5008
rect 3935 5007 3968 5008
rect 2863 5016 2877 5017
rect 2870 5018 3010 5019
rect 2873 5020 3048 5021
rect 2879 5022 3195 5023
rect 2882 5024 3013 5025
rect 2896 5026 3132 5027
rect 2905 5028 3276 5029
rect 2912 5030 3147 5031
rect 2922 5032 3150 5033
rect 2922 5034 3279 5035
rect 2919 5036 3280 5037
rect 2929 5038 3336 5039
rect 2933 5040 3070 5041
rect 2940 5042 3312 5043
rect 2941 5044 2951 5045
rect 2947 5046 3264 5047
rect 2960 5048 3387 5049
rect 2973 5050 3222 5051
rect 2972 5052 3193 5053
rect 2988 5054 2992 5055
rect 2994 5054 2998 5055
rect 3000 5054 3309 5055
rect 3003 5056 3318 5057
rect 3006 5058 3028 5059
rect 3012 5060 3022 5061
rect 3021 5062 3126 5063
rect 3037 5064 3165 5065
rect 3041 5066 3141 5067
rect 2893 5068 3142 5069
rect 3018 5070 3043 5071
rect 3044 5070 3072 5071
rect 3048 5072 3108 5073
rect 3057 5074 3270 5075
rect 2979 5076 3271 5077
rect 3060 5078 3066 5079
rect 3066 5080 3081 5081
rect 3077 5082 3115 5083
rect 3078 5084 3084 5085
rect 3102 5084 3135 5085
rect 3119 5086 3130 5087
rect 3122 5088 3133 5089
rect 3156 5088 3171 5089
rect 3158 5090 3163 5091
rect 3168 5090 3198 5091
rect 3180 5092 3183 5093
rect 3183 5094 3267 5095
rect 3198 5096 3459 5097
rect 3203 5098 3241 5099
rect 3108 5100 3205 5101
rect 3219 5100 3321 5101
rect 3222 5102 3372 5103
rect 3227 5104 3373 5105
rect 3231 5106 3561 5107
rect 3233 5108 3274 5109
rect 3030 5110 3235 5111
rect 3030 5112 3097 5113
rect 3243 5112 3315 5113
rect 3245 5114 3676 5115
rect 3246 5116 3381 5117
rect 3249 5118 3390 5119
rect 3251 5120 3292 5121
rect 3215 5122 3253 5123
rect 3209 5124 3217 5125
rect 3176 5126 3211 5127
rect 3257 5126 3310 5127
rect 3260 5128 3313 5129
rect 3281 5130 3322 5131
rect 2919 5132 3283 5133
rect 3297 5132 3405 5133
rect 3299 5134 3316 5135
rect 3300 5136 3558 5137
rect 3302 5138 3319 5139
rect 3293 5140 3304 5141
rect 3323 5140 3723 5141
rect 3324 5142 3339 5143
rect 3327 5144 3600 5145
rect 3333 5146 3447 5147
rect 3339 5148 3348 5149
rect 3188 5150 3349 5151
rect 3344 5152 3361 5153
rect 3305 5154 3346 5155
rect 3351 5154 3357 5155
rect 3329 5156 3358 5157
rect 3353 5158 3394 5159
rect 3362 5160 3409 5161
rect 3363 5162 3660 5163
rect 3368 5164 3679 5165
rect 3369 5166 3432 5167
rect 3374 5168 3415 5169
rect 3381 5170 3612 5171
rect 3387 5172 3783 5173
rect 3398 5174 3433 5175
rect 3401 5176 3430 5177
rect 3416 5178 3637 5179
rect 3377 5180 3418 5181
rect 3419 5180 3427 5181
rect 3420 5182 3818 5183
rect 3434 5184 3460 5185
rect 3438 5186 3776 5187
rect 3447 5188 3709 5189
rect 3450 5190 3657 5191
rect 3468 5192 3843 5193
rect 3471 5194 3666 5195
rect 3480 5196 3663 5197
rect 3488 5198 3520 5199
rect 3489 5200 3712 5201
rect 3435 5202 3712 5203
rect 3530 5204 3780 5205
rect 3512 5206 3532 5207
rect 3542 5206 3562 5207
rect 3543 5208 3839 5209
rect 3554 5210 3586 5211
rect 3536 5212 3556 5213
rect 3537 5214 3639 5215
rect 3563 5216 3580 5217
rect 3581 5216 3769 5217
rect 3587 5218 3688 5219
rect 3593 5220 3672 5221
rect 3569 5222 3595 5223
rect 3612 5222 3748 5223
rect 3623 5224 3903 5225
rect 3605 5226 3625 5227
rect 3629 5226 3649 5227
rect 3632 5228 3876 5229
rect 3642 5230 3703 5231
rect 3657 5232 3715 5233
rect 3422 5234 3716 5235
rect 3660 5236 3832 5237
rect 3669 5238 3727 5239
rect 3672 5240 3730 5241
rect 3500 5242 3730 5243
rect 3464 5244 3502 5245
rect 3465 5246 3597 5247
rect 3675 5246 3697 5247
rect 3678 5248 3733 5249
rect 3681 5250 3745 5251
rect 3684 5252 3742 5253
rect 3693 5254 3913 5255
rect 3699 5256 3773 5257
rect 3702 5258 3760 5259
rect 3705 5260 3763 5261
rect 3717 5262 3864 5263
rect 3441 5264 3719 5265
rect 3725 5264 3807 5265
rect 3735 5266 3786 5267
rect 3738 5268 3854 5269
rect 3747 5270 3798 5271
rect 3644 5272 3797 5273
rect 3750 5274 3801 5275
rect 3588 5276 3800 5277
rect 3753 5278 3870 5279
rect 3759 5280 3804 5281
rect 3567 5282 3804 5283
rect 3765 5284 3822 5285
rect 3630 5286 3821 5287
rect 3771 5288 3810 5289
rect 3476 5290 3811 5291
rect 3477 5292 3483 5293
rect 3452 5294 3484 5295
rect 3453 5296 3495 5297
rect 3495 5298 3507 5299
rect 3507 5300 3857 5301
rect 3774 5302 3847 5303
rect 3756 5304 3846 5305
rect 3783 5306 3834 5307
rect 3786 5308 3837 5309
rect 3812 5310 3850 5311
rect 3341 5312 3814 5313
rect 3824 5312 3897 5313
rect 3827 5314 3867 5315
rect 3834 5316 3890 5317
rect 2884 5325 3271 5326
rect 2888 5327 3142 5328
rect 2891 5329 2896 5330
rect 2908 5329 3211 5330
rect 2912 5331 2923 5332
rect 2911 5333 3130 5334
rect 2929 5335 2935 5336
rect 2941 5335 3212 5336
rect 2945 5337 3181 5338
rect 2965 5339 3230 5340
rect 2969 5341 3043 5342
rect 2972 5343 3349 5344
rect 2975 5345 3103 5346
rect 2979 5347 3766 5348
rect 2984 5349 2989 5350
rect 2990 5349 2995 5350
rect 2996 5349 3049 5350
rect 2999 5351 3043 5352
rect 3003 5353 3382 5354
rect 3008 5355 3013 5356
rect 3018 5355 3319 5356
rect 3021 5357 3269 5358
rect 3020 5359 3115 5360
rect 3023 5361 3097 5362
rect 3030 5363 3361 5364
rect 3030 5365 3188 5366
rect 3036 5367 3061 5368
rect 3048 5369 3067 5370
rect 3054 5371 3386 5372
rect 3054 5373 3079 5374
rect 3069 5375 3209 5376
rect 3072 5377 3287 5378
rect 3075 5379 3418 5380
rect 3099 5381 3401 5382
rect 3106 5383 3176 5384
rect 3111 5385 3370 5386
rect 3115 5387 3205 5388
rect 2922 5389 3206 5390
rect 3121 5391 3163 5392
rect 3132 5393 3179 5394
rect 3144 5395 3358 5396
rect 3145 5397 3169 5398
rect 3147 5399 3782 5400
rect 3151 5401 3241 5402
rect 2960 5403 3242 5404
rect 3154 5405 3244 5406
rect 3160 5407 3220 5408
rect 3163 5409 3253 5410
rect 3169 5411 3280 5412
rect 3172 5413 3283 5414
rect 3057 5415 3284 5416
rect 3181 5417 3310 5418
rect 3156 5419 3311 5420
rect 3157 5421 3217 5422
rect 3183 5423 3215 5424
rect 3184 5425 3313 5426
rect 3192 5427 3245 5428
rect 3193 5429 3235 5430
rect 3217 5431 3322 5432
rect 3220 5433 3325 5434
rect 3226 5435 3515 5436
rect 3235 5437 3346 5438
rect 3246 5439 3320 5440
rect 3247 5441 3394 5442
rect 3249 5443 3398 5444
rect 3033 5445 3251 5446
rect 3253 5445 3292 5446
rect 3259 5447 3304 5448
rect 3265 5449 3316 5450
rect 3271 5451 3415 5452
rect 3277 5453 3409 5454
rect 3289 5455 3334 5456
rect 3295 5457 3430 5458
rect 3300 5459 3611 5460
rect 3313 5461 3691 5462
rect 3325 5463 3352 5464
rect 3331 5465 3448 5466
rect 3337 5467 3427 5468
rect 3339 5469 3350 5470
rect 3355 5469 3490 5470
rect 3361 5471 3460 5472
rect 3363 5473 3623 5474
rect 3367 5475 3484 5476
rect 3391 5477 3502 5478
rect 3297 5479 3503 5480
rect 3409 5481 3520 5482
rect 3424 5483 3433 5484
rect 3433 5485 3508 5486
rect 3435 5487 3656 5488
rect 3450 5489 3744 5490
rect 3451 5491 3532 5492
rect 3453 5493 3554 5494
rect 3463 5495 3550 5496
rect 3441 5497 3551 5498
rect 3465 5499 3635 5500
rect 3471 5501 3733 5502
rect 3475 5503 3556 5504
rect 3420 5505 3557 5506
rect 3421 5507 3719 5508
rect 3480 5509 3800 5510
rect 3481 5511 3875 5512
rect 3487 5513 3586 5514
rect 3490 5515 3562 5516
rect 3495 5517 3793 5518
rect 3387 5519 3497 5520
rect 3372 5521 3389 5522
rect 3373 5523 3716 5524
rect 3508 5525 3526 5526
rect 3532 5525 3751 5526
rect 3343 5527 3751 5528
rect 3535 5529 3595 5530
rect 3541 5531 3853 5532
rect 3562 5533 3790 5534
rect 3567 5535 3872 5536
rect 3198 5537 3569 5538
rect 3199 5539 3274 5540
rect 3574 5539 3835 5540
rect 3583 5541 3637 5542
rect 3588 5543 3599 5544
rect 3624 5543 3854 5544
rect 3327 5545 3626 5546
rect 3628 5545 3885 5546
rect 3642 5547 3879 5548
rect 3612 5549 3644 5550
rect 3231 5551 3614 5552
rect 3648 5551 3842 5552
rect 3301 5553 3650 5554
rect 3657 5553 3693 5554
rect 3438 5555 3659 5556
rect 3660 5555 3836 5556
rect 3661 5557 3821 5558
rect 3537 5559 3822 5560
rect 3538 5561 3769 5562
rect 3672 5563 3690 5564
rect 3675 5565 3738 5566
rect 3678 5567 3708 5568
rect 3681 5569 3699 5570
rect 3684 5571 3714 5572
rect 3687 5573 3717 5574
rect 3669 5575 3687 5576
rect 3695 5575 3833 5576
rect 3705 5577 3726 5578
rect 3735 5577 3858 5578
rect 3747 5579 3846 5580
rect 3415 5581 3747 5582
rect 3753 5581 3770 5582
rect 3756 5583 3764 5584
rect 3427 5585 3758 5586
rect 3771 5585 3794 5586
rect 3774 5587 3797 5588
rect 3477 5589 3776 5590
rect 3778 5589 3812 5590
rect 3783 5591 3806 5592
rect 3702 5593 3785 5594
rect 3701 5595 3862 5596
rect 3786 5597 3809 5598
rect 3759 5599 3788 5600
rect 3307 5601 3761 5602
rect 3824 5601 3848 5602
rect 3630 5603 3826 5604
rect 3468 5605 3632 5606
rect 3469 5607 3678 5608
rect 3827 5607 3845 5608
rect 3867 5607 3888 5608
rect 3543 5609 3868 5610
rect 3544 5611 3580 5612
rect 3580 5613 3818 5614
rect 3740 5615 3819 5616
rect 2904 5624 3359 5625
rect 2905 5626 3779 5627
rect 2908 5628 3179 5629
rect 2915 5630 3215 5631
rect 2922 5632 3185 5633
rect 2937 5634 2952 5635
rect 2929 5636 2939 5637
rect 2941 5636 3296 5637
rect 2944 5638 3173 5639
rect 2947 5640 3419 5641
rect 2953 5642 3218 5643
rect 2956 5644 3128 5645
rect 2965 5646 3299 5647
rect 2972 5648 2997 5649
rect 2975 5650 3443 5651
rect 2975 5652 3206 5653
rect 2984 5654 3149 5655
rect 2984 5656 2991 5657
rect 2990 5658 3134 5659
rect 3002 5660 3009 5661
rect 3008 5662 3263 5663
rect 3015 5664 3347 5665
rect 3020 5666 3095 5667
rect 3021 5668 3043 5669
rect 3023 5670 3194 5671
rect 3026 5672 3218 5673
rect 3030 5674 3284 5675
rect 3033 5676 3473 5677
rect 3048 5678 3071 5679
rect 3048 5680 3491 5681
rect 3054 5682 3083 5683
rect 3106 5682 3221 5683
rect 3157 5684 3194 5685
rect 3145 5686 3158 5687
rect 3121 5688 3146 5689
rect 3076 5690 3122 5691
rect 3169 5690 3296 5691
rect 3175 5692 3341 5693
rect 3181 5694 3371 5695
rect 3115 5696 3182 5697
rect 3199 5696 3257 5697
rect 3103 5698 3200 5699
rect 3079 5700 3104 5701
rect 3202 5700 3422 5701
rect 3154 5702 3422 5703
rect 3205 5704 3569 5705
rect 3208 5706 3404 5707
rect 3226 5708 3671 5709
rect 3229 5710 3431 5711
rect 3151 5712 3230 5713
rect 3235 5712 3407 5713
rect 3235 5714 3386 5715
rect 3250 5716 3500 5717
rect 3268 5718 3317 5719
rect 2888 5720 3269 5721
rect 3271 5720 3521 5721
rect 3283 5722 3308 5723
rect 3259 5724 3308 5725
rect 3286 5726 3524 5727
rect 3289 5728 3335 5729
rect 3289 5730 3503 5731
rect 3325 5732 3365 5733
rect 3241 5734 3326 5735
rect 2891 5736 3242 5737
rect 3343 5736 3587 5737
rect 2915 5738 3344 5739
rect 3349 5738 3353 5739
rect 3310 5740 3350 5741
rect 3361 5740 3891 5741
rect 3367 5742 3605 5743
rect 3367 5744 3389 5745
rect 3376 5746 3470 5747
rect 3385 5748 3614 5749
rect 3388 5750 3626 5751
rect 3394 5752 3575 5753
rect 3412 5754 3958 5755
rect 3415 5756 3449 5757
rect 3424 5758 3675 5759
rect 3424 5760 3791 5761
rect 3427 5762 3575 5763
rect 3433 5764 3617 5765
rect 3244 5766 3434 5767
rect 3163 5768 3245 5769
rect 3163 5770 3188 5771
rect 3187 5772 3398 5773
rect 3436 5772 3497 5773
rect 3247 5774 3497 5775
rect 3451 5776 3641 5777
rect 3451 5778 3659 5779
rect 3454 5780 3826 5781
rect 3460 5782 3650 5783
rect 3463 5784 3665 5785
rect 3400 5786 3464 5787
rect 2925 5788 3401 5789
rect 3466 5788 3515 5789
rect 3277 5790 3515 5791
rect 3253 5792 3278 5793
rect 3475 5792 3659 5793
rect 3160 5794 3476 5795
rect 3478 5794 3912 5795
rect 3484 5796 3909 5797
rect 3502 5798 3557 5799
rect 3313 5800 3557 5801
rect 3265 5802 3314 5803
rect 3526 5802 3894 5803
rect 3529 5804 3581 5805
rect 3508 5806 3581 5807
rect 3337 5808 3509 5809
rect 3535 5808 4014 5809
rect 3538 5810 3865 5811
rect 3301 5812 3539 5813
rect 3301 5814 3851 5815
rect 3541 5816 3671 5817
rect 3547 5818 3611 5819
rect 3373 5820 3611 5821
rect 3036 5822 3374 5823
rect 3550 5822 3590 5823
rect 3562 5824 3569 5825
rect 3598 5824 3731 5825
rect 3355 5826 3599 5827
rect 3628 5826 4031 5827
rect 3628 5828 3696 5829
rect 3634 5830 3746 5831
rect 3409 5832 3635 5833
rect 3643 5832 3749 5833
rect 3655 5834 3744 5835
rect 3631 5836 3743 5837
rect 3661 5838 3767 5839
rect 3673 5840 3961 5841
rect 3679 5842 3875 5843
rect 3689 5844 3800 5845
rect 3692 5846 3824 5847
rect 3691 5848 3872 5849
rect 3139 5850 3872 5851
rect 3698 5852 3821 5853
rect 3487 5854 3698 5855
rect 3713 5854 3863 5855
rect 3712 5856 4011 5857
rect 3716 5858 3812 5859
rect 3532 5860 3716 5861
rect 3331 5862 3533 5863
rect 3211 5864 3332 5865
rect 3718 5864 4018 5865
rect 3725 5866 4004 5867
rect 3724 5868 3815 5869
rect 3737 5870 3866 5871
rect 3736 5872 3936 5873
rect 3740 5874 3869 5875
rect 3754 5876 3829 5877
rect 3701 5878 3830 5879
rect 3757 5880 3885 5881
rect 3760 5882 3809 5883
rect 3583 5884 3761 5885
rect 3763 5884 3861 5885
rect 3223 5886 3860 5887
rect 3223 5888 3320 5889
rect 3769 5888 3915 5889
rect 3772 5890 3997 5891
rect 3781 5892 3927 5893
rect 3622 5894 3782 5895
rect 3391 5896 3623 5897
rect 3784 5896 3930 5897
rect 3784 5898 3888 5899
rect 3787 5900 3948 5901
rect 3793 5902 3939 5903
rect 3707 5904 3794 5905
rect 3796 5904 3942 5905
rect 3805 5906 3945 5907
rect 3686 5908 3806 5909
rect 3481 5910 3686 5911
rect 3817 5910 4021 5911
rect 3826 5912 3933 5913
rect 3832 5914 3842 5915
rect 3844 5914 3984 5915
rect 3847 5916 3987 5917
rect 3853 5918 3903 5919
rect 3905 5918 3990 5919
rect 2857 5927 3151 5928
rect 2872 5929 2880 5930
rect 2887 5929 3054 5930
rect 2890 5931 3278 5932
rect 2899 5933 3242 5934
rect 2915 5935 3118 5936
rect 2919 5937 3296 5938
rect 2922 5939 2927 5940
rect 2930 5939 2991 5940
rect 2951 5941 3208 5942
rect 2954 5943 3332 5944
rect 2964 5945 2985 5946
rect 2968 5947 3280 5948
rect 2967 5949 2991 5950
rect 2978 5951 3500 5952
rect 2993 5953 3314 5954
rect 2996 5955 3128 5956
rect 3008 5957 3257 5958
rect 3002 5959 3009 5960
rect 3015 5959 3335 5960
rect 3018 5961 3265 5962
rect 3026 5963 3095 5964
rect 3029 5965 3071 5966
rect 3021 5967 3072 5968
rect 3033 5969 3164 5970
rect 3036 5971 3127 5972
rect 3041 5973 3083 5974
rect 3055 5975 3224 5976
rect 3068 5977 3274 5978
rect 3076 5979 3203 5980
rect 3079 5981 3386 5982
rect 2952 5983 3081 5984
rect 3083 5983 3140 5984
rect 3086 5985 3134 5986
rect 2916 5987 3133 5988
rect 3093 5989 3350 5990
rect 3096 5991 3146 5992
rect 3099 5993 3149 5994
rect 3103 5995 3541 5996
rect 2961 5997 3103 5998
rect 3108 5997 3299 5998
rect 3114 5999 3182 6000
rect 3138 6001 3344 6002
rect 3144 6003 3434 6004
rect 3157 6005 3788 6006
rect 3159 6007 3269 6008
rect 3162 6009 3230 6010
rect 3168 6011 3218 6012
rect 3174 6013 3194 6014
rect 3180 6015 3245 6016
rect 3187 6017 3936 6018
rect 2945 6019 3187 6020
rect 3192 6019 3464 6020
rect 3205 6021 3643 6022
rect 3204 6023 3341 6024
rect 3045 6025 3340 6026
rect 3210 6027 3263 6028
rect 3216 6029 3371 6030
rect 3219 6031 3374 6032
rect 3222 6033 3284 6034
rect 3121 6035 3283 6036
rect 2999 6037 3121 6038
rect 3228 6037 3359 6038
rect 3235 6039 3349 6040
rect 3234 6041 3326 6042
rect 3240 6043 3308 6044
rect 3017 6045 3307 6046
rect 3246 6047 3401 6048
rect 3249 6049 3404 6050
rect 3252 6051 3407 6052
rect 3258 6053 3419 6054
rect 3261 6055 3422 6056
rect 3270 6057 3347 6058
rect 3090 6059 3346 6060
rect 3276 6061 3431 6062
rect 3289 6063 3481 6064
rect 3294 6065 3473 6066
rect 3297 6067 3476 6068
rect 3309 6069 3317 6070
rect 3312 6071 3497 6072
rect 3315 6073 3443 6074
rect 3318 6075 3365 6076
rect 3330 6077 3515 6078
rect 3336 6079 3521 6080
rect 3342 6081 3461 6082
rect 3354 6083 3703 6084
rect 3360 6085 3545 6086
rect 3372 6087 3557 6088
rect 3384 6089 3509 6090
rect 3388 6091 3700 6092
rect 3390 6093 3527 6094
rect 3376 6095 3526 6096
rect 3402 6097 3631 6098
rect 3408 6099 3611 6100
rect 3412 6101 3607 6102
rect 3414 6103 3599 6104
rect 3420 6105 3605 6106
rect 3432 6107 3485 6108
rect 3438 6109 3623 6110
rect 3444 6111 3933 6112
rect 3448 6113 3637 6114
rect 3456 6115 3635 6116
rect 3451 6117 3634 6118
rect 3450 6119 3617 6120
rect 3462 6121 3575 6122
rect 3474 6123 3961 6124
rect 3478 6125 3958 6126
rect 3486 6127 3659 6128
rect 3454 6129 3658 6130
rect 3492 6131 3671 6132
rect 3495 6133 3665 6134
rect 3513 6135 3686 6136
rect 3519 6137 3692 6138
rect 3523 6139 3706 6140
rect 3529 6141 3604 6142
rect 3538 6143 3761 6144
rect 3199 6145 3538 6146
rect 3543 6145 3653 6146
rect 3549 6147 3581 6148
rect 3466 6149 3580 6150
rect 3553 6151 3577 6152
rect 3555 6153 3713 6154
rect 3532 6155 3713 6156
rect 3301 6157 3532 6158
rect 3558 6157 3680 6158
rect 3561 6159 3674 6160
rect 3367 6161 3673 6162
rect 3366 6163 3425 6164
rect 3568 6163 3592 6164
rect 3394 6165 3568 6166
rect 3573 6165 3590 6166
rect 3615 6165 3725 6166
rect 3621 6167 3731 6168
rect 3628 6169 3875 6170
rect 3396 6171 3628 6172
rect 3640 6171 3894 6172
rect 3547 6173 3640 6174
rect 3651 6173 3749 6174
rect 3663 6175 4000 6176
rect 3687 6177 3755 6178
rect 3693 6179 3743 6180
rect 3697 6181 4038 6182
rect 3696 6183 3779 6184
rect 3715 6185 4014 6186
rect 3718 6187 4028 6188
rect 3727 6189 3806 6190
rect 3730 6191 3800 6192
rect 3733 6193 3818 6194
rect 3736 6195 3951 6196
rect 3736 6197 3824 6198
rect 3739 6199 3827 6200
rect 3745 6201 3891 6202
rect 3748 6203 3824 6204
rect 3760 6205 3860 6206
rect 3763 6207 3863 6208
rect 3766 6209 3997 6210
rect 3766 6211 3869 6212
rect 3769 6213 3794 6214
rect 3586 6215 3794 6216
rect 3502 6217 3586 6218
rect 3048 6219 3502 6220
rect 3772 6219 3815 6220
rect 3436 6221 3773 6222
rect 3779 6221 3791 6222
rect 3784 6223 4041 6224
rect 3786 6225 3866 6226
rect 3796 6227 3845 6228
rect 3805 6229 3939 6230
rect 3808 6231 3942 6232
rect 3811 6233 3927 6234
rect 3817 6235 3945 6236
rect 3826 6237 3842 6238
rect 3781 6239 3841 6240
rect 3829 6241 3854 6242
rect 3789 6243 3831 6244
rect 3847 6243 3906 6244
rect 3850 6245 3987 6246
rect 3859 6247 3885 6248
rect 3820 6249 3885 6250
rect 3820 6251 3948 6252
rect 3866 6253 3915 6254
rect 3902 6255 3993 6256
rect 3929 6257 4004 6258
rect 3953 6259 3984 6260
rect 2872 6268 3151 6269
rect 2875 6270 3065 6271
rect 2879 6272 2914 6273
rect 2878 6274 3054 6275
rect 2897 6276 3160 6277
rect 2902 6278 3097 6279
rect 2903 6280 3081 6281
rect 2906 6282 3220 6283
rect 2909 6284 3700 6285
rect 2910 6286 3191 6287
rect 2914 6288 3247 6289
rect 2927 6290 3133 6291
rect 2930 6292 3139 6293
rect 2933 6294 2940 6295
rect 2945 6294 3221 6295
rect 2948 6296 3163 6297
rect 2948 6298 3155 6299
rect 2964 6300 3259 6301
rect 2967 6302 3100 6303
rect 2967 6304 3239 6305
rect 2971 6306 3015 6307
rect 2971 6308 3257 6309
rect 2978 6310 3107 6311
rect 2955 6312 2979 6313
rect 2955 6314 2982 6315
rect 2999 6314 3103 6315
rect 3016 6316 3305 6317
rect 3026 6318 3032 6319
rect 3029 6320 3059 6321
rect 3046 6322 3118 6323
rect 3061 6324 3250 6325
rect 3086 6326 3137 6327
rect 3067 6328 3086 6329
rect 3090 6328 3319 6329
rect 2952 6330 3092 6331
rect 2907 6332 2953 6333
rect 3093 6332 3352 6333
rect 3100 6334 3193 6335
rect 3103 6336 3346 6337
rect 3108 6338 3113 6339
rect 3114 6338 3119 6339
rect 3126 6338 3343 6339
rect 3070 6340 3344 6341
rect 3129 6342 3397 6343
rect 3120 6344 3131 6345
rect 2923 6346 3122 6347
rect 3142 6346 3145 6347
rect 3148 6346 3169 6347
rect 3166 6348 3181 6349
rect 3172 6350 3175 6351
rect 3178 6350 3283 6351
rect 3184 6352 3187 6353
rect 3196 6352 3205 6353
rect 3199 6354 3208 6355
rect 3202 6356 3211 6357
rect 3041 6358 3212 6359
rect 3208 6360 3217 6361
rect 3214 6362 3229 6363
rect 3222 6364 3233 6365
rect 3226 6366 3538 6367
rect 3234 6368 3245 6369
rect 3250 6368 3253 6369
rect 3264 6368 3287 6369
rect 3268 6370 3316 6371
rect 3270 6372 3317 6373
rect 3273 6374 3320 6375
rect 3274 6376 3277 6377
rect 3277 6378 3280 6379
rect 3292 6378 3295 6379
rect 3295 6380 3298 6381
rect 3298 6382 3307 6383
rect 3307 6384 3310 6385
rect 3310 6386 3313 6387
rect 2981 6388 3314 6389
rect 3328 6388 3331 6389
rect 3334 6388 3337 6389
rect 3337 6390 3340 6391
rect 3340 6392 3349 6393
rect 3346 6394 3403 6395
rect 3349 6396 3541 6397
rect 3352 6398 3675 6399
rect 3354 6400 3395 6401
rect 3358 6402 3361 6403
rect 3364 6402 3481 6403
rect 3366 6404 3389 6405
rect 3367 6406 3643 6407
rect 3370 6408 3373 6409
rect 3376 6408 3385 6409
rect 3382 6410 3391 6411
rect 3400 6410 3713 6411
rect 3406 6412 3753 6413
rect 3408 6414 3779 6415
rect 3412 6416 3415 6417
rect 3418 6416 3421 6417
rect 3424 6416 3773 6417
rect 3430 6418 3433 6419
rect 3436 6418 3463 6419
rect 3442 6420 3457 6421
rect 3444 6422 3449 6423
rect 3454 6422 3526 6423
rect 3466 6424 3783 6425
rect 3472 6426 3496 6427
rect 3474 6428 3831 6429
rect 3478 6430 3493 6431
rect 3493 6432 3514 6433
rect 3501 6434 3628 6435
rect 3505 6436 3580 6437
rect 3511 6438 3592 6439
rect 3517 6440 3544 6441
rect 3519 6442 3527 6443
rect 3523 6444 3556 6445
rect 3529 6446 3586 6447
rect 3531 6448 3584 6449
rect 3535 6450 3550 6451
rect 3553 6450 3803 6451
rect 3556 6452 3577 6453
rect 3558 6454 3881 6455
rect 3561 6456 3846 6457
rect 3565 6458 3616 6459
rect 3567 6460 3572 6461
rect 3589 6460 3604 6461
rect 3592 6462 3609 6463
rect 3595 6464 3634 6465
rect 3598 6466 3640 6467
rect 3606 6468 3703 6469
rect 3611 6470 3658 6471
rect 3617 6472 3841 6473
rect 3630 6474 3794 6475
rect 3621 6476 3794 6477
rect 3636 6478 3756 6479
rect 3635 6480 3652 6481
rect 3641 6482 3664 6483
rect 3647 6484 3688 6485
rect 3653 6486 3815 6487
rect 3659 6488 3697 6489
rect 3662 6490 3666 6491
rect 3669 6490 3706 6491
rect 3000 6492 3669 6493
rect 3672 6492 3776 6493
rect 3677 6494 3694 6495
rect 3698 6494 3728 6495
rect 3701 6496 3824 6497
rect 3704 6498 3737 6499
rect 3707 6500 3740 6501
rect 3716 6502 3761 6503
rect 3541 6504 3760 6505
rect 3719 6506 3749 6507
rect 3728 6508 3770 6509
rect 3573 6510 3770 6511
rect 3733 6512 3888 6513
rect 3734 6514 3767 6515
rect 3746 6516 3790 6517
rect 3749 6518 3787 6519
rect 3763 6520 3827 6521
rect 3559 6522 3763 6523
rect 3730 6524 3827 6525
rect 3772 6526 3812 6527
rect 3790 6528 3806 6529
rect 3450 6530 3806 6531
rect 3796 6532 3838 6533
rect 3796 6534 3818 6535
rect 3799 6536 3821 6537
rect 3671 6538 3820 6539
rect 3808 6540 3843 6541
rect 3438 6542 3810 6543
rect 3829 6542 3851 6543
rect 3832 6544 3854 6545
rect 3847 6546 3867 6547
rect 3859 6548 3871 6549
rect 3008 6550 3870 6551
rect 3863 6552 3874 6553
rect 2887 6561 2897 6562
rect 2890 6563 3065 6564
rect 2900 6565 3269 6566
rect 2903 6567 3145 6568
rect 2907 6569 2922 6570
rect 2907 6571 3155 6572
rect 2924 6573 3203 6574
rect 2924 6575 3047 6576
rect 2928 6577 3046 6578
rect 2933 6579 2941 6580
rect 2945 6579 3215 6580
rect 2952 6581 3082 6582
rect 2962 6583 2992 6584
rect 2964 6585 3259 6586
rect 2974 6587 3251 6588
rect 2974 6589 3247 6590
rect 2981 6591 3242 6592
rect 2985 6593 3191 6594
rect 2995 6595 3293 6596
rect 3004 6597 3032 6598
rect 3006 6599 3107 6600
rect 2917 6601 3106 6602
rect 3000 6603 3008 6604
rect 3013 6603 3606 6604
rect 3016 6605 3253 6606
rect 3030 6607 3335 6608
rect 3034 6609 3338 6610
rect 3033 6611 3059 6612
rect 3037 6613 3322 6614
rect 3036 6615 3062 6616
rect 3063 6615 3331 6616
rect 3070 6617 3334 6618
rect 3085 6619 3350 6620
rect 3084 6621 3092 6622
rect 3100 6621 3190 6622
rect 3099 6623 3113 6624
rect 3108 6625 3119 6626
rect 3111 6627 3122 6628
rect 3126 6627 3131 6628
rect 3132 6627 3143 6628
rect 3136 6629 3235 6630
rect 3138 6631 3149 6632
rect 3150 6631 3167 6632
rect 3156 6633 3344 6634
rect 3162 6635 3173 6636
rect 3165 6637 3296 6638
rect 3020 6639 3295 6640
rect 3174 6641 3185 6642
rect 3178 6643 3439 6644
rect 3180 6645 3197 6646
rect 3183 6647 3200 6648
rect 3192 6649 3209 6650
rect 3195 6651 3212 6652
rect 3204 6653 3221 6654
rect 3210 6655 3233 6656
rect 3216 6657 3245 6658
rect 3222 6659 3239 6660
rect 3226 6661 3356 6662
rect 2952 6663 3226 6664
rect 3228 6663 3263 6664
rect 3240 6665 3257 6666
rect 3264 6665 3275 6666
rect 3267 6667 3278 6668
rect 3270 6669 3287 6670
rect 3276 6671 3317 6672
rect 3282 6673 3299 6674
rect 3288 6675 3305 6676
rect 3291 6677 3308 6678
rect 3300 6679 3311 6680
rect 3303 6681 3314 6682
rect 3088 6683 3313 6684
rect 2971 6685 3088 6686
rect 2971 6687 3262 6688
rect 3315 6687 3320 6688
rect 3318 6689 3329 6690
rect 3324 6691 3341 6692
rect 3339 6693 3353 6694
rect 3348 6695 3359 6696
rect 3364 6695 3391 6696
rect 3367 6697 3598 6698
rect 3366 6699 3371 6700
rect 3372 6699 3864 6700
rect 3376 6701 3379 6702
rect 3382 6701 3385 6702
rect 3388 6701 3397 6702
rect 3394 6703 3421 6704
rect 3402 6705 3413 6706
rect 3406 6707 3427 6708
rect 3418 6709 3586 6710
rect 3430 6711 3457 6712
rect 3432 6713 3745 6714
rect 3436 6715 3451 6716
rect 3448 6717 3463 6718
rect 3468 6717 3808 6718
rect 3472 6719 3490 6720
rect 3478 6721 3481 6722
rect 3487 6721 3502 6722
rect 3493 6723 3508 6724
rect 3511 6723 3811 6724
rect 3523 6725 3817 6726
rect 3517 6727 3523 6728
rect 3526 6727 3853 6728
rect 3535 6729 3547 6730
rect 3529 6731 3535 6732
rect 3505 6733 3529 6734
rect 3571 6733 3760 6734
rect 3565 6735 3571 6736
rect 3559 6737 3565 6738
rect 3576 6737 3584 6738
rect 3582 6739 3794 6740
rect 3589 6741 3609 6742
rect 3342 6743 3610 6744
rect 3588 6745 3593 6746
rect 3400 6747 3592 6748
rect 3603 6747 3618 6748
rect 3611 6749 3622 6750
rect 3360 6751 3613 6752
rect 3627 6751 3660 6752
rect 3630 6753 3669 6754
rect 3466 6755 3670 6756
rect 3633 6757 3642 6758
rect 3635 6759 3640 6760
rect 3645 6759 3654 6760
rect 3474 6761 3655 6762
rect 3651 6763 3769 6764
rect 3662 6765 3841 6766
rect 3663 6767 3672 6768
rect 3424 6769 3673 6770
rect 3666 6771 3675 6772
rect 3454 6773 3676 6774
rect 3677 6773 3778 6774
rect 3678 6775 3776 6776
rect 3690 6777 3717 6778
rect 3693 6779 3720 6780
rect 3696 6781 3702 6782
rect 3698 6783 3827 6784
rect 3442 6785 3700 6786
rect 3346 6787 3442 6788
rect 3103 6789 3346 6790
rect 3702 6789 3705 6790
rect 3705 6791 3708 6792
rect 3714 6791 3785 6792
rect 3720 6793 3729 6794
rect 3726 6795 3735 6796
rect 3732 6797 3750 6798
rect 3746 6799 3754 6800
rect 3750 6801 3806 6802
rect 3756 6803 3773 6804
rect 3771 6805 3820 6806
rect 3794 6807 3797 6808
rect 3647 6809 3798 6810
rect 3799 6809 3846 6810
rect 3827 6811 3830 6812
rect 3830 6813 3836 6814
rect 3832 6815 3839 6816
rect 3849 6815 3865 6816
rect 3790 6817 3851 6818
rect 3408 6819 3792 6820
rect 2896 6828 3106 6829
rect 2907 6830 3145 6831
rect 2912 6832 3181 6833
rect 2914 6834 3243 6835
rect 2922 6836 3265 6837
rect 2924 6838 3046 6839
rect 2940 6840 2972 6841
rect 2952 6842 3114 6843
rect 2959 6844 2967 6845
rect 2963 6846 3184 6847
rect 2978 6848 3259 6849
rect 2979 6850 3139 6851
rect 2981 6852 3028 6853
rect 2982 6854 3005 6855
rect 2917 6856 3005 6857
rect 2985 6858 3253 6859
rect 2988 6860 3014 6861
rect 2995 6862 3285 6863
rect 3007 6864 3011 6865
rect 3022 6864 3034 6865
rect 3034 6866 3316 6867
rect 3036 6868 3252 6869
rect 3037 6870 3255 6871
rect 3044 6872 3279 6873
rect 3059 6874 3082 6875
rect 3066 6876 3292 6877
rect 3065 6878 3088 6879
rect 3071 6880 3291 6881
rect 3077 6882 3100 6883
rect 3086 6884 3112 6885
rect 3092 6886 3325 6887
rect 3101 6888 3133 6889
rect 3119 6890 3151 6891
rect 3143 6892 3175 6893
rect 3149 6894 3157 6895
rect 3167 6894 3211 6895
rect 3173 6896 3217 6897
rect 3179 6898 3193 6899
rect 2928 6900 3192 6901
rect 2929 6902 3249 6903
rect 3182 6904 3196 6905
rect 3084 6906 3195 6907
rect 3083 6908 3109 6909
rect 3107 6910 3127 6911
rect 3125 6912 3163 6913
rect 3161 6914 3205 6915
rect 2903 6916 3204 6917
rect 3189 6918 3346 6919
rect 3206 6920 3271 6921
rect 3212 6922 3223 6923
rect 3215 6924 3226 6925
rect 2974 6926 3225 6927
rect 3218 6928 3277 6929
rect 3230 6930 3241 6931
rect 3234 6932 3315 6933
rect 3233 6934 3268 6935
rect 3236 6936 3247 6937
rect 3266 6936 3283 6937
rect 3272 6938 3289 6939
rect 3165 6940 3288 6941
rect 3300 6940 3309 6941
rect 3228 6942 3300 6943
rect 3227 6944 3262 6945
rect 3318 6944 3327 6945
rect 3323 6946 3676 6947
rect 3330 6948 3339 6949
rect 3321 6950 3330 6951
rect 3312 6952 3321 6953
rect 3303 6954 3312 6955
rect 3294 6956 3303 6957
rect 3342 6956 3345 6957
rect 3333 6958 3342 6959
rect 3296 6960 3333 6961
rect 3348 6960 3354 6961
rect 3063 6962 3348 6963
rect 3402 6962 3835 6963
rect 3372 6964 3402 6965
rect 3366 6966 3372 6967
rect 3360 6968 3366 6969
rect 3408 6968 3414 6969
rect 3426 6968 3789 6969
rect 3390 6970 3426 6971
rect 3378 6972 3390 6973
rect 3336 6974 3378 6975
rect 3335 6976 3475 6977
rect 3441 6978 3465 6979
rect 3456 6980 3811 6981
rect 3450 6982 3456 6983
rect 3473 6982 3863 6983
rect 3480 6984 3486 6985
rect 3468 6986 3480 6987
rect 3462 6988 3468 6989
rect 3438 6990 3462 6991
rect 3432 6992 3438 6993
rect 3396 6994 3432 6995
rect 3384 6996 3396 6997
rect 3383 6998 3615 6999
rect 3489 7000 3841 7001
rect 3494 7002 3673 7003
rect 3501 7004 3513 7005
rect 3522 7004 3531 7005
rect 3524 7006 3670 7007
rect 3528 7008 3543 7009
rect 3534 7010 3549 7011
rect 3536 7012 3577 7013
rect 3546 7014 3561 7015
rect 3552 7016 3567 7017
rect 3564 7018 3576 7019
rect 3572 7020 3706 7021
rect 3591 7022 3655 7023
rect 3420 7024 3591 7025
rect 3419 7026 3586 7027
rect 3600 7026 3729 7027
rect 3594 7028 3600 7029
rect 3603 7028 3624 7029
rect 3597 7030 3603 7031
rect 3627 7030 3654 7031
rect 3630 7032 3657 7033
rect 3633 7034 3874 7035
rect 3639 7036 3648 7037
rect 3666 7036 3684 7037
rect 3645 7038 3666 7039
rect 3686 7038 3778 7039
rect 3507 7040 3779 7041
rect 3506 7042 3818 7043
rect 3693 7044 3717 7045
rect 2951 7046 3693 7047
rect 3696 7046 3708 7047
rect 3678 7048 3696 7049
rect 3699 7048 3711 7049
rect 3702 7050 3844 7051
rect 3720 7052 3782 7053
rect 3719 7054 3831 7055
rect 3407 7056 3832 7057
rect 3722 7058 3837 7059
rect 3726 7060 3785 7061
rect 3609 7062 3726 7063
rect 3747 7062 3825 7063
rect 3756 7064 3782 7065
rect 3617 7066 3756 7067
rect 3765 7066 3808 7067
rect 3753 7068 3809 7069
rect 3732 7070 3753 7071
rect 3714 7072 3732 7073
rect 3690 7074 3714 7075
rect 3663 7076 3690 7077
rect 3775 7076 3867 7077
rect 3794 7078 3800 7079
rect 3768 7080 3794 7081
rect 3797 7080 3803 7081
rect 3771 7082 3797 7083
rect 3621 7084 3773 7085
rect 3811 7084 3851 7085
rect 3814 7086 3828 7087
rect 3582 7088 3815 7089
rect 3570 7090 3582 7091
rect 3555 7092 3570 7093
rect 3540 7094 3555 7095
rect 3854 7094 3865 7095
rect 2893 7103 3204 7104
rect 2908 7105 3205 7106
rect 2911 7107 2964 7108
rect 2915 7109 3102 7110
rect 2919 7111 3195 7112
rect 2918 7113 3084 7114
rect 2921 7115 3078 7116
rect 2926 7117 3252 7118
rect 2925 7119 3249 7120
rect 2928 7121 3106 7122
rect 2950 7123 3190 7124
rect 2954 7125 3192 7126
rect 2956 7127 2967 7128
rect 2959 7129 3082 7130
rect 2969 7131 3097 7132
rect 2969 7133 3462 7134
rect 2972 7135 3228 7136
rect 2973 7137 3237 7138
rect 2966 7139 3238 7140
rect 2976 7141 3114 7142
rect 2985 7143 3307 7144
rect 2995 7145 3094 7146
rect 2994 7147 3011 7148
rect 3000 7149 3005 7150
rect 3006 7149 3064 7150
rect 3009 7151 3255 7152
rect 3022 7153 3259 7154
rect 3030 7155 3066 7156
rect 3037 7157 3273 7158
rect 2979 7159 3037 7160
rect 2979 7161 2983 7162
rect 3041 7161 3162 7162
rect 3042 7163 3321 7164
rect 3048 7165 3060 7166
rect 3060 7167 3166 7168
rect 3074 7169 3339 7170
rect 3075 7171 3312 7172
rect 3086 7173 3241 7174
rect 3087 7175 3315 7176
rect 3107 7177 3678 7178
rect 3111 7179 3120 7180
rect 3117 7181 3126 7182
rect 3123 7183 3150 7184
rect 3129 7185 3279 7186
rect 3143 7187 3154 7188
rect 3147 7189 3216 7190
rect 3167 7191 3178 7192
rect 3171 7193 3180 7194
rect 3173 7195 3196 7196
rect 3174 7197 3183 7198
rect 3197 7197 3262 7198
rect 3200 7199 3426 7200
rect 3201 7201 3213 7202
rect 3206 7203 3214 7204
rect 3057 7205 3208 7206
rect 3222 7205 3234 7206
rect 3224 7207 3744 7208
rect 3218 7209 3226 7210
rect 3219 7211 3231 7212
rect 3231 7213 3330 7214
rect 3071 7215 3331 7216
rect 3242 7217 3256 7218
rect 3089 7219 3244 7220
rect 3246 7219 3342 7220
rect 3144 7221 3343 7222
rect 3287 7223 3295 7224
rect 3288 7225 3345 7226
rect 3299 7227 3313 7228
rect 3302 7229 3316 7230
rect 3303 7231 3309 7232
rect 3296 7233 3310 7234
rect 3290 7235 3298 7236
rect 3284 7237 3292 7238
rect 3132 7239 3286 7240
rect 3318 7239 3324 7240
rect 3321 7241 3336 7242
rect 3333 7243 3603 7244
rect 3339 7245 3348 7246
rect 3345 7247 3384 7248
rect 3348 7249 3600 7250
rect 3351 7251 3390 7252
rect 3353 7253 3737 7254
rect 3357 7255 3378 7256
rect 3363 7257 3366 7258
rect 3369 7257 3372 7258
rect 3381 7257 3591 7258
rect 3393 7259 3495 7260
rect 3399 7261 3414 7262
rect 3401 7263 3612 7264
rect 3405 7265 3408 7266
rect 3411 7265 3763 7266
rect 3423 7267 3537 7268
rect 3429 7269 3456 7270
rect 3431 7271 3747 7272
rect 3435 7273 3818 7274
rect 3437 7275 3766 7276
rect 3441 7277 3711 7278
rect 3450 7279 3468 7280
rect 3456 7281 3570 7282
rect 3462 7283 3773 7284
rect 3464 7285 3704 7286
rect 3395 7287 3466 7288
rect 3468 7287 3543 7288
rect 3473 7289 3867 7290
rect 3474 7291 3486 7292
rect 3477 7293 3513 7294
rect 3479 7295 3863 7296
rect 3483 7297 3779 7298
rect 3489 7299 3576 7300
rect 3501 7301 3531 7302
rect 3513 7303 3729 7304
rect 3506 7305 3730 7306
rect 3507 7307 3561 7308
rect 3519 7309 3573 7310
rect 3522 7311 3582 7312
rect 3528 7313 3618 7314
rect 3534 7315 3806 7316
rect 3537 7317 3567 7318
rect 3546 7319 3687 7320
rect 3552 7321 3654 7322
rect 3554 7323 3652 7324
rect 3555 7325 3657 7326
rect 3564 7327 3723 7328
rect 3582 7329 3659 7330
rect 3587 7331 3759 7332
rect 3600 7333 3714 7334
rect 3603 7335 3717 7336
rect 3606 7337 3690 7338
rect 3609 7339 3693 7340
rect 3618 7341 3696 7342
rect 3623 7343 3860 7344
rect 3624 7345 3720 7346
rect 3419 7347 3720 7348
rect 3627 7349 3853 7350
rect 3636 7351 3750 7352
rect 3639 7353 3732 7354
rect 3642 7355 3656 7356
rect 3645 7357 3726 7358
rect 3661 7359 3800 7360
rect 3665 7361 3765 7362
rect 3647 7363 3665 7364
rect 3387 7365 3649 7366
rect 3667 7365 3684 7366
rect 3680 7367 3803 7368
rect 3679 7369 3776 7370
rect 3682 7371 3772 7372
rect 3685 7373 3782 7374
rect 3697 7375 3794 7376
rect 3700 7377 3797 7378
rect 3707 7379 3842 7380
rect 3548 7381 3707 7382
rect 3524 7383 3550 7384
rect 3716 7383 3812 7384
rect 3752 7385 3756 7386
rect 3757 7385 3839 7386
rect 3814 7387 3821 7388
rect 2911 7396 2957 7397
rect 2918 7398 3001 7399
rect 2928 7400 3256 7401
rect 2935 7402 3190 7403
rect 2962 7404 3346 7405
rect 2962 7406 3334 7407
rect 2966 7408 3292 7409
rect 2969 7410 3316 7411
rect 2969 7412 3037 7413
rect 2925 7414 3036 7415
rect 2973 7416 3005 7417
rect 2979 7418 2990 7419
rect 2985 7420 3295 7421
rect 2979 7422 2987 7423
rect 2994 7422 3136 7423
rect 3006 7424 3253 7425
rect 3007 7426 3051 7427
rect 3009 7428 3232 7429
rect 3017 7430 3046 7431
rect 3038 7432 3259 7433
rect 3042 7434 3412 7435
rect 3030 7436 3042 7437
rect 3054 7436 3091 7437
rect 2953 7438 3091 7439
rect 3057 7440 3331 7441
rect 3057 7442 3169 7443
rect 3063 7444 3079 7445
rect 3075 7446 3103 7447
rect 3093 7448 3109 7449
rect 3105 7450 3121 7451
rect 3111 7452 3127 7453
rect 3096 7454 3112 7455
rect 3081 7456 3097 7457
rect 3114 7456 3418 7457
rect 3123 7458 3139 7459
rect 3129 7460 3244 7461
rect 3132 7462 3400 7463
rect 3117 7464 3133 7465
rect 3147 7464 3151 7465
rect 3153 7464 3157 7465
rect 3165 7464 3316 7465
rect 3171 7466 3187 7467
rect 3171 7468 3247 7469
rect 3174 7470 3190 7471
rect 2958 7472 3175 7473
rect 3177 7472 3211 7473
rect 3048 7474 3178 7475
rect 3047 7476 3301 7477
rect 3192 7478 3196 7479
rect 3207 7478 3259 7479
rect 3213 7480 3229 7481
rect 3219 7482 3247 7483
rect 2914 7484 3220 7485
rect 2914 7486 3217 7487
rect 3222 7486 3250 7487
rect 3201 7488 3223 7489
rect 3234 7488 3238 7489
rect 3237 7490 3241 7491
rect 3225 7492 3241 7493
rect 3204 7494 3226 7495
rect 2932 7496 3205 7497
rect 3243 7496 3319 7497
rect 3261 7498 3277 7499
rect 3267 7500 3271 7501
rect 3144 7502 3268 7503
rect 3282 7502 3298 7503
rect 3285 7504 3346 7505
rect 3291 7506 3307 7507
rect 3294 7508 3310 7509
rect 3297 7510 3313 7511
rect 3306 7512 3322 7513
rect 3312 7514 3328 7515
rect 3318 7516 3331 7517
rect 3342 7516 3361 7517
rect 3288 7518 3343 7519
rect 3288 7520 3304 7521
rect 3348 7520 3385 7521
rect 3348 7522 3364 7523
rect 3339 7524 3364 7525
rect 3351 7526 3373 7527
rect 3354 7528 3358 7529
rect 3369 7528 3737 7529
rect 3387 7530 3415 7531
rect 3381 7532 3388 7533
rect 3390 7532 3406 7533
rect 3393 7534 3409 7535
rect 3396 7536 3559 7537
rect 3399 7538 3466 7539
rect 3402 7540 3720 7541
rect 3420 7542 3550 7543
rect 3426 7544 3442 7545
rect 3435 7546 3442 7547
rect 3429 7548 3436 7549
rect 3423 7550 3430 7551
rect 3447 7550 3457 7551
rect 3453 7552 3469 7553
rect 3459 7554 3475 7555
rect 3462 7556 3562 7557
rect 3462 7558 3711 7559
rect 3468 7560 3529 7561
rect 3477 7562 3481 7563
rect 3483 7562 3487 7563
rect 3489 7562 3649 7563
rect 3510 7564 3705 7565
rect 3513 7566 3623 7567
rect 3525 7568 3535 7569
rect 3528 7570 3538 7571
rect 3537 7572 3630 7573
rect 3540 7574 3547 7575
rect 3543 7576 3553 7577
rect 3546 7578 3556 7579
rect 3561 7578 3665 7579
rect 3573 7580 3583 7581
rect 3579 7582 3601 7583
rect 3582 7584 3604 7585
rect 3564 7586 3604 7587
rect 3507 7588 3565 7589
rect 3507 7590 3520 7591
rect 3585 7590 3610 7591
rect 3594 7592 3619 7593
rect 3576 7594 3620 7595
rect 3600 7596 3625 7597
rect 3606 7598 3782 7599
rect 3606 7600 3640 7601
rect 3450 7602 3641 7603
rect 3609 7604 3730 7605
rect 3612 7606 3662 7607
rect 3627 7608 3726 7609
rect 3633 7610 3637 7611
rect 3642 7610 3659 7611
rect 3645 7612 3656 7613
rect 3643 7614 3656 7615
rect 3652 7616 3717 7617
rect 3658 7618 3686 7619
rect 3670 7620 3723 7621
rect 3522 7622 3722 7623
rect 3670 7624 3698 7625
rect 3673 7626 3701 7627
rect 3679 7628 3775 7629
rect 3321 7630 3680 7631
rect 3682 7630 3728 7631
rect 3743 7630 3761 7631
rect 2809 7639 3448 7640
rect 2888 7641 2895 7642
rect 2924 7641 3061 7642
rect 2928 7643 3039 7644
rect 2931 7645 3220 7646
rect 2964 7647 3274 7648
rect 2967 7649 3247 7650
rect 2969 7651 3042 7652
rect 2972 7653 3018 7654
rect 2986 7655 3322 7656
rect 2989 7657 3014 7658
rect 3035 7657 3064 7658
rect 3039 7659 3406 7660
rect 3050 7661 3277 7662
rect 3057 7663 3145 7664
rect 2960 7665 3145 7666
rect 3072 7667 3079 7668
rect 3078 7669 3115 7670
rect 3084 7671 3103 7672
rect 3102 7673 3109 7674
rect 3105 7675 3112 7676
rect 3108 7677 3139 7678
rect 3114 7679 3133 7680
rect 3117 7681 3136 7682
rect 3120 7683 3139 7684
rect 3123 7685 3352 7686
rect 3129 7687 3172 7688
rect 3156 7689 3181 7690
rect 2957 7691 3157 7692
rect 3165 7691 3364 7692
rect 3174 7693 3199 7694
rect 3177 7695 3202 7696
rect 3189 7697 3214 7698
rect 3204 7699 3319 7700
rect 3216 7701 3265 7702
rect 3192 7703 3217 7704
rect 3219 7703 3250 7704
rect 3222 7705 3247 7706
rect 3210 7707 3223 7708
rect 3186 7709 3211 7710
rect 3225 7709 3250 7710
rect 3234 7711 3286 7712
rect 3234 7713 3241 7714
rect 3029 7715 3241 7716
rect 3252 7715 3268 7716
rect 3252 7717 3259 7718
rect 3270 7717 3310 7718
rect 3282 7719 3334 7720
rect 3288 7721 3358 7722
rect 2921 7723 3289 7724
rect 2920 7725 3017 7726
rect 3294 7725 3340 7726
rect 3300 7727 3304 7728
rect 3312 7727 3364 7728
rect 3327 7729 3346 7730
rect 3306 7731 3346 7732
rect 3330 7733 3382 7734
rect 3348 7735 3424 7736
rect 3369 7737 3469 7738
rect 3372 7739 3394 7740
rect 3375 7741 3388 7742
rect 3032 7743 3388 7744
rect 3390 7743 3466 7744
rect 3315 7745 3391 7746
rect 3399 7745 3418 7746
rect 3354 7747 3400 7748
rect 3342 7749 3355 7750
rect 3297 7751 3343 7752
rect 3297 7753 3430 7754
rect 3402 7755 3472 7756
rect 3411 7757 3415 7758
rect 3384 7759 3415 7760
rect 3420 7759 3722 7760
rect 3396 7761 3421 7762
rect 3426 7761 3496 7762
rect 3426 7763 3547 7764
rect 3429 7765 3463 7766
rect 3435 7767 3666 7768
rect 3435 7769 3454 7770
rect 3441 7771 3478 7772
rect 3162 7773 3442 7774
rect 3447 7773 3651 7774
rect 3459 7775 3523 7776
rect 3459 7777 3641 7778
rect 3453 7779 3640 7780
rect 3486 7781 3634 7782
rect 3504 7783 3713 7784
rect 3510 7785 3701 7786
rect 3150 7787 3511 7788
rect 3126 7789 3151 7790
rect 3126 7791 3169 7792
rect 3516 7791 3708 7792
rect 3525 7793 3553 7794
rect 3480 7795 3526 7796
rect 3528 7795 3556 7796
rect 3537 7797 3568 7798
rect 3507 7799 3538 7800
rect 3540 7799 3620 7800
rect 3501 7801 3541 7802
rect 3543 7801 3598 7802
rect 3561 7803 3589 7804
rect 3564 7805 3592 7806
rect 3564 7807 3630 7808
rect 3570 7809 3574 7810
rect 3573 7811 3577 7812
rect 3579 7811 3696 7812
rect 3582 7813 3663 7814
rect 3585 7815 3728 7816
rect 3594 7817 3619 7818
rect 3237 7819 3595 7820
rect 3237 7821 3244 7822
rect 3600 7821 3625 7822
rect 3600 7823 3610 7824
rect 3603 7825 3628 7826
rect 3606 7827 3616 7828
rect 3612 7829 3637 7830
rect 3630 7831 3731 7832
rect 3655 7833 3703 7834
rect 3656 7835 3734 7836
rect 3670 7837 3690 7838
rect 3652 7839 3672 7840
rect 3673 7839 3693 7840
rect 3674 7841 3687 7842
rect 3676 7843 3706 7844
rect 3658 7845 3678 7846
rect 3659 7847 3680 7848
rect 2884 7856 2895 7857
rect 2888 7858 2918 7859
rect 2914 7860 3064 7861
rect 2918 7862 3286 7863
rect 2921 7864 3199 7865
rect 2931 7866 3007 7867
rect 2946 7868 3289 7869
rect 2960 7870 3139 7871
rect 2961 7872 3109 7873
rect 2965 7874 3268 7875
rect 2967 7876 3235 7877
rect 2968 7878 3130 7879
rect 2975 7880 3137 7881
rect 2995 7882 3214 7883
rect 2943 7884 2995 7885
rect 2997 7884 3014 7885
rect 3003 7886 3346 7887
rect 3018 7888 3391 7889
rect 3022 7890 3157 7891
rect 3025 7892 3269 7893
rect 3029 7894 3386 7895
rect 3032 7896 3332 7897
rect 3016 7898 3032 7899
rect 3037 7898 3541 7899
rect 3046 7900 3392 7901
rect 3049 7902 3236 7903
rect 3058 7904 3079 7905
rect 3060 7906 3065 7907
rect 3112 7906 3400 7907
rect 3120 7908 3328 7909
rect 3121 7910 3145 7911
rect 3126 7912 3134 7913
rect 3127 7914 3151 7915
rect 3139 7916 3644 7917
rect 3145 7918 3181 7919
rect 3157 7920 3211 7921
rect 3165 7922 3304 7923
rect 3172 7924 3217 7925
rect 3175 7926 3220 7927
rect 3184 7928 3241 7929
rect 3186 7930 3368 7931
rect 3189 7932 3376 7933
rect 3190 7934 3247 7935
rect 3193 7936 3250 7937
rect 3196 7938 3223 7939
rect 3201 7940 3485 7941
rect 3202 7942 3229 7943
rect 3205 7944 3238 7945
rect 3208 7946 3265 7947
rect 3211 7948 3274 7949
rect 3241 7950 3427 7951
rect 3247 7952 3310 7953
rect 3259 7954 3421 7955
rect 3265 7956 3352 7957
rect 3271 7958 3334 7959
rect 3277 7960 3298 7961
rect 3283 7962 3340 7963
rect 3252 7964 3341 7965
rect 3253 7966 3355 7967
rect 3286 7968 3343 7969
rect 3289 7970 3322 7971
rect 3291 7972 3647 7973
rect 3295 7974 3394 7975
rect 3301 7976 3358 7977
rect 3304 7978 3361 7979
rect 3307 7980 3364 7981
rect 3313 7982 3418 7983
rect 3319 7984 3382 7985
rect 3325 7986 3488 7987
rect 3337 7988 3388 7989
rect 3343 7990 3370 7991
rect 3349 7992 3536 7993
rect 3355 7994 3406 7995
rect 3358 7996 3409 7997
rect 3361 7998 3412 7999
rect 3364 8000 3415 8001
rect 3373 8002 3424 8003
rect 3388 8004 3442 8005
rect 3397 8006 3454 8007
rect 3403 8008 3460 8009
rect 3415 8010 3466 8011
rect 3429 8012 3654 8013
rect 3433 8014 3553 8015
rect 3316 8016 3553 8017
rect 3435 8018 3651 8019
rect 3436 8020 3556 8021
rect 3439 8022 3505 8023
rect 3447 8024 3640 8025
rect 3451 8026 3538 8027
rect 3454 8028 3675 8029
rect 3457 8030 3472 8031
rect 3460 8032 3595 8033
rect 3463 8034 3598 8035
rect 3466 8036 3526 8037
rect 3472 8038 3523 8039
rect 3475 8040 3634 8041
rect 3477 8042 3669 8043
rect 3478 8044 3571 8045
rect 3481 8046 3574 8047
rect 3490 8048 3643 8049
rect 3493 8050 3601 8051
rect 3495 8052 3573 8053
rect 3499 8054 3628 8055
rect 3502 8056 3604 8057
rect 3514 8058 3666 8059
rect 3516 8060 3734 8061
rect 3517 8062 3589 8063
rect 3520 8064 3663 8065
rect 3529 8066 3613 8067
rect 3532 8068 3616 8069
rect 3545 8070 3568 8071
rect 3549 8072 3660 8073
rect 3564 8074 3601 8075
rect 3575 8076 3678 8077
rect 3587 8078 3690 8079
rect 3591 8080 3713 8081
rect 3590 8082 3693 8083
rect 3618 8084 3741 8085
rect 3569 8086 3618 8087
rect 3624 8086 3717 8087
rect 3630 8088 3748 8089
rect 3645 8090 3667 8091
rect 3656 8092 3755 8093
rect 3671 8094 3706 8095
rect 3760 8094 3765 8095
rect 2921 8103 3209 8104
rect 2918 8105 2921 8106
rect 2927 8105 3305 8106
rect 2932 8107 3086 8108
rect 2931 8109 3146 8110
rect 2935 8111 3092 8112
rect 2954 8113 3104 8114
rect 2965 8115 3228 8116
rect 2975 8117 3107 8118
rect 2975 8119 2998 8120
rect 2987 8121 3272 8122
rect 2991 8123 3047 8124
rect 2990 8125 3284 8126
rect 2993 8127 3341 8128
rect 3003 8129 3007 8130
rect 3018 8129 3320 8130
rect 3018 8131 3308 8132
rect 3025 8133 3264 8134
rect 3027 8135 3189 8136
rect 3034 8137 3236 8138
rect 3041 8139 3219 8140
rect 3049 8141 3201 8142
rect 3056 8143 3059 8144
rect 3062 8143 3065 8144
rect 2925 8145 3066 8146
rect 3068 8145 3140 8146
rect 2961 8147 3141 8148
rect 3077 8149 3134 8150
rect 3080 8151 3137 8152
rect 3095 8153 3116 8154
rect 3097 8155 3246 8156
rect 3098 8157 3119 8158
rect 3101 8159 3122 8160
rect 3119 8161 3206 8162
rect 3127 8163 3539 8164
rect 3131 8165 3158 8166
rect 3134 8167 3173 8168
rect 3021 8169 3174 8170
rect 3021 8171 3032 8172
rect 3031 8173 3266 8174
rect 3143 8175 3176 8176
rect 3152 8177 3197 8178
rect 3158 8179 3185 8180
rect 3164 8181 3191 8182
rect 3167 8183 3194 8184
rect 3170 8185 3203 8186
rect 3182 8187 3212 8188
rect 3194 8189 3269 8190
rect 3212 8191 3248 8192
rect 3215 8193 3287 8194
rect 3224 8195 3254 8196
rect 3230 8197 3260 8198
rect 3236 8199 3278 8200
rect 3241 8201 3414 8202
rect 3242 8203 3302 8204
rect 3248 8205 3290 8206
rect 3254 8207 3296 8208
rect 3260 8209 3314 8210
rect 3266 8211 3326 8212
rect 3272 8213 3338 8214
rect 3275 8215 3536 8216
rect 3281 8217 3368 8218
rect 3287 8219 3356 8220
rect 3290 8221 3359 8222
rect 3293 8223 3362 8224
rect 3296 8225 3365 8226
rect 3299 8227 3374 8228
rect 3311 8229 3392 8230
rect 3316 8231 3420 8232
rect 3317 8233 3386 8234
rect 3320 8235 3389 8236
rect 3323 8237 3398 8238
rect 3329 8239 3404 8240
rect 3089 8241 3405 8242
rect 3341 8243 3471 8244
rect 3349 8245 3560 8246
rect 3359 8247 3434 8248
rect 3362 8249 3437 8250
rect 3365 8251 3440 8252
rect 3377 8253 3452 8254
rect 3386 8255 3455 8256
rect 3389 8257 3458 8258
rect 3343 8259 3459 8260
rect 3392 8261 3467 8262
rect 3331 8263 3468 8264
rect 3398 8265 3473 8266
rect 3401 8267 3476 8268
rect 3410 8269 3461 8270
rect 3415 8271 3523 8272
rect 3422 8273 3533 8274
rect 3425 8275 3500 8276
rect 3428 8277 3556 8278
rect 3437 8279 3515 8280
rect 3440 8281 3503 8282
rect 3449 8283 3479 8284
rect 3452 8285 3482 8286
rect 3455 8287 3482 8288
rect 3461 8289 3516 8290
rect 3463 8291 3532 8292
rect 3464 8293 3521 8294
rect 3474 8295 3530 8296
rect 3490 8297 3636 8298
rect 3493 8299 3553 8300
rect 3494 8301 3576 8302
rect 3506 8303 3588 8304
rect 3509 8305 3591 8306
rect 3517 8307 3604 8308
rect 3525 8309 3570 8310
rect 3528 8311 3573 8312
rect 3642 8311 3650 8312
rect 3645 8313 3660 8314
rect 2821 8322 2976 8323
rect 2917 8324 3022 8325
rect 2917 8326 3171 8327
rect 2924 8328 3066 8329
rect 2927 8330 3018 8331
rect 2931 8332 3168 8333
rect 2934 8334 3087 8335
rect 2953 8336 3075 8337
rect 2953 8338 3141 8339
rect 2969 8340 3132 8341
rect 2972 8342 2977 8343
rect 2979 8342 3099 8343
rect 2981 8344 3057 8345
rect 2988 8346 3063 8347
rect 2991 8348 3099 8349
rect 2997 8350 3078 8351
rect 2950 8352 3078 8353
rect 2950 8354 3075 8355
rect 3003 8356 3054 8357
rect 3002 8358 3414 8359
rect 3005 8360 3246 8361
rect 3008 8362 3102 8363
rect 3014 8364 3096 8365
rect 3024 8366 3081 8367
rect 3023 8368 3032 8369
rect 3032 8370 3135 8371
rect 3038 8372 3411 8373
rect 2960 8374 3039 8375
rect 3041 8374 3144 8375
rect 3044 8376 3159 8377
rect 3050 8378 3165 8379
rect 3056 8380 3120 8381
rect 3062 8382 3153 8383
rect 3068 8384 3405 8385
rect 3092 8386 3243 8387
rect 3095 8388 3183 8389
rect 3104 8390 3213 8391
rect 3107 8392 3216 8393
rect 3110 8394 3228 8395
rect 3089 8396 3229 8397
rect 3089 8398 3174 8399
rect 3113 8400 3151 8401
rect 3120 8402 3288 8403
rect 3123 8404 3273 8405
rect 3132 8406 3219 8407
rect 3138 8408 3225 8409
rect 3144 8410 3294 8411
rect 3153 8412 3195 8413
rect 3156 8414 3255 8415
rect 3162 8416 3300 8417
rect 3174 8418 3291 8419
rect 3183 8420 3231 8421
rect 3186 8422 3261 8423
rect 3188 8424 3417 8425
rect 3195 8426 3321 8427
rect 3200 8428 3523 8429
rect 3210 8430 3293 8431
rect 3213 8432 3237 8433
rect 3216 8434 3324 8435
rect 3234 8436 3366 8437
rect 3246 8438 3378 8439
rect 3189 8440 3377 8441
rect 3248 8442 3326 8443
rect 3249 8444 3399 8445
rect 3252 8446 3402 8447
rect 3255 8448 3360 8449
rect 3258 8450 3363 8451
rect 3263 8452 3420 8453
rect 3266 8454 3478 8455
rect 3267 8456 3345 8457
rect 3270 8458 3390 8459
rect 3273 8460 3297 8461
rect 3275 8462 3456 8463
rect 3276 8464 3408 8465
rect 3279 8466 3426 8467
rect 3281 8468 3338 8469
rect 3177 8470 3283 8471
rect 3295 8470 3423 8471
rect 3304 8472 3438 8473
rect 3307 8474 3441 8475
rect 3311 8476 3320 8477
rect 3317 8478 3475 8479
rect 3316 8480 3450 8481
rect 3329 8482 3482 8483
rect 3328 8484 3462 8485
rect 3331 8486 3465 8487
rect 3341 8488 3384 8489
rect 3358 8490 3516 8491
rect 3367 8492 3507 8493
rect 3370 8494 3510 8495
rect 3386 8496 3492 8497
rect 3386 8498 3526 8499
rect 3392 8500 3560 8501
rect 3406 8502 3529 8503
rect 3417 8504 3495 8505
rect 3428 8506 3563 8507
rect 3452 8508 3471 8509
rect 3548 8508 3553 8509
rect 2815 8517 2822 8518
rect 2881 8517 2892 8518
rect 2917 8517 3124 8518
rect 2920 8519 3042 8520
rect 2933 8521 3143 8522
rect 2941 8523 3108 8524
rect 2945 8525 3175 8526
rect 2952 8527 3075 8528
rect 2960 8529 3033 8530
rect 2962 8531 3078 8532
rect 2968 8533 3093 8534
rect 2972 8535 2994 8536
rect 2991 8537 3054 8538
rect 2990 8539 3015 8540
rect 2995 8541 3090 8542
rect 3002 8543 3018 8544
rect 2931 8545 3018 8546
rect 3005 8547 3154 8548
rect 3005 8549 3039 8550
rect 3008 8551 3024 8552
rect 3008 8553 3045 8554
rect 2998 8555 3045 8556
rect 2924 8557 3000 8558
rect 3014 8557 3051 8558
rect 3026 8559 3057 8560
rect 3032 8561 3063 8562
rect 3038 8563 3096 8564
rect 3041 8565 3087 8566
rect 3053 8567 3105 8568
rect 3056 8569 3099 8570
rect 3059 8571 3133 8572
rect 3062 8573 3184 8574
rect 3065 8575 3139 8576
rect 3068 8577 3271 8578
rect 3071 8579 3253 8580
rect 3074 8581 3145 8582
rect 3080 8583 3349 8584
rect 3086 8585 3157 8586
rect 3092 8587 3163 8588
rect 3101 8589 3335 8590
rect 3104 8591 3293 8592
rect 3107 8593 3187 8594
rect 3117 8595 3126 8596
rect 3116 8597 3277 8598
rect 3119 8599 3190 8600
rect 3122 8601 3342 8602
rect 3128 8603 3151 8604
rect 3132 8605 3178 8606
rect 3145 8607 3259 8608
rect 3151 8609 3320 8610
rect 3161 8611 3268 8612
rect 3167 8613 3329 8614
rect 3171 8615 3332 8616
rect 3174 8617 3217 8618
rect 3178 8619 3274 8620
rect 3184 8621 3280 8622
rect 3187 8623 3296 8624
rect 3190 8625 3317 8626
rect 3193 8627 3387 8628
rect 3195 8629 3345 8630
rect 3210 8631 3326 8632
rect 3213 8633 3323 8634
rect 3228 8635 3286 8636
rect 3234 8637 3384 8638
rect 3246 8639 3400 8640
rect 3249 8641 3381 8642
rect 3255 8643 3377 8644
rect 3304 8645 3390 8646
rect 3307 8647 3414 8648
rect 3367 8649 3421 8650
rect 3370 8651 3418 8652
rect 2884 8660 2892 8661
rect 2881 8662 2892 8663
rect 2882 8664 2889 8665
rect 2923 8664 3003 8665
rect 2930 8666 3015 8667
rect 2933 8668 3009 8669
rect 2942 8670 3000 8671
rect 2949 8672 2963 8673
rect 2956 8674 3039 8675
rect 2959 8676 3006 8677
rect 2965 8678 2991 8679
rect 2968 8680 3001 8681
rect 2972 8682 3045 8683
rect 2981 8684 3057 8685
rect 2993 8686 3042 8687
rect 2984 8688 2994 8689
rect 2984 8690 3027 8691
rect 2996 8692 3033 8693
rect 2987 8694 2998 8695
rect 3003 8694 3016 8695
rect 3006 8696 3075 8697
rect 3017 8698 3143 8699
rect 3018 8700 3129 8701
rect 3030 8702 3052 8703
rect 3042 8704 3120 8705
rect 3045 8706 3081 8707
rect 3053 8708 3072 8709
rect 3055 8710 3087 8711
rect 3059 8712 3066 8713
rect 3058 8714 3108 8715
rect 3092 8716 3140 8717
rect 3101 8718 3168 8719
rect 3104 8720 3126 8721
rect 3116 8722 3159 8723
rect 3122 8724 3165 8725
rect 3145 8726 3172 8727
rect 3161 8728 3188 8729
rect 3184 8730 3207 8731
rect 3193 8732 3200 8733
rect 2875 8741 2889 8742
rect 2882 8743 2892 8744
rect 2917 8743 2925 8744
rect 2962 8743 2966 8744
rect 2968 8743 3007 8744
rect 2971 8745 2982 8746
rect 2975 8747 2985 8748
rect 2987 8747 2994 8748
rect 2997 8747 3004 8748
rect 3012 8747 3031 8748
rect 3015 8749 3028 8750
rect 3018 8751 3056 8752
rect 3042 8753 3052 8754
rect 3045 8755 3049 8756
<< metal2 >>
rect 2941 1415 2942 1435
rect 2963 1415 2964 1435
rect 2944 1417 2945 1435
rect 3035 1417 3036 1435
rect 2947 1419 2948 1435
rect 2953 1419 2954 1435
rect 2957 1419 2958 1435
rect 2978 1419 2979 1435
rect 2960 1421 2961 1435
rect 2999 1421 3000 1435
rect 2966 1423 2967 1435
rect 3005 1423 3006 1435
rect 2984 1425 2985 1435
rect 3002 1425 3003 1435
rect 2987 1427 2988 1435
rect 2996 1427 2997 1435
rect 3011 1427 3012 1435
rect 3014 1427 3015 1435
rect 3017 1427 3018 1435
rect 3020 1427 3021 1435
rect 3026 1427 3027 1435
rect 3032 1427 3033 1435
rect 3044 1427 3045 1435
rect 3050 1427 3051 1435
rect 3047 1429 3048 1435
rect 3059 1429 3060 1435
rect 3056 1431 3057 1435
rect 3068 1431 3069 1435
rect 2809 1441 2810 1506
rect 3242 1441 3243 1506
rect 2938 1443 2939 1506
rect 2990 1443 2991 1506
rect 2944 1439 2945 1446
rect 3114 1445 3115 1506
rect 2947 1439 2948 1448
rect 2967 1447 2968 1506
rect 2953 1439 2954 1450
rect 2980 1449 2981 1506
rect 2973 1451 2974 1506
rect 3084 1451 3085 1506
rect 2978 1439 2979 1454
rect 3030 1453 3031 1506
rect 2984 1455 2985 1506
rect 3017 1439 3018 1456
rect 2987 1439 2988 1458
rect 3102 1457 3103 1506
rect 2987 1459 2988 1506
rect 3054 1459 3055 1506
rect 2993 1461 2994 1506
rect 3174 1461 3175 1506
rect 2996 1439 2997 1464
rect 3060 1463 3061 1506
rect 2999 1439 3000 1466
rect 3063 1465 3064 1506
rect 3000 1467 3001 1506
rect 3014 1439 3015 1468
rect 2950 1439 2951 1470
rect 3015 1469 3016 1506
rect 3002 1439 3003 1472
rect 3066 1471 3067 1506
rect 3005 1439 3006 1474
rect 3069 1473 3070 1506
rect 3011 1439 3012 1476
rect 3018 1475 3019 1506
rect 2963 1439 2964 1478
rect 3012 1477 3013 1506
rect 2952 1479 2953 1506
rect 2964 1479 2965 1506
rect 3023 1439 3024 1480
rect 3087 1479 3088 1506
rect 3026 1439 3027 1482
rect 3093 1481 3094 1506
rect 2931 1483 2932 1506
rect 3027 1483 3028 1506
rect 3035 1439 3036 1484
rect 3120 1483 3121 1506
rect 3036 1485 3037 1506
rect 3129 1485 3130 1506
rect 3039 1487 3040 1506
rect 3090 1487 3091 1506
rect 3044 1439 3045 1490
rect 3111 1489 3112 1506
rect 3047 1439 3048 1492
rect 3126 1491 3127 1506
rect 3056 1439 3057 1494
rect 3144 1493 3145 1506
rect 3150 1493 3151 1506
rect 3236 1493 3237 1506
rect 3153 1495 3154 1506
rect 3183 1495 3184 1506
rect 3156 1497 3157 1506
rect 3211 1497 3212 1506
rect 3165 1499 3166 1506
rect 3225 1499 3226 1506
rect 3177 1501 3178 1506
rect 3229 1501 3230 1506
rect 3190 1503 3191 1506
rect 3197 1503 3198 1506
rect 3204 1503 3205 1506
rect 3251 1503 3252 1506
rect 2920 1510 2921 1513
rect 2986 1512 2987 1631
rect 2920 1514 2921 1631
rect 2993 1510 2994 1515
rect 2936 1516 2937 1631
rect 3124 1516 3125 1631
rect 2938 1510 2939 1519
rect 3256 1518 3257 1631
rect 2934 1510 2935 1521
rect 2939 1520 2940 1631
rect 2933 1522 2934 1631
rect 2948 1510 2949 1523
rect 2917 1510 2918 1525
rect 2948 1524 2949 1631
rect 2941 1510 2942 1527
rect 3253 1526 3254 1631
rect 2955 1510 2956 1529
rect 3001 1528 3002 1631
rect 2809 1510 2810 1531
rect 2954 1530 2955 1631
rect 2957 1530 2958 1631
rect 3063 1510 3064 1531
rect 2924 1510 2925 1533
rect 3064 1532 3065 1631
rect 2960 1534 2961 1631
rect 3076 1534 3077 1631
rect 2964 1510 2965 1537
rect 2973 1510 2974 1537
rect 2970 1510 2971 1539
rect 3007 1538 3008 1631
rect 2971 1540 2972 1631
rect 3331 1540 3332 1631
rect 2990 1510 2991 1543
rect 3058 1542 3059 1631
rect 3015 1510 3016 1545
rect 3079 1544 3080 1631
rect 2967 1510 2968 1547
rect 3016 1546 3017 1631
rect 3018 1510 3019 1547
rect 3042 1546 3043 1631
rect 3025 1548 3026 1631
rect 3030 1510 3031 1549
rect 3035 1548 3036 1631
rect 3343 1548 3344 1631
rect 3046 1550 3047 1631
rect 3160 1550 3161 1631
rect 3069 1510 3070 1553
rect 3133 1552 3134 1631
rect 3072 1510 3073 1555
rect 3093 1510 3094 1555
rect 2984 1510 2985 1557
rect 3094 1556 3095 1631
rect 2917 1558 2918 1631
rect 2983 1558 2984 1631
rect 3084 1510 3085 1559
rect 3169 1558 3170 1631
rect 3087 1510 3088 1561
rect 3181 1560 3182 1631
rect 3102 1510 3103 1563
rect 3196 1562 3197 1631
rect 3111 1510 3112 1565
rect 3277 1564 3278 1631
rect 3114 1510 3115 1567
rect 3205 1566 3206 1631
rect 2931 1510 2932 1569
rect 3115 1568 3116 1631
rect 2930 1570 2931 1631
rect 3215 1510 3216 1571
rect 3120 1510 3121 1573
rect 3211 1572 3212 1631
rect 3027 1510 3028 1575
rect 3121 1574 3122 1631
rect 3126 1510 3127 1575
rect 3229 1574 3230 1631
rect 3032 1576 3033 1631
rect 3127 1576 3128 1631
rect 3129 1510 3130 1577
rect 3346 1576 3347 1631
rect 2977 1510 2978 1579
rect 3130 1578 3131 1631
rect 3141 1510 3142 1579
rect 3202 1578 3203 1631
rect 3142 1580 3143 1631
rect 3361 1580 3362 1631
rect 3144 1510 3145 1583
rect 3399 1582 3400 1631
rect 3054 1510 3055 1585
rect 3145 1584 3146 1631
rect 3150 1510 3151 1585
rect 3355 1584 3356 1631
rect 3066 1510 3067 1587
rect 3151 1586 3152 1631
rect 3153 1510 3154 1587
rect 3358 1586 3359 1631
rect 2998 1588 2999 1631
rect 3154 1588 3155 1631
rect 3156 1510 3157 1589
rect 3283 1588 3284 1631
rect 3060 1510 3061 1591
rect 3157 1590 3158 1631
rect 2902 1592 2903 1631
rect 3061 1592 3062 1631
rect 3162 1510 3163 1593
rect 3217 1592 3218 1631
rect 3165 1510 3166 1595
rect 3271 1594 3272 1631
rect 3174 1510 3175 1597
rect 3310 1596 3311 1631
rect 3175 1598 3176 1631
rect 3378 1598 3379 1631
rect 3177 1510 3178 1601
rect 3313 1600 3314 1631
rect 3178 1602 3179 1631
rect 3193 1602 3194 1631
rect 3183 1510 3184 1605
rect 3247 1604 3248 1631
rect 3090 1510 3091 1607
rect 3184 1606 3185 1631
rect 3012 1510 3013 1609
rect 3091 1608 3092 1631
rect 2974 1610 2975 1631
rect 3013 1610 3014 1631
rect 3187 1610 3188 1631
rect 3375 1610 3376 1631
rect 3222 1510 3223 1613
rect 3325 1612 3326 1631
rect 3225 1510 3226 1615
rect 3316 1614 3317 1631
rect 3236 1510 3237 1617
rect 3328 1616 3329 1631
rect 3241 1618 3242 1631
rect 3385 1618 3386 1631
rect 3259 1620 3260 1631
rect 3417 1620 3418 1631
rect 3274 1622 3275 1631
rect 3406 1622 3407 1631
rect 3295 1624 3296 1631
rect 3434 1624 3435 1631
rect 3319 1626 3320 1631
rect 3382 1626 3383 1631
rect 3322 1628 3323 1631
rect 3403 1628 3404 1631
rect 2894 1637 2895 1784
rect 3450 1637 3451 1784
rect 2917 1635 2918 1640
rect 2941 1639 2942 1784
rect 2933 1635 2934 1642
rect 2977 1641 2978 1784
rect 2932 1643 2933 1784
rect 3145 1635 3146 1644
rect 2944 1645 2945 1784
rect 2971 1635 2972 1646
rect 2930 1635 2931 1648
rect 2971 1647 2972 1784
rect 2954 1635 2955 1650
rect 3005 1649 3006 1784
rect 2948 1635 2949 1652
rect 2953 1651 2954 1784
rect 2974 1635 2975 1652
rect 3053 1651 3054 1784
rect 2881 1653 2882 1784
rect 2974 1653 2975 1784
rect 2983 1635 2984 1654
rect 3032 1653 3033 1784
rect 2990 1655 2991 1784
rect 3138 1655 3139 1784
rect 3010 1635 3011 1658
rect 3207 1657 3208 1784
rect 3011 1659 3012 1784
rect 3160 1635 3161 1660
rect 3035 1635 3036 1662
rect 3501 1661 3502 1784
rect 2986 1635 2987 1664
rect 3035 1663 3036 1784
rect 2987 1665 2988 1784
rect 3079 1635 3080 1666
rect 2929 1667 2930 1784
rect 3080 1667 3081 1784
rect 3039 1635 3040 1670
rect 3225 1669 3226 1784
rect 2922 1671 2923 1784
rect 3038 1671 3039 1784
rect 3041 1671 3042 1784
rect 3070 1635 3071 1672
rect 3007 1635 3008 1674
rect 3071 1673 3072 1784
rect 3046 1635 3047 1676
rect 3178 1635 3179 1676
rect 3049 1635 3050 1678
rect 3144 1677 3145 1784
rect 2902 1635 2903 1680
rect 3050 1679 3051 1784
rect 3058 1635 3059 1680
rect 3105 1679 3106 1784
rect 3013 1635 3014 1682
rect 3059 1681 3060 1784
rect 3001 1635 3002 1684
rect 3014 1683 3015 1784
rect 3061 1635 3062 1684
rect 3147 1683 3148 1784
rect 3016 1635 3017 1686
rect 3062 1685 3063 1784
rect 3064 1635 3065 1686
rect 3117 1685 3118 1784
rect 3083 1687 3084 1784
rect 3448 1635 3449 1688
rect 3124 1635 3125 1690
rect 3171 1689 3172 1784
rect 3076 1635 3077 1692
rect 3123 1691 3124 1784
rect 2915 1693 2916 1784
rect 3077 1693 3078 1784
rect 3130 1635 3131 1694
rect 3213 1693 3214 1784
rect 3151 1635 3152 1696
rect 3198 1695 3199 1784
rect 3089 1697 3090 1784
rect 3150 1697 3151 1784
rect 3175 1635 3176 1698
rect 3222 1697 3223 1784
rect 3127 1635 3128 1700
rect 3174 1699 3175 1784
rect 3184 1635 3185 1700
rect 3234 1699 3235 1784
rect 3190 1635 3191 1702
rect 3352 1635 3353 1702
rect 3142 1635 3143 1704
rect 3351 1703 3352 1784
rect 3094 1635 3095 1706
rect 3141 1705 3142 1784
rect 3093 1707 3094 1784
rect 3121 1635 3122 1708
rect 3193 1635 3194 1708
rect 3358 1635 3359 1708
rect 3202 1635 3203 1710
rect 3357 1709 3358 1784
rect 3154 1635 3155 1712
rect 3201 1711 3202 1784
rect 3205 1635 3206 1712
rect 3306 1711 3307 1784
rect 3157 1635 3158 1714
rect 3204 1713 3205 1784
rect 3211 1635 3212 1714
rect 3264 1713 3265 1784
rect 2998 1635 2999 1716
rect 3210 1715 3211 1784
rect 3229 1635 3230 1716
rect 3349 1635 3350 1716
rect 3181 1635 3182 1718
rect 3228 1717 3229 1784
rect 3133 1635 3134 1720
rect 3180 1719 3181 1784
rect 3091 1635 3092 1722
rect 3132 1721 3133 1784
rect 3187 1635 3188 1722
rect 3348 1721 3349 1784
rect 3025 1635 3026 1724
rect 3186 1723 3187 1784
rect 2925 1725 2926 1784
rect 3026 1725 3027 1784
rect 3231 1725 3232 1784
rect 3360 1725 3361 1784
rect 3247 1635 3248 1728
rect 3465 1727 3466 1784
rect 3196 1635 3197 1730
rect 3246 1729 3247 1784
rect 3253 1635 3254 1730
rect 3336 1729 3337 1784
rect 3256 1635 3257 1732
rect 3339 1731 3340 1784
rect 3271 1635 3272 1734
rect 3406 1635 3407 1734
rect 3270 1735 3271 1784
rect 3371 1635 3372 1736
rect 3274 1635 3275 1738
rect 3514 1737 3515 1784
rect 3283 1635 3284 1740
rect 3384 1739 3385 1784
rect 3295 1635 3296 1742
rect 3375 1741 3376 1784
rect 3217 1635 3218 1744
rect 3294 1743 3295 1784
rect 3028 1635 3029 1746
rect 3216 1745 3217 1784
rect 3300 1745 3301 1784
rect 3417 1635 3418 1746
rect 3310 1635 3311 1748
rect 3402 1747 3403 1784
rect 3313 1635 3314 1750
rect 3405 1749 3406 1784
rect 3312 1751 3313 1784
rect 3525 1751 3526 1784
rect 3316 1635 3317 1754
rect 3471 1753 3472 1784
rect 3315 1755 3316 1784
rect 3389 1635 3390 1756
rect 3319 1635 3320 1758
rect 3420 1757 3421 1784
rect 3255 1759 3256 1784
rect 3318 1759 3319 1784
rect 3322 1635 3323 1760
rect 3423 1759 3424 1784
rect 3325 1635 3326 1762
rect 3408 1761 3409 1784
rect 3241 1635 3242 1764
rect 3324 1763 3325 1784
rect 3073 1635 3074 1766
rect 3240 1765 3241 1784
rect 3331 1635 3332 1766
rect 3432 1765 3433 1784
rect 3343 1635 3344 1768
rect 3453 1767 3454 1784
rect 3259 1635 3260 1770
rect 3342 1769 3343 1784
rect 3346 1635 3347 1770
rect 3438 1769 3439 1784
rect 3355 1635 3356 1772
rect 3456 1771 3457 1784
rect 3354 1773 3355 1784
rect 3363 1773 3364 1784
rect 3372 1773 3373 1784
rect 3410 1635 3411 1774
rect 3328 1635 3329 1776
rect 3411 1775 3412 1784
rect 3378 1635 3379 1778
rect 3459 1777 3460 1784
rect 3277 1635 3278 1780
rect 3378 1779 3379 1784
rect 3276 1781 3277 1784
rect 3392 1635 3393 1782
rect 3468 1781 3469 1784
rect 3477 1781 3478 1784
rect 3552 1781 3553 1784
rect 3572 1781 3573 1784
rect 2863 1790 2864 1991
rect 2974 1788 2975 1791
rect 2866 1792 2867 1991
rect 2870 1792 2871 1991
rect 2884 1788 2885 1793
rect 2888 1788 2889 1793
rect 2894 1788 2895 1793
rect 2932 1788 2933 1793
rect 2901 1788 2902 1795
rect 3067 1794 3068 1991
rect 2904 1788 2905 1797
rect 3050 1788 3051 1797
rect 2914 1798 2915 1991
rect 3077 1788 3078 1799
rect 2918 1788 2919 1801
rect 3123 1788 3124 1801
rect 2922 1788 2923 1803
rect 3043 1802 3044 1991
rect 2925 1788 2926 1805
rect 3041 1788 3042 1805
rect 2928 1806 2929 1991
rect 3064 1806 3065 1991
rect 2953 1788 2954 1809
rect 2998 1808 2999 1991
rect 2959 1788 2960 1811
rect 3196 1810 3197 1991
rect 2962 1788 2963 1813
rect 2987 1788 2988 1813
rect 2968 1814 2969 1991
rect 3168 1788 3169 1815
rect 2971 1788 2972 1817
rect 2995 1816 2996 1991
rect 2983 1788 2984 1819
rect 3062 1788 3063 1819
rect 2990 1788 2991 1821
rect 3132 1788 3133 1821
rect 2989 1822 2990 1991
rect 3035 1788 3036 1823
rect 3007 1824 3008 1991
rect 3038 1788 3039 1825
rect 3014 1788 3015 1827
rect 3073 1826 3074 1991
rect 3026 1788 3027 1829
rect 3055 1828 3056 1991
rect 3032 1788 3033 1831
rect 3049 1830 3050 1991
rect 3005 1788 3006 1833
rect 3031 1832 3032 1991
rect 3004 1834 3005 1991
rect 3178 1834 3179 1991
rect 3034 1836 3035 1991
rect 3171 1788 3172 1837
rect 3053 1788 3054 1839
rect 3085 1838 3086 1991
rect 2941 1788 2942 1841
rect 3052 1840 3053 1991
rect 2940 1842 2941 1991
rect 3011 1788 3012 1843
rect 2977 1788 2978 1845
rect 3010 1844 3011 1991
rect 2977 1846 2978 1991
rect 3130 1846 3131 1991
rect 3059 1788 3060 1849
rect 3091 1848 3092 1991
rect 3061 1850 3062 1991
rect 3577 1850 3578 1991
rect 3080 1788 3081 1853
rect 3100 1852 3101 1991
rect 3079 1854 3080 1991
rect 3511 1788 3512 1855
rect 3089 1788 3090 1857
rect 3213 1788 3214 1857
rect 3096 1788 3097 1859
rect 3334 1858 3335 1991
rect 2917 1860 2918 1991
rect 3097 1860 3098 1991
rect 3111 1788 3112 1861
rect 3274 1860 3275 1991
rect 3136 1862 3137 1991
rect 3225 1788 3226 1863
rect 2911 1788 2912 1865
rect 3226 1864 3227 1991
rect 2910 1866 2911 1991
rect 3070 1866 3071 1991
rect 3138 1788 3139 1867
rect 3160 1866 3161 1991
rect 3141 1788 3142 1869
rect 3163 1868 3164 1991
rect 2897 1788 2898 1871
rect 3142 1870 3143 1991
rect 3144 1788 3145 1871
rect 3184 1870 3185 1991
rect 2903 1872 2904 1991
rect 3145 1872 3146 1991
rect 3166 1872 3167 1991
rect 3216 1788 3217 1873
rect 3169 1874 3170 1991
rect 3180 1788 3181 1875
rect 3174 1788 3175 1877
rect 3214 1876 3215 1991
rect 3186 1788 3187 1879
rect 3220 1878 3221 1991
rect 3190 1880 3191 1991
rect 3201 1788 3202 1881
rect 3112 1882 3113 1991
rect 3202 1882 3203 1991
rect 3204 1788 3205 1883
rect 3238 1882 3239 1991
rect 3210 1788 3211 1885
rect 3244 1884 3245 1991
rect 3222 1788 3223 1887
rect 3262 1886 3263 1991
rect 3231 1788 3232 1889
rect 3298 1888 3299 1991
rect 3198 1788 3199 1891
rect 3232 1890 3233 1991
rect 3147 1788 3148 1893
rect 3199 1892 3200 1991
rect 3117 1788 3118 1895
rect 3148 1894 3149 1991
rect 2921 1896 2922 1991
rect 3118 1896 3119 1991
rect 3234 1788 3235 1897
rect 3268 1896 3269 1991
rect 3235 1898 3236 1991
rect 3474 1788 3475 1899
rect 3240 1788 3241 1901
rect 3286 1900 3287 1991
rect 3207 1788 3208 1903
rect 3241 1902 3242 1991
rect 3109 1904 3110 1991
rect 3208 1904 3209 1991
rect 3246 1788 3247 1905
rect 3280 1904 3281 1991
rect 3150 1788 3151 1907
rect 3247 1906 3248 1991
rect 3255 1788 3256 1907
rect 3351 1788 3352 1907
rect 3264 1788 3265 1909
rect 3544 1908 3545 1991
rect 3016 1910 3017 1991
rect 3265 1910 3266 1991
rect 3270 1788 3271 1911
rect 3304 1910 3305 1991
rect 3276 1788 3277 1913
rect 3310 1912 3311 1991
rect 3294 1788 3295 1915
rect 3328 1914 3329 1991
rect 3300 1788 3301 1917
rect 3525 1788 3526 1917
rect 3114 1788 3115 1919
rect 3301 1918 3302 1991
rect 3083 1788 3084 1921
rect 3115 1920 3116 1991
rect 3306 1788 3307 1921
rect 3352 1920 3353 1991
rect 3322 1922 3323 1991
rect 3339 1788 3340 1923
rect 3312 1788 3313 1925
rect 3340 1924 3341 1991
rect 3324 1788 3325 1927
rect 3382 1926 3383 1991
rect 3336 1788 3337 1929
rect 3415 1928 3416 1991
rect 3348 1788 3349 1931
rect 3400 1930 3401 1991
rect 3354 1788 3355 1933
rect 3430 1932 3431 1991
rect 3370 1934 3371 1991
rect 3481 1788 3482 1935
rect 3384 1788 3385 1937
rect 3565 1936 3566 1991
rect 3402 1788 3403 1939
rect 3484 1938 3485 1991
rect 3318 1788 3319 1941
rect 3403 1940 3404 1991
rect 3405 1788 3406 1941
rect 3487 1940 3488 1991
rect 3408 1788 3409 1943
rect 3490 1942 3491 1991
rect 3411 1788 3412 1945
rect 3493 1944 3494 1991
rect 3412 1946 3413 1991
rect 3547 1946 3548 1991
rect 3420 1788 3421 1949
rect 3496 1948 3497 1991
rect 3375 1788 3376 1951
rect 3421 1950 3422 1991
rect 2896 1952 2897 1991
rect 3376 1952 3377 1991
rect 3423 1788 3424 1953
rect 3499 1952 3500 1991
rect 3342 1788 3343 1955
rect 3424 1954 3425 1991
rect 3315 1788 3316 1957
rect 3343 1956 3344 1991
rect 3438 1788 3439 1957
rect 3508 1956 3509 1991
rect 3448 1958 3449 1991
rect 3646 1958 3647 1991
rect 3450 1788 3451 1961
rect 3520 1960 3521 1991
rect 3372 1788 3373 1963
rect 3451 1962 3452 1991
rect 3453 1788 3454 1963
rect 3523 1962 3524 1991
rect 3378 1788 3379 1965
rect 3454 1964 3455 1991
rect 3456 1788 3457 1965
rect 3526 1964 3527 1991
rect 3459 1788 3460 1967
rect 3529 1966 3530 1991
rect 3468 1788 3469 1969
rect 3538 1968 3539 1991
rect 3471 1788 3472 1971
rect 3541 1970 3542 1991
rect 3552 1788 3553 1971
rect 3636 1970 3637 1991
rect 3418 1972 3419 1991
rect 3551 1972 3552 1991
rect 3558 1788 3559 1973
rect 3583 1972 3584 1991
rect 3228 1788 3229 1975
rect 3558 1974 3559 1991
rect 2980 1788 2981 1977
rect 3229 1976 3230 1991
rect 2980 1978 2981 1991
rect 3105 1788 3106 1979
rect 3562 1788 3563 1979
rect 3574 1978 3575 1991
rect 3572 1788 3573 1981
rect 3633 1980 3634 1991
rect 3501 1788 3502 1983
rect 3571 1982 3572 1991
rect 3432 1788 3433 1985
rect 3502 1984 3503 1991
rect 3357 1788 3358 1987
rect 3433 1986 3434 1991
rect 3358 1988 3359 1991
rect 3603 1988 3604 1991
rect 2866 1995 2867 1998
rect 3010 1995 3011 1998
rect 2896 1995 2897 2000
rect 3175 1999 3176 2212
rect 2903 1995 2904 2002
rect 2958 1995 2959 2002
rect 2870 1995 2871 2004
rect 2957 2003 2958 2212
rect 2902 2005 2903 2212
rect 3070 1995 3071 2006
rect 2909 2007 2910 2212
rect 3034 1995 3035 2008
rect 2915 2009 2916 2212
rect 3052 1995 3053 2010
rect 2921 1995 2922 2012
rect 3064 1995 3065 2012
rect 2924 1995 2925 2014
rect 3196 1995 3197 2014
rect 2934 2015 2935 2212
rect 3055 1995 3056 2016
rect 2940 1995 2941 2018
rect 3039 2017 3040 2212
rect 2961 1995 2962 2020
rect 3247 1995 3248 2020
rect 2960 2021 2961 2212
rect 3157 2021 3158 2212
rect 2963 2023 2964 2212
rect 3073 1995 3074 2024
rect 2966 2025 2967 2212
rect 2989 1995 2990 2026
rect 2968 1995 2969 2028
rect 3283 2027 3284 2212
rect 2972 2029 2973 2212
rect 2998 1995 2999 2030
rect 2977 1995 2978 2032
rect 3199 1995 3200 2032
rect 2984 2033 2985 2212
rect 3145 1995 3146 2034
rect 2995 1995 2996 2036
rect 3002 2035 3003 2212
rect 3005 2035 3006 2212
rect 3130 1995 3131 2036
rect 3016 1995 3017 2038
rect 3067 1995 3068 2038
rect 3017 2039 3018 2212
rect 3079 1995 3080 2040
rect 3020 2041 3021 2212
rect 3241 1995 3242 2042
rect 3023 2043 3024 2212
rect 3112 2043 3113 2212
rect 3025 1995 3026 2046
rect 3238 1995 3239 2046
rect 3028 1995 3029 2048
rect 3151 2047 3152 2212
rect 3033 2049 3034 2212
rect 3289 2049 3290 2212
rect 3036 2051 3037 2212
rect 3049 1995 3050 2052
rect 3043 1995 3044 2054
rect 3054 2053 3055 2212
rect 3031 1995 3032 2056
rect 3042 2055 3043 2212
rect 3030 2057 3031 2212
rect 3295 2057 3296 2212
rect 3051 2059 3052 2212
rect 3061 1995 3062 2060
rect 3070 2059 3071 2212
rect 3085 1995 3086 2060
rect 3076 2061 3077 2212
rect 3091 1995 3092 2062
rect 3100 1995 3101 2062
rect 3121 2061 3122 2212
rect 3109 1995 3110 2064
rect 3190 1995 3191 2064
rect 3118 1995 3119 2066
rect 3130 2065 3131 2212
rect 3097 1995 3098 2068
rect 3118 2067 3119 2212
rect 3124 2067 3125 2212
rect 3148 1995 3149 2068
rect 3142 1995 3143 2070
rect 3199 2069 3200 2212
rect 2931 2071 2932 2212
rect 3142 2071 3143 2212
rect 3160 1995 3161 2072
rect 3181 2071 3182 2212
rect 3166 1995 3167 2074
rect 3433 1995 3434 2074
rect 3169 1995 3170 2076
rect 3349 2075 3350 2212
rect 3169 2077 3170 2212
rect 3454 1995 3455 2078
rect 3178 1995 3179 2080
rect 3193 2079 3194 2212
rect 3115 1995 3116 2082
rect 3178 2081 3179 2212
rect 3184 1995 3185 2082
rect 3241 2081 3242 2212
rect 3163 1995 3164 2084
rect 3184 2083 3185 2212
rect 3139 1995 3140 2086
rect 3163 2085 3164 2212
rect 3187 2085 3188 2212
rect 3403 1995 3404 2086
rect 3202 1995 3203 2088
rect 3211 2087 3212 2212
rect 2900 1995 2901 2090
rect 3202 2089 3203 2212
rect 3208 1995 3209 2090
rect 3217 2089 3218 2212
rect 3226 1995 3227 2090
rect 3337 2089 3338 2212
rect 3232 1995 3233 2092
rect 3313 2091 3314 2212
rect 3235 1995 3236 2094
rect 3316 2093 3317 2212
rect 3220 1995 3221 2096
rect 3235 2095 3236 2212
rect 3244 1995 3245 2096
rect 3277 2095 3278 2212
rect 3244 2097 3245 2212
rect 3301 1995 3302 2098
rect 3250 1995 3251 2100
rect 3274 1995 3275 2100
rect 3250 2101 3251 2212
rect 3253 1995 3254 2102
rect 3253 2103 3254 2212
rect 3298 1995 3299 2104
rect 3214 1995 3215 2106
rect 3298 2105 3299 2212
rect 3256 2107 3257 2212
rect 3430 1995 3431 2108
rect 3262 1995 3263 2110
rect 3331 2109 3332 2212
rect 3265 1995 3266 2112
rect 3346 2111 3347 2212
rect 3268 1995 3269 2114
rect 3364 2113 3365 2212
rect 3286 1995 3287 2116
rect 3319 2115 3320 2212
rect 3307 2117 3308 2212
rect 3382 1995 3383 2118
rect 3280 1995 3281 2120
rect 3382 2119 3383 2212
rect 3310 1995 3311 2122
rect 3639 1995 3640 2122
rect 3322 1995 3323 2124
rect 3388 2123 3389 2212
rect 3340 1995 3341 2126
rect 3403 2125 3404 2212
rect 3229 1995 3230 2128
rect 3340 2127 3341 2212
rect 3229 2129 3230 2212
rect 3523 1995 3524 2130
rect 3343 1995 3344 2132
rect 3409 2131 3410 2212
rect 3103 2133 3104 2212
rect 3343 2133 3344 2212
rect 3352 1995 3353 2134
rect 3535 1995 3536 2134
rect 3358 1995 3359 2136
rect 3433 2135 3434 2212
rect 3328 1995 3329 2138
rect 3358 2137 3359 2212
rect 3367 2137 3368 2212
rect 3400 1995 3401 2138
rect 3376 1995 3377 2140
rect 3427 2139 3428 2212
rect 3376 2141 3377 2212
rect 3526 1995 3527 2142
rect 3379 2143 3380 2212
rect 3529 1995 3530 2144
rect 3385 2145 3386 2212
rect 3520 1995 3521 2146
rect 3400 2147 3401 2212
rect 3412 1995 3413 2148
rect 3418 1995 3419 2148
rect 3545 2147 3546 2212
rect 3418 2149 3419 2212
rect 3548 2149 3549 2212
rect 3424 1995 3425 2152
rect 3442 2151 3443 2212
rect 3439 2153 3440 2212
rect 3496 1995 3497 2154
rect 3448 1995 3449 2156
rect 3523 2155 3524 2212
rect 3415 1995 3416 2158
rect 3448 2157 3449 2212
rect 3415 2159 3416 2212
rect 3577 1995 3578 2160
rect 3445 2161 3446 2212
rect 3578 2161 3579 2212
rect 3481 2163 3482 2212
rect 3670 2163 3671 2212
rect 3484 1995 3485 2166
rect 3496 2165 3497 2212
rect 3451 1995 3452 2168
rect 3484 2167 3485 2212
rect 3451 2169 3452 2212
rect 3618 2169 3619 2212
rect 3490 1995 3491 2172
rect 3532 2171 3533 2212
rect 3421 1995 3422 2174
rect 3490 2173 3491 2212
rect 3370 1995 3371 2176
rect 3421 2175 3422 2212
rect 3304 1995 3305 2178
rect 3370 2177 3371 2212
rect 3493 1995 3494 2178
rect 3535 2177 3536 2212
rect 3493 2179 3494 2212
rect 3639 2179 3640 2212
rect 3499 1995 3500 2182
rect 3565 1995 3566 2182
rect 3487 1995 3488 2184
rect 3499 2183 3500 2212
rect 3502 1995 3503 2184
rect 3526 2183 3527 2212
rect 3508 1995 3509 2186
rect 3529 2185 3530 2212
rect 3514 2187 3515 2212
rect 3653 1995 3654 2188
rect 3520 2189 3521 2212
rect 3664 2189 3665 2212
rect 3538 1995 3539 2192
rect 3558 2191 3559 2212
rect 3325 2193 3326 2212
rect 3538 2193 3539 2212
rect 3555 2193 3556 2212
rect 3612 2193 3613 2212
rect 3561 1995 3562 2196
rect 3567 2195 3568 2212
rect 3541 1995 3542 2198
rect 3561 2197 3562 2212
rect 3265 2199 3266 2212
rect 3541 2199 3542 2212
rect 3571 1995 3572 2200
rect 3603 2199 3604 2212
rect 3574 1995 3575 2202
rect 3606 2201 3607 2212
rect 3583 1995 3584 2204
rect 3609 2203 3610 2212
rect 3591 2205 3592 2212
rect 3654 2205 3655 2212
rect 3633 1995 3634 2208
rect 3648 2207 3649 2212
rect 3636 1995 3637 2210
rect 3651 2209 3652 2212
rect 2899 2218 2900 2455
rect 2899 2216 2900 2219
rect 2902 2216 2903 2219
rect 3130 2216 3131 2219
rect 2915 2216 2916 2221
rect 3039 2216 3040 2221
rect 2924 2216 2925 2223
rect 3073 2222 3074 2455
rect 2923 2224 2924 2455
rect 3046 2224 3047 2455
rect 2927 2216 2928 2227
rect 3227 2226 3228 2455
rect 2927 2228 2928 2455
rect 3118 2216 3119 2229
rect 2934 2216 2935 2231
rect 3248 2230 3249 2455
rect 2933 2232 2934 2455
rect 2957 2216 2958 2233
rect 2961 2232 2962 2455
rect 2984 2216 2985 2233
rect 2964 2234 2965 2455
rect 3202 2216 3203 2235
rect 2966 2216 2967 2237
rect 3040 2236 3041 2455
rect 2972 2216 2973 2239
rect 2979 2238 2980 2455
rect 2985 2238 2986 2455
rect 3283 2216 3284 2239
rect 2988 2240 2989 2455
rect 3112 2216 3113 2241
rect 2993 2216 2994 2243
rect 3092 2242 3093 2455
rect 2992 2244 2993 2455
rect 3036 2216 3037 2245
rect 2920 2246 2921 2455
rect 3037 2246 3038 2455
rect 3004 2248 3005 2455
rect 3311 2248 3312 2455
rect 3007 2250 3008 2455
rect 3100 2216 3101 2251
rect 3020 2216 3021 2253
rect 3095 2252 3096 2455
rect 3017 2216 3018 2255
rect 3019 2254 3020 2455
rect 3002 2216 3003 2257
rect 3016 2256 3017 2455
rect 3023 2216 3024 2257
rect 3316 2216 3317 2257
rect 3030 2216 3031 2259
rect 3277 2216 3278 2259
rect 3031 2260 3032 2455
rect 3054 2216 3055 2261
rect 3042 2216 3043 2263
rect 3049 2262 3050 2455
rect 3043 2264 3044 2455
rect 3051 2216 3052 2265
rect 2906 2216 2907 2267
rect 3052 2266 3053 2455
rect 2906 2268 2907 2455
rect 3199 2216 3200 2269
rect 2967 2270 2968 2455
rect 3200 2270 3201 2455
rect 3060 2216 3061 2273
rect 3346 2216 3347 2273
rect 3061 2274 3062 2455
rect 3070 2216 3071 2275
rect 3067 2216 3068 2277
rect 3250 2216 3251 2277
rect 3067 2278 3068 2455
rect 3076 2216 3077 2279
rect 3076 2280 3077 2455
rect 3121 2216 3122 2281
rect 2995 2282 2996 2455
rect 3122 2282 3123 2455
rect 3079 2284 3080 2455
rect 3313 2216 3314 2285
rect 3098 2286 3099 2455
rect 3548 2286 3549 2455
rect 3103 2216 3104 2289
rect 3193 2216 3194 2289
rect 2902 2290 2903 2455
rect 3104 2290 3105 2455
rect 3116 2290 3117 2455
rect 3124 2216 3125 2291
rect 3128 2290 3129 2455
rect 3151 2216 3152 2291
rect 3140 2292 3141 2455
rect 3175 2216 3176 2293
rect 3142 2216 3143 2295
rect 3146 2294 3147 2455
rect 3143 2296 3144 2455
rect 3178 2216 3179 2297
rect 3157 2216 3158 2299
rect 3161 2298 3162 2455
rect 3169 2216 3170 2299
rect 3530 2298 3531 2455
rect 3173 2300 3174 2455
rect 3367 2216 3368 2301
rect 3176 2302 3177 2455
rect 3305 2302 3306 2455
rect 3179 2304 3180 2455
rect 3181 2216 3182 2305
rect 3182 2306 3183 2455
rect 3184 2216 3185 2307
rect 3187 2216 3188 2307
rect 3272 2306 3273 2455
rect 3197 2308 3198 2455
rect 3241 2216 3242 2309
rect 3203 2310 3204 2455
rect 3211 2216 3212 2311
rect 3163 2216 3164 2313
rect 3212 2312 3213 2455
rect 3209 2314 3210 2455
rect 3217 2216 3218 2315
rect 3215 2316 3216 2455
rect 3298 2216 3299 2317
rect 3229 2216 3230 2319
rect 3526 2216 3527 2319
rect 3233 2320 3234 2455
rect 3244 2216 3245 2321
rect 3239 2322 3240 2455
rect 3289 2216 3290 2323
rect 3245 2324 3246 2455
rect 3295 2216 3296 2325
rect 3251 2326 3252 2455
rect 3349 2216 3350 2327
rect 3256 2216 3257 2329
rect 3287 2328 3288 2455
rect 3088 2216 3089 2331
rect 3257 2330 3258 2455
rect 3089 2332 3090 2455
rect 3235 2216 3236 2333
rect 3236 2334 3237 2455
rect 3253 2216 3254 2335
rect 3263 2334 3264 2455
rect 3319 2216 3320 2335
rect 3265 2216 3266 2337
rect 3539 2336 3540 2455
rect 3275 2338 3276 2455
rect 3331 2216 3332 2339
rect 3281 2340 3282 2455
rect 3337 2216 3338 2341
rect 3284 2342 3285 2455
rect 3340 2216 3341 2343
rect 3290 2344 3291 2455
rect 3579 2344 3580 2455
rect 3296 2346 3297 2455
rect 3358 2216 3359 2347
rect 3302 2348 3303 2455
rect 3364 2216 3365 2349
rect 3307 2216 3308 2351
rect 3320 2350 3321 2455
rect 3325 2216 3326 2351
rect 3479 2350 3480 2455
rect 3326 2352 3327 2455
rect 3382 2216 3383 2353
rect 3332 2354 3333 2455
rect 3567 2216 3568 2355
rect 3338 2356 3339 2455
rect 3388 2216 3389 2357
rect 3343 2216 3344 2359
rect 3555 2216 3556 2359
rect 3350 2360 3351 2455
rect 3576 2360 3577 2455
rect 3353 2362 3354 2455
rect 3403 2216 3404 2363
rect 3359 2364 3360 2455
rect 3409 2216 3410 2365
rect 3365 2366 3366 2455
rect 3415 2216 3416 2367
rect 3370 2216 3371 2369
rect 3555 2368 3556 2455
rect 3371 2370 3372 2455
rect 3421 2216 3422 2371
rect 3379 2216 3380 2373
rect 3541 2216 3542 2373
rect 3383 2374 3384 2455
rect 3433 2216 3434 2375
rect 3385 2216 3386 2377
rect 3527 2376 3528 2455
rect 3392 2378 3393 2455
rect 3545 2216 3546 2379
rect 3400 2216 3401 2381
rect 3585 2216 3586 2381
rect 3401 2382 3402 2455
rect 3451 2216 3452 2383
rect 3057 2216 3058 2385
rect 3452 2384 3453 2455
rect 3437 2386 3438 2455
rect 3484 2216 3485 2387
rect 3439 2216 3440 2389
rect 3586 2388 3587 2455
rect 3442 2216 3443 2391
rect 3458 2390 3459 2455
rect 3445 2216 3446 2393
rect 3542 2392 3543 2455
rect 3448 2216 3449 2395
rect 3545 2394 3546 2455
rect 3418 2216 3419 2397
rect 3449 2396 3450 2455
rect 3455 2396 3456 2455
rect 3583 2396 3584 2455
rect 3473 2398 3474 2455
rect 3493 2216 3494 2399
rect 3476 2400 3477 2455
rect 3581 2216 3582 2401
rect 3481 2216 3482 2403
rect 3677 2216 3678 2403
rect 3485 2404 3486 2455
rect 3520 2216 3521 2405
rect 3490 2216 3491 2407
rect 3643 2406 3644 2455
rect 3496 2216 3497 2409
rect 3497 2408 3498 2455
rect 3499 2216 3500 2409
rect 3500 2408 3501 2455
rect 3503 2408 3504 2455
rect 3561 2216 3562 2409
rect 3509 2410 3510 2455
rect 3567 2410 3568 2455
rect 3514 2216 3515 2413
rect 3661 2216 3662 2413
rect 3521 2414 3522 2455
rect 3532 2216 3533 2415
rect 3523 2216 3524 2417
rect 3664 2216 3665 2417
rect 3524 2418 3525 2455
rect 3535 2216 3536 2419
rect 3376 2216 3377 2421
rect 3536 2420 3537 2455
rect 3377 2422 3378 2455
rect 3427 2216 3428 2423
rect 3533 2422 3534 2455
rect 3629 2422 3630 2455
rect 3558 2216 3559 2425
rect 3617 2424 3618 2455
rect 3314 2426 3315 2455
rect 3558 2426 3559 2455
rect 3564 2216 3565 2427
rect 3614 2426 3615 2455
rect 3571 2216 3572 2429
rect 3674 2216 3675 2429
rect 3488 2430 3489 2455
rect 3673 2430 3674 2455
rect 3573 2432 3574 2455
rect 3663 2432 3664 2455
rect 3603 2216 3604 2435
rect 3620 2434 3621 2455
rect 3602 2436 3603 2455
rect 3654 2216 3655 2437
rect 3606 2216 3607 2439
rect 3623 2438 3624 2455
rect 3591 2216 3592 2441
rect 3605 2440 3606 2455
rect 3609 2216 3610 2441
rect 3625 2216 3626 2441
rect 3608 2442 3609 2455
rect 3651 2216 3652 2443
rect 3425 2444 3426 2455
rect 3650 2444 3651 2455
rect 3612 2216 3613 2447
rect 3657 2216 3658 2447
rect 3611 2448 3612 2455
rect 3626 2448 3627 2455
rect 3636 2216 3637 2449
rect 3670 2448 3671 2455
rect 3308 2450 3309 2455
rect 3636 2450 3637 2455
rect 3648 2216 3649 2451
rect 3653 2450 3654 2455
rect 3413 2452 3414 2455
rect 3647 2452 3648 2455
rect 2894 2461 2895 2668
rect 3106 2461 3107 2668
rect 2899 2459 2900 2464
rect 2933 2459 2934 2464
rect 2901 2465 2902 2668
rect 3278 2465 3279 2668
rect 2904 2467 2905 2668
rect 3109 2467 3110 2668
rect 2906 2459 2907 2470
rect 3230 2469 3231 2668
rect 2913 2459 2914 2472
rect 3058 2471 3059 2668
rect 2916 2459 2917 2474
rect 3073 2459 3074 2474
rect 2918 2475 2919 2668
rect 3076 2459 3077 2476
rect 2934 2477 2935 2668
rect 3046 2459 3047 2478
rect 2943 2459 2944 2480
rect 3242 2479 3243 2668
rect 2951 2481 2952 2668
rect 2988 2459 2989 2482
rect 2955 2483 2956 2668
rect 3028 2483 3029 2668
rect 2992 2459 2993 2486
rect 3116 2459 3117 2486
rect 2995 2459 2996 2488
rect 3323 2487 3324 2668
rect 3010 2489 3011 2668
rect 3293 2489 3294 2668
rect 3013 2491 3014 2668
rect 3179 2459 3180 2492
rect 3016 2459 3017 2494
rect 3076 2493 3077 2668
rect 3019 2459 3020 2496
rect 3034 2495 3035 2668
rect 3022 2497 3023 2668
rect 3254 2497 3255 2668
rect 3037 2459 3038 2500
rect 3070 2499 3071 2668
rect 3043 2459 3044 2502
rect 3079 2501 3080 2668
rect 3052 2459 3053 2504
rect 3118 2503 3119 2668
rect 3061 2459 3062 2506
rect 3064 2505 3065 2668
rect 2974 2507 2975 2668
rect 3061 2507 3062 2668
rect 3095 2459 3096 2508
rect 3130 2507 3131 2668
rect 3094 2509 3095 2668
rect 3392 2459 3393 2510
rect 3101 2459 3102 2512
rect 3227 2459 3228 2512
rect 3104 2459 3105 2514
rect 3164 2513 3165 2668
rect 3049 2459 3050 2516
rect 3103 2515 3104 2668
rect 3128 2459 3129 2516
rect 3194 2515 3195 2668
rect 3092 2459 3093 2518
rect 3127 2517 3128 2668
rect 3146 2459 3147 2518
rect 3206 2517 3207 2668
rect 3152 2459 3153 2520
rect 3236 2459 3237 2520
rect 3091 2521 3092 2668
rect 3236 2521 3237 2668
rect 3158 2523 3159 2668
rect 3212 2459 3213 2524
rect 3161 2459 3162 2526
rect 3224 2525 3225 2668
rect 3170 2527 3171 2668
rect 3200 2459 3201 2528
rect 3140 2459 3141 2530
rect 3200 2529 3201 2668
rect 3140 2531 3141 2668
rect 3362 2531 3363 2668
rect 3188 2533 3189 2668
rect 3305 2459 3306 2534
rect 3212 2535 3213 2668
rect 3272 2459 3273 2536
rect 3197 2459 3198 2538
rect 3272 2537 3273 2668
rect 3182 2459 3183 2540
rect 3197 2539 3198 2668
rect 3233 2459 3234 2540
rect 3576 2459 3577 2540
rect 2964 2459 2965 2542
rect 3233 2541 3234 2668
rect 3248 2459 3249 2542
rect 3260 2541 3261 2668
rect 3266 2541 3267 2668
rect 3287 2459 3288 2542
rect 3281 2459 3282 2544
rect 3344 2543 3345 2668
rect 2927 2545 2928 2668
rect 3281 2545 3282 2668
rect 3284 2459 3285 2546
rect 3347 2545 3348 2668
rect 3203 2459 3204 2548
rect 3284 2547 3285 2668
rect 3143 2459 3144 2550
rect 3203 2549 3204 2668
rect 3143 2551 3144 2668
rect 3251 2459 3252 2552
rect 3296 2459 3297 2552
rect 3555 2459 3556 2552
rect 3215 2459 3216 2554
rect 3296 2553 3297 2668
rect 3302 2459 3303 2554
rect 3368 2553 3369 2668
rect 3086 2459 3087 2556
rect 3302 2555 3303 2668
rect 3067 2459 3068 2558
rect 3085 2557 3086 2668
rect 3308 2459 3309 2558
rect 3374 2557 3375 2668
rect 3257 2459 3258 2560
rect 3308 2559 3309 2668
rect 3314 2459 3315 2560
rect 3386 2559 3387 2668
rect 3239 2459 3240 2562
rect 3314 2561 3315 2668
rect 3320 2459 3321 2562
rect 3380 2561 3381 2668
rect 3245 2459 3246 2564
rect 3320 2563 3321 2668
rect 3031 2459 3032 2566
rect 3245 2565 3246 2668
rect 3326 2459 3327 2566
rect 3392 2565 3393 2668
rect 2985 2459 2986 2568
rect 3326 2567 3327 2668
rect 2961 2459 2962 2570
rect 2986 2569 2987 2668
rect 3332 2459 3333 2570
rect 3398 2569 3399 2668
rect 3290 2459 3291 2572
rect 3332 2571 3333 2668
rect 3209 2459 3210 2574
rect 3290 2573 3291 2668
rect 3004 2459 3005 2576
rect 3209 2575 3210 2668
rect 3004 2577 3005 2668
rect 3040 2459 3041 2578
rect 3338 2459 3339 2578
rect 3410 2577 3411 2668
rect 3263 2459 3264 2580
rect 3338 2579 3339 2668
rect 3350 2459 3351 2580
rect 3692 2579 3693 2668
rect 3275 2459 3276 2582
rect 3350 2581 3351 2668
rect 2915 2583 2916 2668
rect 3275 2583 3276 2668
rect 3353 2459 3354 2584
rect 3482 2583 3483 2668
rect 3356 2585 3357 2668
rect 3551 2459 3552 2586
rect 3365 2459 3366 2588
rect 3431 2587 3432 2668
rect 3371 2459 3372 2590
rect 3443 2589 3444 2668
rect 3176 2459 3177 2592
rect 3371 2591 3372 2668
rect 3122 2459 3123 2594
rect 3176 2593 3177 2668
rect 2979 2459 2980 2596
rect 3121 2595 3122 2668
rect 3401 2459 3402 2596
rect 3467 2595 3468 2668
rect 3416 2597 3417 2668
rect 3419 2597 3420 2668
rect 3422 2597 3423 2668
rect 3661 2597 3662 2668
rect 3425 2459 3426 2600
rect 3667 2599 3668 2668
rect 3359 2459 3360 2602
rect 3425 2601 3426 2668
rect 3452 2459 3453 2602
rect 3593 2459 3594 2602
rect 3458 2459 3459 2604
rect 3506 2603 3507 2668
rect 3479 2459 3480 2606
rect 3515 2605 3516 2668
rect 3449 2459 3450 2608
rect 3479 2607 3480 2668
rect 3485 2459 3486 2608
rect 3551 2607 3552 2668
rect 3413 2459 3414 2610
rect 3485 2609 3486 2668
rect 3488 2459 3489 2610
rect 3554 2609 3555 2668
rect 3497 2459 3498 2612
rect 3611 2459 3612 2612
rect 3500 2459 3501 2614
rect 3608 2459 3609 2614
rect 3509 2459 3510 2616
rect 3557 2615 3558 2668
rect 3437 2459 3438 2618
rect 3509 2617 3510 2668
rect 3521 2459 3522 2618
rect 3578 2617 3579 2668
rect 3524 2459 3525 2620
rect 3581 2619 3582 2668
rect 3527 2459 3528 2622
rect 3563 2621 3564 2668
rect 3533 2459 3534 2624
rect 3656 2459 3657 2624
rect 3545 2459 3546 2626
rect 3567 2459 3568 2626
rect 3503 2459 3504 2628
rect 3545 2627 3546 2668
rect 3455 2459 3456 2630
rect 3503 2629 3504 2668
rect 3383 2459 3384 2632
rect 3455 2631 3456 2668
rect 3530 2459 3531 2632
rect 3566 2631 3567 2668
rect 3569 2631 3570 2668
rect 3586 2459 3587 2632
rect 3536 2459 3537 2634
rect 3587 2633 3588 2668
rect 3573 2459 3574 2636
rect 3637 2635 3638 2668
rect 3377 2459 3378 2638
rect 3572 2637 3573 2668
rect 3311 2459 3312 2640
rect 3377 2639 3378 2668
rect 3575 2639 3576 2668
rect 3743 2639 3744 2668
rect 3584 2641 3585 2668
rect 3590 2459 3591 2642
rect 3539 2459 3540 2644
rect 3590 2643 3591 2668
rect 3473 2459 3474 2646
rect 3539 2645 3540 2668
rect 3599 2645 3600 2668
rect 3650 2459 3651 2646
rect 3605 2459 3606 2648
rect 3655 2647 3656 2668
rect 3329 2649 3330 2668
rect 3605 2649 3606 2668
rect 3617 2459 3618 2650
rect 3679 2649 3680 2668
rect 3404 2651 3405 2668
rect 3617 2651 3618 2668
rect 3620 2459 3621 2652
rect 3664 2651 3665 2668
rect 3623 2459 3624 2654
rect 3647 2459 3648 2654
rect 3542 2459 3543 2656
rect 3624 2655 3625 2668
rect 3476 2459 3477 2658
rect 3542 2657 3543 2668
rect 3653 2459 3654 2658
rect 3695 2657 3696 2668
rect 3602 2459 3603 2660
rect 3652 2659 3653 2668
rect 3602 2661 3603 2668
rect 3640 2661 3641 2668
rect 3670 2661 3671 2668
rect 3689 2661 3690 2668
rect 3677 2459 3678 2664
rect 3733 2663 3734 2668
rect 3614 2459 3615 2666
rect 3676 2665 3677 2668
rect 2890 2672 2891 2675
rect 3200 2672 3201 2675
rect 2897 2672 2898 2677
rect 3109 2672 3110 2677
rect 2905 2678 2906 2925
rect 3133 2678 3134 2925
rect 2915 2672 2916 2681
rect 3006 2680 3007 2925
rect 2931 2682 2932 2925
rect 3070 2672 3071 2683
rect 2934 2684 2935 2925
rect 3281 2672 3282 2685
rect 2908 2672 2909 2687
rect 3280 2686 3281 2925
rect 2937 2672 2938 2689
rect 2967 2672 2968 2689
rect 2941 2672 2942 2691
rect 3206 2672 3207 2691
rect 2944 2672 2945 2693
rect 3268 2692 3269 2925
rect 2943 2694 2944 2925
rect 2948 2672 2949 2695
rect 2946 2696 2947 2925
rect 3209 2672 3210 2697
rect 2965 2698 2966 2925
rect 3433 2698 3434 2925
rect 2974 2672 2975 2701
rect 3197 2672 3198 2701
rect 2976 2702 2977 2925
rect 3194 2672 3195 2703
rect 2986 2672 2987 2705
rect 3018 2704 3019 2925
rect 2997 2706 2998 2925
rect 3212 2672 3213 2707
rect 3004 2672 3005 2709
rect 3358 2708 3359 2925
rect 3028 2672 3029 2711
rect 3055 2710 3056 2925
rect 3027 2712 3028 2925
rect 3158 2672 3159 2713
rect 3034 2672 3035 2715
rect 3049 2714 3050 2925
rect 3036 2716 3037 2925
rect 3064 2672 3065 2717
rect 3046 2718 3047 2925
rect 3302 2672 3303 2719
rect 3061 2672 3062 2721
rect 3088 2720 3089 2925
rect 3073 2722 3074 2925
rect 3245 2672 3246 2723
rect 3076 2672 3077 2725
rect 3112 2724 3113 2925
rect 3079 2672 3080 2727
rect 3097 2726 3098 2925
rect 3079 2728 3080 2925
rect 3109 2728 3110 2925
rect 3082 2730 3083 2925
rect 3314 2672 3315 2731
rect 3085 2672 3086 2733
rect 3091 2732 3092 2925
rect 3058 2672 3059 2735
rect 3085 2734 3086 2925
rect 3094 2672 3095 2735
rect 3136 2672 3137 2735
rect 3103 2672 3104 2737
rect 3148 2736 3149 2925
rect 3103 2738 3104 2925
rect 3460 2738 3461 2925
rect 3106 2672 3107 2741
rect 3121 2740 3122 2925
rect 3106 2742 3107 2925
rect 3266 2672 3267 2743
rect 3115 2744 3116 2925
rect 3127 2672 3128 2745
rect 3124 2672 3125 2747
rect 3308 2672 3309 2747
rect 3140 2672 3141 2749
rect 3617 2672 3618 2749
rect 3151 2750 3152 2925
rect 3188 2672 3189 2751
rect 3022 2672 3023 2753
rect 3187 2752 3188 2925
rect 3164 2672 3165 2755
rect 3181 2754 3182 2925
rect 3170 2672 3171 2757
rect 3205 2756 3206 2925
rect 3176 2672 3177 2759
rect 3193 2758 3194 2925
rect 3199 2758 3200 2925
rect 3566 2672 3567 2759
rect 3217 2760 3218 2925
rect 3254 2672 3255 2761
rect 3224 2672 3225 2763
rect 3244 2762 3245 2925
rect 2979 2764 2980 2925
rect 3223 2764 3224 2925
rect 3230 2672 3231 2765
rect 3298 2764 3299 2925
rect 3229 2766 3230 2925
rect 3515 2672 3516 2767
rect 3233 2672 3234 2769
rect 3301 2768 3302 2925
rect 3236 2672 3237 2771
rect 3250 2770 3251 2925
rect 3203 2672 3204 2773
rect 3235 2772 3236 2925
rect 3238 2772 3239 2925
rect 3590 2672 3591 2773
rect 3242 2672 3243 2775
rect 3286 2774 3287 2925
rect 3256 2776 3257 2925
rect 3326 2672 3327 2777
rect 3262 2778 3263 2925
rect 3404 2672 3405 2779
rect 3275 2672 3276 2781
rect 3325 2780 3326 2925
rect 3260 2672 3261 2783
rect 3274 2782 3275 2925
rect 3259 2784 3260 2925
rect 3329 2672 3330 2785
rect 2969 2786 2970 2925
rect 3328 2786 3329 2925
rect 3284 2672 3285 2789
rect 3316 2788 3317 2925
rect 3293 2672 3294 2791
rect 3334 2790 3335 2925
rect 3292 2792 3293 2925
rect 3587 2672 3588 2793
rect 3296 2672 3297 2795
rect 3310 2794 3311 2925
rect 3323 2672 3324 2795
rect 3394 2794 3395 2925
rect 3272 2672 3273 2797
rect 3322 2796 3323 2925
rect 3332 2672 3333 2797
rect 3620 2672 3621 2797
rect 3290 2672 3291 2799
rect 3331 2798 3332 2925
rect 2915 2800 2916 2925
rect 3289 2800 3290 2925
rect 3344 2672 3345 2801
rect 3427 2800 3428 2925
rect 3356 2672 3357 2803
rect 3687 2802 3688 2925
rect 3278 2672 3279 2805
rect 3355 2804 3356 2925
rect 3368 2672 3369 2805
rect 3451 2804 3452 2925
rect 3367 2806 3368 2925
rect 3661 2672 3662 2807
rect 3374 2672 3375 2809
rect 3463 2808 3464 2925
rect 3362 2672 3363 2811
rect 3373 2810 3374 2925
rect 3380 2672 3381 2811
rect 3403 2810 3404 2925
rect 2950 2812 2951 2925
rect 3379 2812 3380 2925
rect 3386 2672 3387 2813
rect 3457 2812 3458 2925
rect 3160 2814 3161 2925
rect 3385 2814 3386 2925
rect 3398 2672 3399 2815
rect 3487 2814 3488 2925
rect 3397 2816 3398 2925
rect 3605 2672 3606 2817
rect 3410 2672 3411 2819
rect 3662 2818 3663 2925
rect 3409 2820 3410 2925
rect 3754 2820 3755 2925
rect 3425 2672 3426 2823
rect 3517 2822 3518 2925
rect 3431 2672 3432 2825
rect 3523 2824 3524 2925
rect 3347 2672 3348 2827
rect 3430 2826 3431 2925
rect 3439 2826 3440 2925
rect 3672 2826 3673 2925
rect 3443 2672 3444 2829
rect 3493 2828 3494 2925
rect 2972 2830 2973 2925
rect 3442 2830 3443 2925
rect 3455 2672 3456 2831
rect 3547 2830 3548 2925
rect 3371 2672 3372 2833
rect 3454 2832 3455 2925
rect 3467 2672 3468 2833
rect 3559 2832 3560 2925
rect 3377 2672 3378 2835
rect 3466 2834 3467 2925
rect 3475 2834 3476 2925
rect 3624 2672 3625 2835
rect 3479 2672 3480 2837
rect 3691 2836 3692 2925
rect 3482 2672 3483 2839
rect 3658 2672 3659 2839
rect 3392 2672 3393 2841
rect 3481 2840 3482 2925
rect 3320 2672 3321 2843
rect 3391 2842 3392 2925
rect 3415 2842 3416 2925
rect 3658 2842 3659 2925
rect 3490 2844 3491 2925
rect 3563 2672 3564 2845
rect 3496 2846 3497 2925
rect 3503 2672 3504 2847
rect 3499 2848 3500 2925
rect 3557 2672 3558 2849
rect 3506 2672 3507 2851
rect 3640 2672 3641 2851
rect 3505 2852 3506 2925
rect 3631 2672 3632 2853
rect 3509 2672 3510 2855
rect 3595 2854 3596 2925
rect 3422 2672 3423 2857
rect 3508 2856 3509 2925
rect 3350 2672 3351 2859
rect 3421 2858 3422 2925
rect 2922 2860 2923 2925
rect 3349 2860 3350 2925
rect 3526 2860 3527 2925
rect 3684 2860 3685 2925
rect 3529 2862 3530 2925
rect 3572 2672 3573 2863
rect 3485 2672 3486 2865
rect 3571 2864 3572 2925
rect 3532 2866 3533 2925
rect 3569 2672 3570 2867
rect 3535 2868 3536 2925
rect 3545 2672 3546 2869
rect 3539 2672 3540 2871
rect 3607 2870 3608 2925
rect 3542 2672 3543 2873
rect 3610 2872 3611 2925
rect 3541 2874 3542 2925
rect 3682 2672 3683 2875
rect 3551 2672 3552 2877
rect 3625 2876 3626 2925
rect 3554 2672 3555 2879
rect 3628 2878 3629 2925
rect 3565 2880 3566 2925
rect 3581 2672 3582 2881
rect 3575 2672 3576 2883
rect 3768 2882 3769 2925
rect 3578 2672 3579 2885
rect 3640 2884 3641 2925
rect 3589 2886 3590 2925
rect 3599 2672 3600 2887
rect 3592 2888 3593 2925
rect 3602 2672 3603 2889
rect 3652 2672 3653 2889
rect 3681 2888 3682 2925
rect 3655 2672 3656 2891
rect 3718 2890 3719 2925
rect 3338 2672 3339 2893
rect 3655 2892 3656 2925
rect 3039 2894 3040 2925
rect 3337 2894 3338 2925
rect 3676 2672 3677 2895
rect 3712 2894 3713 2925
rect 3679 2672 3680 2897
rect 3715 2896 3716 2925
rect 3584 2672 3585 2899
rect 3678 2898 3679 2925
rect 3583 2900 3584 2925
rect 3667 2672 3668 2901
rect 3689 2672 3690 2901
rect 3758 2900 3759 2925
rect 3695 2672 3696 2903
rect 3738 2902 3739 2925
rect 3708 2672 3709 2905
rect 3726 2672 3727 2905
rect 3637 2672 3638 2907
rect 3709 2906 3710 2925
rect 3637 2908 3638 2925
rect 3698 2672 3699 2909
rect 3664 2672 3665 2911
rect 3697 2910 3698 2925
rect 3361 2912 3362 2925
rect 3665 2912 3666 2925
rect 3729 2672 3730 2913
rect 3736 2672 3737 2913
rect 3601 2914 3602 2925
rect 3735 2914 3736 2925
rect 3675 2916 3676 2925
rect 3728 2916 3729 2925
rect 3733 2672 3734 2917
rect 3786 2916 3787 2925
rect 3740 2672 3741 2919
rect 3747 2672 3748 2919
rect 3700 2920 3701 2925
rect 3747 2920 3748 2925
rect 3741 2922 3742 2925
rect 3772 2922 3773 2925
rect 2914 2931 2915 3154
rect 3085 2929 3086 2932
rect 2931 2929 2932 2934
rect 3286 2929 3287 2934
rect 2950 2929 2951 2936
rect 3363 2935 3364 3154
rect 2953 2929 2954 2938
rect 3358 2929 3359 2938
rect 2962 2929 2963 2940
rect 3073 2929 3074 2940
rect 2934 2929 2935 2942
rect 3072 2941 3073 3154
rect 2921 2943 2922 3154
rect 2933 2943 2934 3154
rect 2961 2943 2962 3154
rect 2994 2929 2995 2944
rect 2971 2945 2972 3154
rect 3427 2929 3428 2946
rect 2976 2929 2977 2948
rect 3193 2929 3194 2948
rect 2993 2949 2994 3154
rect 3468 2949 3469 3154
rect 3006 2929 3007 2952
rect 3029 2951 3030 3154
rect 3014 2953 3015 3154
rect 3244 2929 3245 2954
rect 3018 2929 3019 2956
rect 3023 2955 3024 3154
rect 3027 2929 3028 2956
rect 3187 2929 3188 2956
rect 3043 2929 3044 2958
rect 3421 2929 3422 2958
rect 3045 2959 3046 3154
rect 3162 2959 3163 3154
rect 3048 2961 3049 3154
rect 3049 2929 3050 2962
rect 3055 2929 3056 2962
rect 3060 2961 3061 3154
rect 3069 2961 3070 3154
rect 3103 2929 3104 2962
rect 3079 2929 3080 2964
rect 3303 2963 3304 3154
rect 2979 2929 2980 2966
rect 3078 2965 3079 3154
rect 2978 2967 2979 3154
rect 3379 2929 3380 2968
rect 3087 2969 3088 3154
rect 3088 2929 3089 2970
rect 3097 2929 3098 2970
rect 3099 2969 3100 3154
rect 3096 2971 3097 3154
rect 3112 2929 3113 2972
rect 3091 2929 3092 2974
rect 3111 2973 3112 3154
rect 3106 2929 3107 2976
rect 3259 2929 3260 2976
rect 3109 2929 3110 2978
rect 3123 2977 3124 3154
rect 3115 2929 3116 2980
rect 3144 2979 3145 3154
rect 3126 2981 3127 3154
rect 3148 2929 3149 2982
rect 3118 2929 3119 2984
rect 3147 2983 3148 3154
rect 3117 2985 3118 3154
rect 3475 2929 3476 2986
rect 3130 2929 3131 2988
rect 3138 2987 3139 3154
rect 3121 2929 3122 2990
rect 3129 2989 3130 3154
rect 3120 2991 3121 3154
rect 3378 2991 3379 3154
rect 3133 2929 3134 2994
rect 3141 2993 3142 3154
rect 3151 2929 3152 2994
rect 3174 2993 3175 3154
rect 3157 2929 3158 2996
rect 3238 2929 3239 2996
rect 3160 2929 3161 2998
rect 3373 2929 3374 2998
rect 3181 2929 3182 3000
rect 3186 2999 3187 3154
rect 3180 3001 3181 3154
rect 3442 2929 3443 3002
rect 3210 3003 3211 3154
rect 3223 2929 3224 3004
rect 3222 3005 3223 3154
rect 3229 2929 3230 3006
rect 3228 3007 3229 3154
rect 3250 2929 3251 3008
rect 2899 3009 2900 3154
rect 3249 3009 3250 3154
rect 3234 3011 3235 3154
rect 3235 2929 3236 3012
rect 3237 3011 3238 3154
rect 3765 2929 3766 3012
rect 3240 3013 3241 3154
rect 3262 2929 3263 3014
rect 3246 3015 3247 3154
rect 3256 2929 3257 3016
rect 3255 3017 3256 3154
rect 3274 2929 3275 3018
rect 3261 3019 3262 3154
rect 3658 2929 3659 3020
rect 3268 2929 3269 3022
rect 3273 3021 3274 3154
rect 3267 3023 3268 3154
rect 3310 2929 3311 3024
rect 3038 3025 3039 3154
rect 3309 3025 3310 3154
rect 3280 2929 3281 3028
rect 3285 3027 3286 3154
rect 3279 3029 3280 3154
rect 3316 2929 3317 3030
rect 3288 3031 3289 3154
rect 3289 2929 3290 3032
rect 3292 2929 3293 3032
rect 3357 3031 3358 3154
rect 3291 3033 3292 3154
rect 3298 2929 3299 3034
rect 2975 3035 2976 3154
rect 3297 3035 3298 3154
rect 3294 3037 3295 3154
rect 3301 2929 3302 3038
rect 3312 3037 3313 3154
rect 3430 2929 3431 3038
rect 3315 3039 3316 3154
rect 3331 2929 3332 3040
rect 3318 3041 3319 3154
rect 3334 2929 3335 3042
rect 3325 2929 3326 3044
rect 3369 3043 3370 3154
rect 2943 2929 2944 3046
rect 3324 3045 3325 3154
rect 3333 3045 3334 3154
rect 3337 2929 3338 3046
rect 3349 2929 3350 3046
rect 3351 3045 3352 3154
rect 3372 3045 3373 3154
rect 3685 3045 3686 3154
rect 3384 3047 3385 3154
rect 3385 2929 3386 3048
rect 3390 3047 3391 3154
rect 3391 2929 3392 3048
rect 3393 3047 3394 3154
rect 3394 2929 3395 3048
rect 3403 2929 3404 3048
rect 3660 3047 3661 3154
rect 3397 2929 3398 3050
rect 3402 3049 3403 3154
rect 2912 2929 2913 3052
rect 3396 3051 3397 3154
rect 2911 3053 2912 3154
rect 3084 3053 3085 3154
rect 3409 2929 3410 3054
rect 3420 3053 3421 3154
rect 3367 2929 3368 3056
rect 3408 3055 3409 3154
rect 2965 2929 2966 3058
rect 3366 3057 3367 3154
rect 2964 3059 2965 3154
rect 3205 2929 3206 3060
rect 3415 2929 3416 3060
rect 3426 3059 3427 3154
rect 3439 2929 3440 3060
rect 3444 3059 3445 3154
rect 3361 2929 3362 3062
rect 3438 3061 3439 3154
rect 3454 2929 3455 3062
rect 3483 3061 3484 3154
rect 2946 2929 2947 3064
rect 3453 3063 3454 3154
rect 3466 2929 3467 3064
rect 3471 3063 3472 3154
rect 3460 2929 3461 3066
rect 3465 3065 3466 3154
rect 3499 2929 3500 3066
rect 3756 3065 3757 3154
rect 3505 2929 3506 3068
rect 3510 3067 3511 3154
rect 3493 2929 3494 3070
rect 3504 3069 3505 3154
rect 3487 2929 3488 3072
rect 3492 3071 3493 3154
rect 3481 2929 3482 3074
rect 3486 3073 3487 3154
rect 3082 2929 3083 3076
rect 3480 3075 3481 3154
rect 3508 2929 3509 3076
rect 3513 3075 3514 3154
rect 3496 2929 3497 3078
rect 3507 3077 3508 3154
rect 3490 2929 3491 3080
rect 3495 3079 3496 3154
rect 3535 2929 3536 3080
rect 3728 2929 3729 3080
rect 3523 2929 3524 3082
rect 3534 3081 3535 3154
rect 3517 2929 3518 3084
rect 3522 3083 3523 3154
rect 3433 2929 3434 3086
rect 3516 3085 3517 3154
rect 3432 3087 3433 3154
rect 3451 2929 3452 3088
rect 3450 3089 3451 3154
rect 3669 2929 3670 3090
rect 3541 2929 3542 3092
rect 3687 2929 3688 3092
rect 3526 2929 3527 3094
rect 3540 3093 3541 3154
rect 3543 3093 3544 3154
rect 3691 2929 3692 3094
rect 3585 3095 3586 3154
rect 3703 2929 3704 3096
rect 3589 2929 3590 3098
rect 3621 3097 3622 3154
rect 3571 2929 3572 3100
rect 3588 3099 3589 3154
rect 3559 2929 3560 3102
rect 3570 3101 3571 3154
rect 3547 2929 3548 3104
rect 3558 3103 3559 3154
rect 3529 2929 3530 3106
rect 3546 3105 3547 3154
rect 3528 3107 3529 3154
rect 3727 3107 3728 3154
rect 3595 2929 3596 3110
rect 3615 3109 3616 3154
rect 3610 2929 3611 3112
rect 3630 3111 3631 3154
rect 3612 3113 3613 3154
rect 3796 2929 3797 3114
rect 3625 2929 3626 3116
rect 3791 3115 3792 3154
rect 3592 2929 3593 3118
rect 3624 3117 3625 3154
rect 3628 2929 3629 3118
rect 3793 2929 3794 3118
rect 3607 2929 3608 3120
rect 3627 3119 3628 3154
rect 3565 2929 3566 3122
rect 3606 3121 3607 3154
rect 3637 2929 3638 3122
rect 3746 3121 3747 3154
rect 3640 2929 3641 3124
rect 3645 3123 3646 3154
rect 3657 3123 3658 3154
rect 3749 3123 3750 3154
rect 3669 3125 3670 3154
rect 3779 2929 3780 3126
rect 3601 2929 3602 3128
rect 3778 3127 3779 3154
rect 3583 2929 3584 3130
rect 3600 3129 3601 3154
rect 3532 2929 3533 3132
rect 3582 3131 3583 3154
rect 3678 2929 3679 3132
rect 3718 2929 3719 3132
rect 3681 2929 3682 3134
rect 3703 3133 3704 3154
rect 3700 2929 3701 3136
rect 3718 3135 3719 3154
rect 3694 2929 3695 3138
rect 3700 3137 3701 3154
rect 3706 3137 3707 3154
rect 3794 3137 3795 3154
rect 3709 2929 3710 3140
rect 3721 3139 3722 3154
rect 3738 2929 3739 3140
rect 3762 3139 3763 3154
rect 3712 2929 3713 3142
rect 3737 3141 3738 3154
rect 3741 2929 3742 3142
rect 3765 3141 3766 3154
rect 3715 2929 3716 3144
rect 3740 3143 3741 3154
rect 3697 2929 3698 3146
rect 3715 3145 3716 3154
rect 3675 2929 3676 3148
rect 3697 3147 3698 3154
rect 3772 2929 3773 3148
rect 3789 2929 3790 3148
rect 3743 3149 3744 3154
rect 3771 3149 3772 3154
rect 3788 3149 3789 3154
rect 3808 3149 3809 3154
rect 3797 3151 3798 3154
rect 3801 3151 3802 3154
rect 3824 3151 3825 3154
rect 3831 3151 3832 3154
rect 2906 3160 2907 3453
rect 3069 3160 3070 3453
rect 2909 3162 2910 3453
rect 3129 3158 3130 3163
rect 2913 3164 2914 3453
rect 3141 3158 3142 3165
rect 2916 3166 2917 3453
rect 3075 3166 3076 3453
rect 2933 3158 2934 3169
rect 2949 3158 2950 3169
rect 2935 3170 2936 3453
rect 3258 3170 3259 3453
rect 2945 3158 2946 3173
rect 3029 3158 3030 3173
rect 2944 3174 2945 3453
rect 3321 3158 3322 3175
rect 2951 3176 2952 3453
rect 3363 3158 3364 3177
rect 2958 3178 2959 3453
rect 3369 3158 3370 3179
rect 2961 3158 2962 3181
rect 3312 3158 3313 3181
rect 2968 3158 2969 3183
rect 2980 3182 2981 3453
rect 2968 3184 2969 3453
rect 3309 3158 3310 3185
rect 2977 3186 2978 3453
rect 3501 3186 3502 3453
rect 2984 3188 2985 3453
rect 3156 3188 3157 3453
rect 2987 3190 2988 3453
rect 3144 3158 3145 3191
rect 2993 3158 2994 3193
rect 3002 3192 3003 3453
rect 3014 3158 3015 3193
rect 3105 3158 3106 3193
rect 3014 3194 3015 3453
rect 3023 3158 3024 3195
rect 3020 3196 3021 3453
rect 3306 3196 3307 3453
rect 3023 3198 3024 3453
rect 3414 3198 3415 3453
rect 3030 3200 3031 3453
rect 3468 3158 3469 3201
rect 3033 3202 3034 3453
rect 3048 3158 3049 3203
rect 3042 3158 3043 3205
rect 3168 3204 3169 3453
rect 3045 3158 3046 3207
rect 3471 3158 3472 3207
rect 3051 3208 3052 3453
rect 3060 3158 3061 3209
rect 3057 3210 3058 3453
rect 3727 3158 3728 3211
rect 3063 3212 3064 3453
rect 3072 3158 3073 3213
rect 3078 3158 3079 3213
rect 3339 3212 3340 3453
rect 3084 3158 3085 3215
rect 3102 3214 3103 3453
rect 3087 3158 3088 3217
rect 3105 3216 3106 3453
rect 3093 3218 3094 3453
rect 3096 3158 3097 3219
rect 2911 3158 2912 3221
rect 3096 3220 3097 3453
rect 3099 3158 3100 3221
rect 3114 3220 3115 3453
rect 3108 3158 3109 3223
rect 3117 3158 3118 3223
rect 3111 3158 3112 3225
rect 3129 3224 3130 3453
rect 3123 3158 3124 3227
rect 3165 3226 3166 3453
rect 3123 3228 3124 3453
rect 3150 3228 3151 3453
rect 3138 3158 3139 3231
rect 3141 3230 3142 3453
rect 3174 3158 3175 3231
rect 3429 3230 3430 3453
rect 3162 3158 3163 3233
rect 3174 3232 3175 3453
rect 3066 3158 3067 3235
rect 3162 3234 3163 3453
rect 3198 3234 3199 3453
rect 3198 3158 3199 3235
rect 3201 3234 3202 3453
rect 3276 3234 3277 3453
rect 3207 3236 3208 3453
rect 3324 3158 3325 3237
rect 3213 3238 3214 3453
rect 3237 3158 3238 3239
rect 3147 3158 3148 3241
rect 3237 3240 3238 3453
rect 3222 3158 3223 3243
rect 3633 3242 3634 3453
rect 3243 3244 3244 3453
rect 3294 3158 3295 3245
rect 3255 3158 3256 3247
rect 3300 3246 3301 3453
rect 3264 3248 3265 3453
rect 3285 3158 3286 3249
rect 3267 3158 3268 3251
rect 3342 3250 3343 3453
rect 3270 3252 3271 3453
rect 3273 3158 3274 3253
rect 3273 3254 3274 3453
rect 3288 3158 3289 3255
rect 3282 3256 3283 3453
rect 3354 3158 3355 3257
rect 3288 3258 3289 3453
rect 3351 3158 3352 3259
rect 3294 3260 3295 3453
rect 3327 3158 3328 3261
rect 3297 3158 3298 3263
rect 3336 3262 3337 3453
rect 3303 3158 3304 3265
rect 3330 3264 3331 3453
rect 3312 3266 3313 3453
rect 3366 3158 3367 3267
rect 3279 3158 3280 3269
rect 3366 3268 3367 3453
rect 3318 3158 3319 3271
rect 3381 3270 3382 3453
rect 3120 3158 3121 3273
rect 3318 3272 3319 3453
rect 3120 3274 3121 3453
rect 3126 3158 3127 3275
rect 3324 3274 3325 3453
rect 3396 3158 3397 3275
rect 3252 3276 3253 3453
rect 3396 3276 3397 3453
rect 3348 3278 3349 3453
rect 3444 3158 3445 3279
rect 3354 3280 3355 3453
rect 3450 3158 3451 3281
rect 3360 3282 3361 3453
rect 3390 3158 3391 3283
rect 3372 3158 3373 3285
rect 3756 3284 3757 3453
rect 3372 3286 3373 3453
rect 3456 3158 3457 3287
rect 3375 3288 3376 3453
rect 3712 3158 3713 3289
rect 3378 3158 3379 3291
rect 3660 3158 3661 3291
rect 3315 3158 3316 3293
rect 3378 3292 3379 3453
rect 2961 3294 2962 3453
rect 3315 3294 3316 3453
rect 3390 3294 3391 3453
rect 3480 3158 3481 3295
rect 3393 3158 3394 3297
rect 3423 3296 3424 3453
rect 3402 3158 3403 3299
rect 3688 3158 3689 3299
rect 3402 3300 3403 3453
rect 3486 3158 3487 3301
rect 3408 3158 3409 3303
rect 3657 3158 3658 3303
rect 3333 3158 3334 3305
rect 3408 3304 3409 3453
rect 3426 3158 3427 3305
rect 3681 3158 3682 3305
rect 3027 3306 3028 3453
rect 3426 3306 3427 3453
rect 3435 3306 3436 3453
rect 3528 3158 3529 3307
rect 3441 3308 3442 3453
rect 3462 3158 3463 3309
rect 3459 3310 3460 3453
rect 3534 3158 3535 3311
rect 3240 3158 3241 3313
rect 3534 3312 3535 3453
rect 3240 3314 3241 3453
rect 3291 3158 3292 3315
rect 2921 3158 2922 3317
rect 3291 3316 3292 3453
rect 2920 3318 2921 3453
rect 3483 3158 3484 3319
rect 3471 3320 3472 3453
rect 3540 3158 3541 3321
rect 3477 3322 3478 3453
rect 3797 3158 3798 3323
rect 3483 3324 3484 3453
rect 3706 3158 3707 3325
rect 3489 3326 3490 3453
rect 3570 3158 3571 3327
rect 3492 3158 3493 3329
rect 3723 3328 3724 3453
rect 3504 3158 3505 3331
rect 3709 3158 3710 3331
rect 3246 3158 3247 3333
rect 3504 3332 3505 3453
rect 3210 3158 3211 3335
rect 3246 3334 3247 3453
rect 3210 3336 3211 3453
rect 3234 3158 3235 3337
rect 3234 3338 3235 3453
rect 3785 3158 3786 3339
rect 3507 3158 3508 3341
rect 3642 3340 3643 3453
rect 3507 3342 3508 3453
rect 3546 3158 3547 3343
rect 3513 3158 3514 3345
rect 3685 3158 3686 3345
rect 3216 3158 3217 3347
rect 3513 3346 3514 3453
rect 3516 3158 3517 3347
rect 3648 3346 3649 3453
rect 3522 3158 3523 3349
rect 3784 3348 3785 3453
rect 3525 3350 3526 3453
rect 3612 3158 3613 3351
rect 3420 3158 3421 3353
rect 3612 3352 3613 3453
rect 3228 3158 3229 3355
rect 3420 3354 3421 3453
rect 3228 3356 3229 3453
rect 3249 3158 3250 3357
rect 3540 3356 3541 3453
rect 3600 3158 3601 3357
rect 3552 3358 3553 3453
rect 3585 3158 3586 3359
rect 3564 3360 3565 3453
rect 3897 3360 3898 3453
rect 3570 3362 3571 3453
rect 3627 3158 3628 3363
rect 3573 3364 3574 3453
rect 3630 3158 3631 3365
rect 3465 3158 3466 3367
rect 3630 3366 3631 3453
rect 3465 3368 3466 3453
rect 3780 3368 3781 3453
rect 3576 3370 3577 3453
rect 3827 3370 3828 3453
rect 3582 3158 3583 3373
rect 3687 3372 3688 3453
rect 3582 3374 3583 3453
rect 3791 3158 3792 3375
rect 3594 3376 3595 3453
rect 3606 3158 3607 3377
rect 3621 3158 3622 3377
rect 3693 3376 3694 3453
rect 3645 3158 3646 3379
rect 3660 3378 3661 3453
rect 3438 3158 3439 3381
rect 3645 3380 3646 3453
rect 3666 3380 3667 3453
rect 3669 3158 3670 3381
rect 3669 3382 3670 3453
rect 3746 3158 3747 3383
rect 3192 3158 3193 3385
rect 3747 3384 3748 3453
rect 3186 3158 3187 3387
rect 3192 3386 3193 3453
rect 3180 3158 3181 3389
rect 3186 3388 3187 3453
rect 2964 3158 2965 3391
rect 3180 3390 3181 3453
rect 2965 3392 2966 3453
rect 3204 3392 3205 3453
rect 3681 3392 3682 3453
rect 3765 3158 3766 3393
rect 3690 3394 3691 3453
rect 3766 3394 3767 3453
rect 3697 3158 3698 3397
rect 3732 3396 3733 3453
rect 3624 3158 3625 3399
rect 3696 3398 3697 3453
rect 3543 3158 3544 3401
rect 3624 3400 3625 3453
rect 3700 3158 3701 3401
rect 3735 3400 3736 3453
rect 3495 3158 3496 3403
rect 3699 3402 3700 3453
rect 3261 3158 3262 3405
rect 3495 3404 3496 3453
rect 3705 3404 3706 3453
rect 3721 3158 3722 3405
rect 3715 3158 3716 3407
rect 3844 3406 3845 3453
rect 3678 3158 3679 3409
rect 3714 3408 3715 3453
rect 3737 3158 3738 3409
rect 3790 3408 3791 3453
rect 3703 3158 3704 3411
rect 3738 3410 3739 3453
rect 3195 3158 3196 3413
rect 3702 3412 3703 3453
rect 3743 3158 3744 3413
rect 3796 3412 3797 3453
rect 3357 3158 3358 3415
rect 3744 3414 3745 3453
rect 3357 3416 3358 3453
rect 3453 3158 3454 3417
rect 3384 3158 3385 3419
rect 3453 3418 3454 3453
rect 3384 3420 3385 3453
rect 3432 3158 3433 3421
rect 3432 3422 3433 3453
rect 3510 3158 3511 3423
rect 3750 3422 3751 3453
rect 3841 3422 3842 3453
rect 3752 3158 3753 3425
rect 3794 3158 3795 3425
rect 3718 3158 3719 3427
rect 3753 3426 3754 3453
rect 3717 3428 3718 3453
rect 3851 3428 3852 3453
rect 3740 3158 3741 3431
rect 3793 3430 3794 3453
rect 3741 3432 3742 3453
rect 3866 3432 3867 3453
rect 3762 3158 3763 3435
rect 3863 3434 3864 3453
rect 3768 3158 3769 3437
rect 3817 3436 3818 3453
rect 3788 3158 3789 3439
rect 3854 3438 3855 3453
rect 3588 3158 3589 3441
rect 3787 3440 3788 3453
rect 3804 3158 3805 3441
rect 3887 3440 3888 3453
rect 3811 3158 3812 3443
rect 3876 3442 3877 3453
rect 3815 3158 3816 3445
rect 3857 3444 3858 3453
rect 3771 3158 3772 3447
rect 3814 3446 3815 3453
rect 3831 3158 3832 3447
rect 3838 3158 3839 3447
rect 3558 3158 3559 3449
rect 3830 3448 3831 3453
rect 3558 3450 3559 3453
rect 3615 3158 3616 3451
rect 3860 3450 3861 3453
rect 3880 3450 3881 3453
rect 2815 3459 2816 3776
rect 2822 3459 2823 3776
rect 2878 3457 2879 3460
rect 3219 3459 3220 3776
rect 2884 3461 2885 3776
rect 3216 3461 3217 3776
rect 2899 3457 2900 3464
rect 3084 3463 3085 3776
rect 2908 3465 2909 3776
rect 3102 3457 3103 3466
rect 2913 3457 2914 3468
rect 3069 3457 3070 3468
rect 2916 3457 2917 3470
rect 3063 3457 3064 3470
rect 2915 3471 2916 3776
rect 3075 3457 3076 3472
rect 2918 3473 2919 3776
rect 3282 3457 3283 3474
rect 2920 3457 2921 3476
rect 3291 3457 3292 3476
rect 2935 3457 2936 3478
rect 3264 3457 3265 3478
rect 2939 3479 2940 3776
rect 3204 3457 3205 3480
rect 2942 3481 2943 3776
rect 3129 3457 3130 3482
rect 2949 3483 2950 3776
rect 2954 3457 2955 3484
rect 2958 3457 2959 3484
rect 2972 3483 2973 3776
rect 2961 3457 2962 3486
rect 3267 3485 3268 3776
rect 2965 3457 2966 3488
rect 3330 3457 3331 3488
rect 2968 3457 2969 3490
rect 3336 3457 3337 3490
rect 2978 3491 2979 3776
rect 3315 3457 3316 3492
rect 2980 3457 2981 3494
rect 3324 3457 3325 3494
rect 2987 3457 2988 3496
rect 3162 3457 3163 3496
rect 2990 3497 2991 3776
rect 3357 3457 3358 3498
rect 2993 3499 2994 3776
rect 3315 3499 3316 3776
rect 3008 3501 3009 3776
rect 3014 3457 3015 3502
rect 3014 3503 3015 3776
rect 3027 3457 3028 3504
rect 3033 3457 3034 3504
rect 3075 3503 3076 3776
rect 3039 3505 3040 3776
rect 3093 3457 3094 3506
rect 3042 3507 3043 3776
rect 3168 3457 3169 3508
rect 3048 3509 3049 3776
rect 3096 3457 3097 3510
rect 3051 3457 3052 3512
rect 3060 3511 3061 3776
rect 3051 3513 3052 3776
rect 3105 3457 3106 3514
rect 3054 3515 3055 3776
rect 3252 3457 3253 3516
rect 3057 3457 3058 3518
rect 3138 3517 3139 3776
rect 3066 3519 3067 3776
rect 3114 3457 3115 3520
rect 3072 3521 3073 3776
rect 3120 3457 3121 3522
rect 3081 3523 3082 3776
rect 3141 3457 3142 3524
rect 3087 3525 3088 3776
rect 3207 3457 3208 3526
rect 3114 3527 3115 3776
rect 3156 3457 3157 3528
rect 3120 3529 3121 3776
rect 3180 3457 3181 3530
rect 3036 3531 3037 3776
rect 3180 3531 3181 3776
rect 3126 3457 3127 3534
rect 3165 3457 3166 3534
rect 3126 3535 3127 3776
rect 3186 3457 3187 3536
rect 3132 3537 3133 3776
rect 3192 3457 3193 3538
rect 2960 3539 2961 3776
rect 3192 3539 3193 3776
rect 3144 3541 3145 3776
rect 3234 3457 3235 3542
rect 2947 3457 2948 3544
rect 3234 3543 3235 3776
rect 3147 3545 3148 3776
rect 3237 3457 3238 3546
rect 3156 3547 3157 3776
rect 3210 3457 3211 3548
rect 3159 3549 3160 3776
rect 3213 3457 3214 3550
rect 3168 3551 3169 3776
rect 3246 3457 3247 3552
rect 2891 3553 2892 3776
rect 3246 3553 3247 3776
rect 3186 3555 3187 3776
rect 3240 3457 3241 3556
rect 3189 3557 3190 3776
rect 3243 3457 3244 3558
rect 3198 3457 3199 3560
rect 3426 3457 3427 3560
rect 3198 3561 3199 3776
rect 3420 3457 3421 3562
rect 3020 3457 3021 3564
rect 3420 3563 3421 3776
rect 3201 3457 3202 3566
rect 3450 3565 3451 3776
rect 3204 3567 3205 3776
rect 3258 3457 3259 3568
rect 3222 3569 3223 3776
rect 3270 3457 3271 3570
rect 3225 3571 3226 3776
rect 3273 3457 3274 3572
rect 3240 3573 3241 3776
rect 3294 3457 3295 3574
rect 3249 3575 3250 3776
rect 3288 3457 3289 3576
rect 3252 3577 3253 3776
rect 3300 3457 3301 3578
rect 3255 3457 3256 3580
rect 3432 3457 3433 3580
rect 3258 3581 3259 3776
rect 3342 3457 3343 3582
rect 3264 3583 3265 3776
rect 3312 3457 3313 3584
rect 3270 3585 3271 3776
rect 3408 3457 3409 3586
rect 3276 3457 3277 3588
rect 3766 3457 3767 3588
rect 3276 3589 3277 3776
rect 3318 3457 3319 3590
rect 3023 3457 3024 3592
rect 3318 3591 3319 3776
rect 3279 3593 3280 3776
rect 3339 3457 3340 3594
rect 3282 3595 3283 3776
rect 3366 3457 3367 3596
rect 3174 3457 3175 3598
rect 3366 3597 3367 3776
rect 3174 3599 3175 3776
rect 3228 3457 3229 3600
rect 3228 3601 3229 3776
rect 3306 3457 3307 3602
rect 3288 3603 3289 3776
rect 3378 3457 3379 3604
rect 3291 3605 3292 3776
rect 3381 3457 3382 3606
rect 3294 3607 3295 3776
rect 3360 3457 3361 3608
rect 3300 3609 3301 3776
rect 3414 3457 3415 3610
rect 3306 3611 3307 3776
rect 3348 3457 3349 3612
rect 3312 3613 3313 3776
rect 3354 3457 3355 3614
rect 3321 3615 3322 3776
rect 3423 3457 3424 3616
rect 3324 3617 3325 3776
rect 3363 3617 3364 3776
rect 3330 3619 3331 3776
rect 3372 3457 3373 3620
rect 3348 3621 3349 3776
rect 3390 3457 3391 3622
rect 3354 3623 3355 3776
rect 3396 3457 3397 3624
rect 3369 3625 3370 3776
rect 3375 3457 3376 3626
rect 3378 3625 3379 3776
rect 3453 3457 3454 3626
rect 3384 3457 3385 3628
rect 3453 3627 3454 3776
rect 3150 3457 3151 3630
rect 3384 3629 3385 3776
rect 2956 3631 2957 3776
rect 3150 3631 3151 3776
rect 3390 3631 3391 3776
rect 3723 3457 3724 3632
rect 3396 3633 3397 3776
rect 3459 3457 3460 3634
rect 3402 3457 3403 3636
rect 3720 3457 3721 3636
rect 3408 3637 3409 3776
rect 3777 3457 3778 3638
rect 3414 3639 3415 3776
rect 3504 3457 3505 3640
rect 3417 3641 3418 3776
rect 3501 3457 3502 3642
rect 3426 3643 3427 3776
rect 3489 3457 3490 3644
rect 3429 3457 3430 3646
rect 3748 3645 3749 3776
rect 3432 3647 3433 3776
rect 3477 3457 3478 3648
rect 3435 3457 3436 3650
rect 3894 3457 3895 3650
rect 3444 3651 3445 3776
rect 3507 3457 3508 3652
rect 3456 3653 3457 3776
rect 3552 3457 3553 3654
rect 3465 3457 3466 3656
rect 3787 3457 3788 3656
rect 3468 3657 3469 3776
rect 3540 3457 3541 3658
rect 3471 3457 3472 3660
rect 3780 3457 3781 3660
rect 3474 3661 3475 3776
rect 3525 3457 3526 3662
rect 3483 3457 3484 3664
rect 3723 3663 3724 3776
rect 3489 3665 3490 3776
rect 3558 3457 3559 3666
rect 3045 3667 3046 3776
rect 3558 3667 3559 3776
rect 3495 3457 3496 3670
rect 3531 3669 3532 3776
rect 3501 3671 3502 3776
rect 3576 3457 3577 3672
rect 3507 3673 3508 3776
rect 3570 3457 3571 3674
rect 3510 3675 3511 3776
rect 3573 3457 3574 3676
rect 3513 3457 3514 3678
rect 3567 3677 3568 3776
rect 3513 3679 3514 3776
rect 3594 3457 3595 3680
rect 3441 3457 3442 3682
rect 3594 3681 3595 3776
rect 3519 3683 3520 3776
rect 3582 3457 3583 3684
rect 3525 3685 3526 3776
rect 3763 3457 3764 3686
rect 3534 3457 3535 3688
rect 3591 3687 3592 3776
rect 3537 3689 3538 3776
rect 3857 3457 3858 3690
rect 3543 3691 3544 3776
rect 3897 3457 3898 3692
rect 3549 3693 3550 3776
rect 3821 3693 3822 3776
rect 3561 3695 3562 3776
rect 3624 3457 3625 3696
rect 3573 3697 3574 3776
rect 3612 3457 3613 3698
rect 3579 3699 3580 3776
rect 3756 3457 3757 3700
rect 3585 3701 3586 3776
rect 3759 3457 3760 3702
rect 3597 3703 3598 3776
rect 3753 3457 3754 3704
rect 3600 3705 3601 3776
rect 3835 3705 3836 3776
rect 3615 3707 3616 3776
rect 3660 3457 3661 3708
rect 3621 3709 3622 3776
rect 3699 3457 3700 3710
rect 3387 3711 3388 3776
rect 3699 3711 3700 3776
rect 3624 3713 3625 3776
rect 3702 3457 3703 3714
rect 3627 3715 3628 3776
rect 3669 3457 3670 3716
rect 3630 3457 3631 3718
rect 3744 3457 3745 3718
rect 3645 3457 3646 3720
rect 3755 3719 3756 3776
rect 3645 3721 3646 3776
rect 3705 3457 3706 3722
rect 3651 3723 3652 3776
rect 3752 3723 3753 3776
rect 3666 3457 3667 3726
rect 3857 3725 3858 3776
rect 3648 3457 3649 3728
rect 3666 3727 3667 3776
rect 3642 3457 3643 3730
rect 3648 3729 3649 3776
rect 3672 3729 3673 3776
rect 3687 3457 3688 3730
rect 3675 3731 3676 3776
rect 3690 3457 3691 3732
rect 3684 3733 3685 3776
rect 3693 3457 3694 3734
rect 3687 3735 3688 3776
rect 3696 3457 3697 3736
rect 3633 3457 3634 3738
rect 3696 3737 3697 3776
rect 3633 3739 3634 3776
rect 3681 3457 3682 3740
rect 3702 3739 3703 3776
rect 3714 3457 3715 3740
rect 3705 3741 3706 3776
rect 3717 3457 3718 3742
rect 3720 3741 3721 3776
rect 3738 3457 3739 3742
rect 3654 3743 3655 3776
rect 3738 3743 3739 3776
rect 3726 3745 3727 3776
rect 3732 3457 3733 3746
rect 3741 3457 3742 3746
rect 3842 3745 3843 3776
rect 3660 3747 3661 3776
rect 3741 3747 3742 3776
rect 3750 3457 3751 3748
rect 3873 3457 3874 3748
rect 3770 3457 3771 3750
rect 3851 3749 3852 3776
rect 3778 3751 3779 3776
rect 3831 3751 3832 3776
rect 3784 3753 3785 3776
rect 3790 3457 3791 3754
rect 3787 3755 3788 3776
rect 3793 3457 3794 3756
rect 3790 3757 3791 3776
rect 3796 3457 3797 3758
rect 3796 3759 3797 3776
rect 3863 3457 3864 3760
rect 3799 3761 3800 3776
rect 3868 3761 3869 3776
rect 3808 3763 3809 3776
rect 3814 3457 3815 3764
rect 3735 3457 3736 3766
rect 3814 3765 3815 3776
rect 3811 3767 3812 3776
rect 3817 3457 3818 3768
rect 3729 3769 3730 3776
rect 3817 3769 3818 3776
rect 3838 3769 3839 3776
rect 3848 3457 3849 3770
rect 3848 3771 3849 3776
rect 3854 3457 3855 3772
rect 3860 3457 3861 3772
rect 3887 3457 3888 3772
rect 3564 3457 3565 3774
rect 3861 3773 3862 3776
rect 2881 3780 2882 3783
rect 3219 3780 3220 3783
rect 2893 3784 2894 4069
rect 3246 3780 3247 3785
rect 2900 3786 2901 4069
rect 2901 3780 2902 3787
rect 2904 3780 2905 3787
rect 3361 3786 3362 4069
rect 2908 3780 2909 3789
rect 3430 3788 3431 4069
rect 2915 3780 2916 3791
rect 2926 3790 2927 4069
rect 2942 3780 2943 3791
rect 3238 3790 3239 4069
rect 2946 3780 2947 3793
rect 2957 3792 2958 4069
rect 2949 3780 2950 3795
rect 3346 3794 3347 4069
rect 2960 3780 2961 3797
rect 3198 3780 3199 3797
rect 2963 3780 2964 3799
rect 3008 3780 3009 3799
rect 2918 3780 2919 3801
rect 3008 3800 3009 4069
rect 2953 3780 2954 3803
rect 2964 3802 2965 4069
rect 2953 3804 2954 4069
rect 3189 3780 3190 3805
rect 2967 3806 2968 4069
rect 3412 3806 3413 4069
rect 2972 3780 2973 3809
rect 2990 3808 2991 4069
rect 2971 3810 2972 4069
rect 3279 3780 3280 3811
rect 2884 3780 2885 3813
rect 3280 3812 3281 4069
rect 2978 3780 2979 3815
rect 2996 3814 2997 4069
rect 2978 3816 2979 4069
rect 3163 3816 3164 4069
rect 2981 3818 2982 4069
rect 3132 3780 3133 3819
rect 3014 3820 3015 4069
rect 3382 3820 3383 4069
rect 3017 3780 3018 3823
rect 3436 3822 3437 4069
rect 2950 3824 2951 4069
rect 3017 3824 3018 4069
rect 3036 3780 3037 3825
rect 3321 3780 3322 3825
rect 3039 3780 3040 3827
rect 3130 3826 3131 4069
rect 3038 3828 3039 4069
rect 3315 3780 3316 3829
rect 3042 3780 3043 3831
rect 3472 3830 3473 4069
rect 3045 3780 3046 3833
rect 3324 3780 3325 3833
rect 3048 3780 3049 3835
rect 3058 3834 3059 4069
rect 3048 3836 3049 4069
rect 3310 3836 3311 4069
rect 3060 3780 3061 3839
rect 3064 3838 3065 4069
rect 3066 3780 3067 3839
rect 3070 3838 3071 4069
rect 3081 3780 3082 3839
rect 3106 3838 3107 4069
rect 3084 3780 3085 3841
rect 3364 3840 3365 4069
rect 3112 3842 3113 4069
rect 3138 3780 3139 3843
rect 3114 3780 3115 3845
rect 3118 3844 3119 4069
rect 3120 3780 3121 3845
rect 3190 3844 3191 4069
rect 3124 3846 3125 4069
rect 3648 3780 3649 3847
rect 3126 3780 3127 3849
rect 3487 3848 3488 4069
rect 3139 3850 3140 4069
rect 3366 3780 3367 3851
rect 3144 3780 3145 3853
rect 3232 3852 3233 4069
rect 3156 3780 3157 3855
rect 3274 3854 3275 4069
rect 2922 3856 2923 4069
rect 3157 3856 3158 4069
rect 3168 3780 3169 3857
rect 3244 3856 3245 4069
rect 3174 3780 3175 3859
rect 3298 3858 3299 4069
rect 3072 3780 3073 3861
rect 3175 3860 3176 4069
rect 3180 3780 3181 3861
rect 3184 3860 3185 4069
rect 3186 3780 3187 3861
rect 3328 3860 3329 4069
rect 3204 3780 3205 3863
rect 3334 3862 3335 4069
rect 3208 3864 3209 4069
rect 3567 3780 3568 3865
rect 3222 3780 3223 3867
rect 3316 3866 3317 4069
rect 3223 3868 3224 4069
rect 3624 3780 3625 3869
rect 3225 3780 3226 3871
rect 3337 3870 3338 4069
rect 3150 3780 3151 3873
rect 3226 3872 3227 4069
rect 3228 3780 3229 3873
rect 3262 3872 3263 4069
rect 3234 3780 3235 3875
rect 3304 3874 3305 4069
rect 3240 3780 3241 3877
rect 3367 3876 3368 4069
rect 3087 3780 3088 3879
rect 3241 3878 3242 4069
rect 3075 3780 3076 3881
rect 3088 3880 3089 4069
rect 3054 3780 3055 3883
rect 3076 3882 3077 4069
rect 3055 3884 3056 4069
rect 3439 3884 3440 4069
rect 3256 3886 3257 4069
rect 3480 3780 3481 3887
rect 3258 3780 3259 3889
rect 3340 3888 3341 4069
rect 3264 3780 3265 3891
rect 3394 3890 3395 4069
rect 3276 3780 3277 3893
rect 3406 3892 3407 4069
rect 3282 3780 3283 3895
rect 3373 3894 3374 4069
rect 3159 3780 3160 3897
rect 3283 3896 3284 4069
rect 3286 3896 3287 4069
rect 3300 3780 3301 3897
rect 3288 3780 3289 3899
rect 3755 3898 3756 4069
rect 3291 3780 3292 3901
rect 3376 3900 3377 4069
rect 3252 3780 3253 3903
rect 3292 3902 3293 4069
rect 3294 3780 3295 3903
rect 3442 3902 3443 4069
rect 3306 3780 3307 3905
rect 3478 3904 3479 4069
rect 3312 3780 3313 3907
rect 3484 3906 3485 4069
rect 3318 3780 3319 3909
rect 3322 3908 3323 4069
rect 3369 3780 3370 3909
rect 3505 3908 3506 4069
rect 3378 3780 3379 3911
rect 3448 3910 3449 4069
rect 3249 3780 3250 3913
rect 3379 3912 3380 4069
rect 3250 3914 3251 4069
rect 3531 3780 3532 3915
rect 3384 3780 3385 3917
rect 3403 3916 3404 4069
rect 3387 3780 3388 3919
rect 3400 3918 3401 4069
rect 3390 3780 3391 3921
rect 3553 3920 3554 4069
rect 3396 3780 3397 3923
rect 3547 3922 3548 4069
rect 3408 3780 3409 3925
rect 3762 3780 3763 3925
rect 2939 3780 2940 3927
rect 3409 3926 3410 4069
rect 2929 3928 2930 4069
rect 2938 3928 2939 4069
rect 3417 3780 3418 3929
rect 3424 3928 3425 4069
rect 3418 3930 3419 4069
rect 3585 3780 3586 3931
rect 3420 3780 3421 3933
rect 3466 3932 3467 4069
rect 3444 3780 3445 3935
rect 3571 3934 3572 4069
rect 3033 3780 3034 3937
rect 3445 3936 3446 4069
rect 3032 3938 3033 4069
rect 3147 3780 3148 3939
rect 3450 3780 3451 3939
rect 3523 3938 3524 4069
rect 3456 3780 3457 3941
rect 3589 3940 3590 4069
rect 3468 3780 3469 3943
rect 3613 3942 3614 4069
rect 3469 3944 3470 4069
rect 3621 3780 3622 3945
rect 3474 3780 3475 3947
rect 3943 3946 3944 4069
rect 3489 3780 3490 3949
rect 3637 3948 3638 4069
rect 3453 3780 3454 3951
rect 3490 3950 3491 4069
rect 3454 3952 3455 4069
rect 3708 3780 3709 3953
rect 3496 3954 3497 4069
rect 3654 3780 3655 3955
rect 3501 3780 3502 3957
rect 3619 3956 3620 4069
rect 3330 3780 3331 3959
rect 3502 3958 3503 4069
rect 2897 3780 2898 3961
rect 3331 3960 3332 4069
rect 2896 3962 2897 4069
rect 3216 3780 3217 3963
rect 3507 3780 3508 3963
rect 3649 3962 3650 4069
rect 3354 3780 3355 3965
rect 3508 3964 3509 4069
rect 3510 3780 3511 3965
rect 3896 3964 3897 4069
rect 3414 3780 3415 3967
rect 3511 3966 3512 4069
rect 3267 3780 3268 3969
rect 3415 3968 3416 4069
rect 3192 3780 3193 3971
rect 3268 3970 3269 4069
rect 3513 3780 3514 3971
rect 3655 3970 3656 4069
rect 3525 3780 3526 3973
rect 3882 3972 3883 4069
rect 3526 3974 3527 4069
rect 3731 3974 3732 4069
rect 3529 3976 3530 4069
rect 3594 3780 3595 3977
rect 3532 3978 3533 4069
rect 3660 3780 3661 3979
rect 3519 3780 3520 3981
rect 3661 3980 3662 4069
rect 3348 3780 3349 3983
rect 3520 3982 3521 4069
rect 3270 3780 3271 3985
rect 3349 3984 3350 4069
rect 3537 3780 3538 3985
rect 3915 3984 3916 4069
rect 3538 3986 3539 4069
rect 3734 3986 3735 4069
rect 3541 3988 3542 4069
rect 3558 3780 3559 3989
rect 3543 3780 3544 3991
rect 3918 3990 3919 4069
rect 3549 3780 3550 3993
rect 3770 3992 3771 4069
rect 3555 3780 3556 3995
rect 3591 3780 3592 3995
rect 3559 3996 3560 4069
rect 3842 3780 3843 3997
rect 3561 3780 3562 3999
rect 3631 3998 3632 4069
rect 3573 3780 3574 4001
rect 3577 4000 3578 4069
rect 3579 3780 3580 4001
rect 3711 3780 3712 4001
rect 3580 4002 3581 4069
rect 3752 3780 3753 4003
rect 3597 3780 3598 4005
rect 3764 4004 3765 4069
rect 3600 3780 3601 4007
rect 3625 4006 3626 4069
rect 3432 3780 3433 4009
rect 3601 4008 3602 4069
rect 3051 3780 3052 4011
rect 3433 4010 3434 4069
rect 3607 4010 3608 4069
rect 3675 3780 3676 4011
rect 3627 3780 3628 4013
rect 3868 4012 3869 4069
rect 3633 3780 3634 4015
rect 3743 4014 3744 4069
rect 3643 4016 3644 4069
rect 3861 3780 3862 4017
rect 3645 3780 3646 4019
rect 3773 4018 3774 4069
rect 3651 3780 3652 4021
rect 3821 3780 3822 4021
rect 3426 3780 3427 4023
rect 3652 4022 3653 4069
rect 3666 3780 3667 4023
rect 3741 3780 3742 4023
rect 3667 4024 3668 4069
rect 3946 4024 3947 4069
rect 3670 4026 3671 4069
rect 3885 4026 3886 4069
rect 3684 3780 3685 4029
rect 3691 4028 3692 4069
rect 3687 3780 3688 4031
rect 3688 4030 3689 4069
rect 3694 4030 3695 4069
rect 3857 3780 3858 4031
rect 3705 3780 3706 4033
rect 3752 4032 3753 4069
rect 3615 3780 3616 4035
rect 3706 4034 3707 4069
rect 3720 3780 3721 4035
rect 3776 4034 3777 4069
rect 3721 4036 3722 4069
rect 3766 3780 3767 4037
rect 3726 3780 3727 4039
rect 3817 3780 3818 4039
rect 3696 3780 3697 4041
rect 3727 4040 3728 4069
rect 3729 3780 3730 4041
rect 3767 4040 3768 4069
rect 3737 4042 3738 4069
rect 3787 3780 3788 4043
rect 3748 3780 3749 4045
rect 3759 3780 3760 4045
rect 3460 4046 3461 4069
rect 3758 4046 3759 4069
rect 3702 3780 3703 4049
rect 3749 4048 3750 4069
rect 3761 4048 3762 4069
rect 3889 4048 3890 4069
rect 3778 3780 3779 4051
rect 3814 4050 3815 4069
rect 3723 3780 3724 4053
rect 3779 4052 3780 4069
rect 3784 3780 3785 4053
rect 3862 4052 3863 4069
rect 3790 3780 3791 4055
rect 3838 4054 3839 4069
rect 3796 3780 3797 4057
rect 3844 4056 3845 4069
rect 3808 3780 3809 4059
rect 3856 4058 3857 4069
rect 3718 4060 3719 4069
rect 3808 4060 3809 4069
rect 3811 3780 3812 4061
rect 3859 4060 3860 4069
rect 3672 3780 3673 4063
rect 3811 4062 3812 4069
rect 3820 4062 3821 4069
rect 3831 3780 3832 4063
rect 3848 3780 3849 4063
rect 3902 4062 3903 4069
rect 3799 3780 3800 4065
rect 3847 4064 3848 4069
rect 3851 3780 3852 4065
rect 3905 4064 3906 4069
rect 3865 4066 3866 4069
rect 3878 4066 3879 4069
rect 3925 4066 3926 4069
rect 3929 4066 3930 4069
rect 2809 4075 2810 4346
rect 3175 4073 3176 4076
rect 2887 4077 2888 4346
rect 3280 4073 3281 4078
rect 2907 4073 2908 4080
rect 3058 4073 3059 4080
rect 2918 4081 2919 4346
rect 3433 4073 3434 4082
rect 2922 4073 2923 4084
rect 3430 4073 3431 4084
rect 2926 4073 2927 4086
rect 3457 4085 3458 4346
rect 2925 4087 2926 4346
rect 3394 4073 3395 4088
rect 2928 4089 2929 4346
rect 3391 4089 3392 4346
rect 2935 4091 2936 4346
rect 3316 4073 3317 4092
rect 2941 4073 2942 4094
rect 3298 4073 3299 4094
rect 2944 4095 2945 4346
rect 3385 4095 3386 4346
rect 2947 4097 2948 4346
rect 3286 4073 3287 4098
rect 2954 4099 2955 4346
rect 3346 4073 3347 4100
rect 2961 4101 2962 4346
rect 3190 4073 3191 4102
rect 2971 4073 2972 4104
rect 3430 4103 3431 4346
rect 2981 4073 2982 4106
rect 3487 4073 3488 4106
rect 2984 4107 2985 4346
rect 2990 4073 2991 4108
rect 2996 4073 2997 4108
rect 3739 4107 3740 4346
rect 2996 4109 2997 4346
rect 3172 4073 3173 4110
rect 3008 4109 3009 4346
rect 3008 4073 3009 4110
rect 3026 4111 3027 4346
rect 3032 4073 3033 4112
rect 3038 4073 3039 4112
rect 3472 4073 3473 4112
rect 3041 4073 3042 4114
rect 3436 4073 3437 4114
rect 3042 4115 3043 4346
rect 3382 4073 3383 4116
rect 3045 4073 3046 4118
rect 3064 4073 3065 4118
rect 2899 4119 2900 4346
rect 3045 4119 3046 4346
rect 3048 4073 3049 4120
rect 3292 4073 3293 4120
rect 2896 4073 2897 4122
rect 3292 4121 3293 4346
rect 3052 4073 3053 4124
rect 3403 4073 3404 4124
rect 2903 4073 2904 4126
rect 3051 4125 3052 4346
rect 3057 4125 3058 4346
rect 3310 4073 3311 4126
rect 3076 4073 3077 4128
rect 3081 4127 3082 4346
rect 3070 4073 3071 4130
rect 3075 4129 3076 4346
rect 3088 4073 3089 4130
rect 3093 4129 3094 4346
rect 3105 4129 3106 4346
rect 3106 4073 3107 4130
rect 3112 4073 3113 4130
rect 3132 4129 3133 4346
rect 3111 4131 3112 4346
rect 3147 4131 3148 4346
rect 3117 4133 3118 4346
rect 3118 4073 3119 4134
rect 3124 4073 3125 4134
rect 3517 4133 3518 4346
rect 3129 4135 3130 4346
rect 3130 4073 3131 4136
rect 3138 4135 3139 4346
rect 3139 4073 3140 4136
rect 3151 4135 3152 4346
rect 3487 4135 3488 4346
rect 3154 4137 3155 4346
rect 3286 4137 3287 4346
rect 3157 4137 3158 4346
rect 3157 4073 3158 4138
rect 3160 4139 3161 4346
rect 3163 4073 3164 4140
rect 3178 4139 3179 4346
rect 3184 4073 3185 4140
rect 2958 4141 2959 4346
rect 3184 4141 3185 4346
rect 3190 4141 3191 4346
rect 3523 4073 3524 4142
rect 3196 4143 3197 4346
rect 3211 4143 3212 4346
rect 3202 4145 3203 4346
rect 3409 4073 3410 4146
rect 3214 4147 3215 4346
rect 3232 4073 3233 4148
rect 3220 4149 3221 4346
rect 3226 4073 3227 4150
rect 3014 4073 3015 4152
rect 3226 4151 3227 4346
rect 3229 4151 3230 4346
rect 3439 4073 3440 4152
rect 3232 4153 3233 4346
rect 3238 4073 3239 4154
rect 3238 4155 3239 4346
rect 3244 4073 3245 4156
rect 3208 4073 3209 4158
rect 3244 4157 3245 4346
rect 3208 4159 3209 4346
rect 3424 4073 3425 4160
rect 3250 4073 3251 4162
rect 3727 4073 3728 4162
rect 3256 4073 3257 4164
rect 3316 4163 3317 4346
rect 3256 4165 3257 4346
rect 3262 4073 3263 4166
rect 3262 4167 3263 4346
rect 3274 4073 3275 4168
rect 3265 4169 3266 4346
rect 3283 4073 3284 4170
rect 3268 4073 3269 4172
rect 3274 4171 3275 4346
rect 2950 4073 2951 4174
rect 3268 4173 3269 4346
rect 3280 4173 3281 4346
rect 3322 4073 3323 4174
rect 3298 4175 3299 4346
rect 3304 4073 3305 4176
rect 2910 4073 2911 4178
rect 3304 4177 3305 4346
rect 3310 4177 3311 4346
rect 3334 4073 3335 4178
rect 3223 4073 3224 4180
rect 3334 4179 3335 4346
rect 3322 4181 3323 4346
rect 3328 4073 3329 4182
rect 2951 4183 2952 4346
rect 3328 4183 3329 4346
rect 3325 4185 3326 4346
rect 3331 4073 3332 4186
rect 3337 4073 3338 4186
rect 3352 4185 3353 4346
rect 2906 4187 2907 4346
rect 3337 4187 3338 4346
rect 3340 4073 3341 4188
rect 3343 4187 3344 4346
rect 3355 4187 3356 4346
rect 3367 4073 3368 4188
rect 3349 4073 3350 4190
rect 3367 4189 3368 4346
rect 2938 4073 2939 4192
rect 3349 4191 3350 4346
rect 3361 4191 3362 4346
rect 3361 4073 3362 4192
rect 3364 4191 3365 4346
rect 3364 4073 3365 4192
rect 3373 4073 3374 4192
rect 3397 4191 3398 4346
rect 3379 4073 3380 4194
rect 3394 4193 3395 4346
rect 3403 4193 3404 4346
rect 3496 4073 3497 4194
rect 3406 4073 3407 4196
rect 3427 4195 3428 4346
rect 3412 4073 3413 4198
rect 3421 4197 3422 4346
rect 3415 4073 3416 4200
rect 3424 4199 3425 4346
rect 3169 4073 3170 4202
rect 3415 4201 3416 4346
rect 3433 4201 3434 4346
rect 3466 4073 3467 4202
rect 3439 4203 3440 4346
rect 3442 4073 3443 4204
rect 3442 4205 3443 4346
rect 3445 4073 3446 4206
rect 3448 4073 3449 4206
rect 3734 4073 3735 4206
rect 3451 4207 3452 4346
rect 3460 4073 3461 4208
rect 3241 4073 3242 4210
rect 3460 4209 3461 4346
rect 3454 4073 3455 4212
rect 3463 4211 3464 4346
rect 3466 4211 3467 4346
rect 3469 4073 3470 4212
rect 3475 4211 3476 4346
rect 3526 4073 3527 4212
rect 3478 4073 3479 4214
rect 3493 4213 3494 4346
rect 3481 4215 3482 4346
rect 3490 4073 3491 4216
rect 3484 4073 3485 4218
rect 3499 4217 3500 4346
rect 3505 4073 3506 4218
rect 3526 4217 3527 4346
rect 3505 4219 3506 4346
rect 3529 4073 3530 4220
rect 3508 4073 3509 4222
rect 3529 4221 3530 4346
rect 3508 4223 3509 4346
rect 3797 4223 3798 4346
rect 3520 4073 3521 4226
rect 3535 4225 3536 4346
rect 3400 4073 3401 4228
rect 3520 4227 3521 4346
rect 3376 4073 3377 4230
rect 3400 4229 3401 4346
rect 3532 4073 3533 4230
rect 3709 4229 3710 4346
rect 3511 4073 3512 4232
rect 3532 4231 3533 4346
rect 3502 4073 3503 4234
rect 3511 4233 3512 4346
rect 2975 4235 2976 4346
rect 3502 4235 3503 4346
rect 3538 4073 3539 4236
rect 3782 4073 3783 4236
rect 3032 4237 3033 4346
rect 3538 4237 3539 4346
rect 3541 4073 3542 4238
rect 3562 4237 3563 4346
rect 3547 4073 3548 4240
rect 3568 4239 3569 4346
rect 3547 4241 3548 4346
rect 3801 4073 3802 4242
rect 3418 4073 3419 4244
rect 3800 4243 3801 4346
rect 3553 4073 3554 4246
rect 3574 4245 3575 4346
rect 3553 4247 3554 4346
rect 3577 4073 3578 4248
rect 3571 4073 3572 4250
rect 3586 4249 3587 4346
rect 3577 4251 3578 4346
rect 3580 4073 3581 4252
rect 3559 4073 3560 4254
rect 3580 4253 3581 4346
rect 3559 4255 3560 4346
rect 3816 4255 3817 4346
rect 3589 4073 3590 4258
rect 3598 4257 3599 4346
rect 3601 4073 3602 4258
rect 3616 4257 3617 4346
rect 3604 4259 3605 4346
rect 3652 4073 3653 4260
rect 3607 4073 3608 4262
rect 3610 4261 3611 4346
rect 3613 4073 3614 4262
rect 3628 4261 3629 4346
rect 3619 4073 3620 4264
rect 3622 4263 3623 4346
rect 3625 4073 3626 4264
rect 3634 4263 3635 4346
rect 3631 4073 3632 4266
rect 3755 4073 3756 4266
rect 3637 4073 3638 4268
rect 3652 4267 3653 4346
rect 3643 4073 3644 4270
rect 3658 4269 3659 4346
rect 3646 4271 3647 4346
rect 3649 4073 3650 4272
rect 3655 4073 3656 4272
rect 3664 4271 3665 4346
rect 3667 4073 3668 4272
rect 3685 4271 3686 4346
rect 3682 4273 3683 4346
rect 3941 4273 3942 4346
rect 3694 4073 3695 4276
rect 3712 4275 3713 4346
rect 3694 4277 3695 4346
rect 3871 4073 3872 4278
rect 3706 4073 3707 4280
rect 3724 4279 3725 4346
rect 3691 4073 3692 4282
rect 3706 4281 3707 4346
rect 3718 4281 3719 4346
rect 3718 4073 3719 4282
rect 3721 4073 3722 4282
rect 3808 4073 3809 4282
rect 3721 4283 3722 4346
rect 3915 4073 3916 4284
rect 3731 4073 3732 4286
rect 3826 4285 3827 4346
rect 3743 4073 3744 4288
rect 3922 4073 3923 4288
rect 3749 4073 3750 4290
rect 3758 4289 3759 4346
rect 3749 4291 3750 4346
rect 3951 4291 3952 4346
rect 3767 4073 3768 4294
rect 3788 4293 3789 4346
rect 3773 4073 3774 4296
rect 3794 4295 3795 4346
rect 3776 4073 3777 4298
rect 3874 4297 3875 4346
rect 3761 4073 3762 4300
rect 3776 4299 3777 4346
rect 3752 4073 3753 4302
rect 3761 4301 3762 4346
rect 3779 4073 3780 4302
rect 3908 4073 3909 4302
rect 3764 4073 3765 4304
rect 3779 4303 3780 4346
rect 3782 4303 3783 4346
rect 3927 4303 3928 4346
rect 3785 4073 3786 4306
rect 3792 4073 3793 4306
rect 3770 4073 3771 4308
rect 3791 4307 3792 4346
rect 3688 4073 3689 4310
rect 3770 4309 3771 4346
rect 3661 4073 3662 4312
rect 3688 4311 3689 4346
rect 3785 4311 3786 4346
rect 3931 4311 3932 4346
rect 3814 4073 3815 4314
rect 3889 4073 3890 4314
rect 3670 4073 3671 4316
rect 3888 4315 3889 4346
rect 3670 4317 3671 4346
rect 3899 4073 3900 4318
rect 3820 4073 3821 4320
rect 3835 4319 3836 4346
rect 3523 4321 3524 4346
rect 3819 4321 3820 4346
rect 3838 4073 3839 4322
rect 3871 4321 3872 4346
rect 3844 4073 3845 4324
rect 3868 4073 3869 4324
rect 3847 4073 3848 4326
rect 3850 4325 3851 4346
rect 3847 4327 3848 4346
rect 3918 4073 3919 4328
rect 3853 4329 3854 4346
rect 3865 4073 3866 4330
rect 3856 4073 3857 4332
rect 3865 4331 3866 4346
rect 3737 4073 3738 4334
rect 3856 4333 3857 4346
rect 3859 4073 3860 4334
rect 3868 4333 3869 4346
rect 3862 4073 3863 4336
rect 3878 4073 3879 4336
rect 3882 4073 3883 4336
rect 3924 4335 3925 4346
rect 3885 4335 3886 4346
rect 3885 4073 3886 4336
rect 3898 4337 3899 4346
rect 3936 4073 3937 4338
rect 3905 4073 3906 4340
rect 3907 4339 3908 4346
rect 3902 4073 3903 4342
rect 3904 4341 3905 4346
rect 3901 4343 3902 4346
rect 3917 4343 3918 4346
rect 2882 4352 2883 4659
rect 2991 4352 2992 4659
rect 2890 4350 2891 4355
rect 3262 4350 3263 4355
rect 2896 4356 2897 4659
rect 3322 4350 3323 4357
rect 2899 4350 2900 4359
rect 2921 4350 2922 4359
rect 2906 4360 2907 4659
rect 3364 4350 3365 4361
rect 2909 4350 2910 4363
rect 3340 4362 3341 4659
rect 2925 4350 2926 4365
rect 2972 4350 2973 4365
rect 2924 4366 2925 4659
rect 3406 4366 3407 4659
rect 2928 4350 2929 4369
rect 3385 4350 3386 4369
rect 2932 4350 2933 4371
rect 3292 4350 3293 4371
rect 2933 4372 2934 4659
rect 3310 4350 3311 4373
rect 2947 4350 2948 4375
rect 3349 4350 3350 4375
rect 2954 4376 2955 4659
rect 3238 4350 3239 4377
rect 2957 4378 2958 4659
rect 3427 4350 3428 4379
rect 2961 4350 2962 4381
rect 3331 4380 3332 4659
rect 2961 4382 2962 4659
rect 3493 4350 3494 4383
rect 2964 4384 2965 4659
rect 3181 4384 3182 4659
rect 2973 4386 2974 4659
rect 2984 4350 2985 4387
rect 2975 4350 2976 4389
rect 3211 4350 3212 4389
rect 2979 4390 2980 4659
rect 2996 4350 2997 4391
rect 2994 4392 2995 4659
rect 3265 4350 3266 4393
rect 2876 4394 2877 4659
rect 3265 4394 3266 4659
rect 2997 4396 2998 4659
rect 3008 4350 3009 4397
rect 2872 4398 2873 4659
rect 3009 4398 3010 4659
rect 3003 4400 3004 4659
rect 3226 4350 3227 4401
rect 3017 4350 3018 4403
rect 3502 4350 3503 4403
rect 3018 4404 3019 4659
rect 3026 4350 3027 4405
rect 3024 4406 3025 4659
rect 3256 4350 3257 4407
rect 3032 4350 3033 4409
rect 3421 4350 3422 4409
rect 3035 4350 3036 4411
rect 3583 4410 3584 4659
rect 2943 4412 2944 4659
rect 3036 4412 3037 4659
rect 3045 4350 3046 4413
rect 3048 4412 3049 4659
rect 3051 4350 3052 4413
rect 3054 4412 3055 4659
rect 3057 4350 3058 4413
rect 3502 4412 3503 4659
rect 3057 4414 3058 4659
rect 3325 4350 3326 4415
rect 3075 4350 3076 4417
rect 3078 4416 3079 4659
rect 3090 4416 3091 4659
rect 3093 4350 3094 4417
rect 3096 4416 3097 4659
rect 3111 4350 3112 4417
rect 3105 4350 3106 4419
rect 3108 4418 3109 4659
rect 3117 4350 3118 4419
rect 3120 4418 3121 4659
rect 3126 4418 3127 4659
rect 3132 4350 3133 4419
rect 3132 4420 3133 4659
rect 3160 4350 3161 4421
rect 3135 4422 3136 4659
rect 3814 4422 3815 4659
rect 3138 4350 3139 4425
rect 3934 4350 3935 4425
rect 3139 4426 3140 4659
rect 3196 4350 3197 4427
rect 2892 4428 2893 4659
rect 3196 4428 3197 4659
rect 3142 4430 3143 4659
rect 3199 4430 3200 4659
rect 3144 4350 3145 4433
rect 3217 4432 3218 4659
rect 3129 4350 3130 4435
rect 3145 4434 3146 4659
rect 3151 4350 3152 4435
rect 3816 4350 3817 4435
rect 3154 4350 3155 4437
rect 3481 4350 3482 4437
rect 3166 4438 3167 4659
rect 3190 4350 3191 4439
rect 3178 4350 3179 4441
rect 3190 4440 3191 4659
rect 3157 4350 3158 4443
rect 3178 4442 3179 4659
rect 3157 4444 3158 4659
rect 3310 4444 3311 4659
rect 3184 4350 3185 4447
rect 3205 4446 3206 4659
rect 3214 4350 3215 4447
rect 3253 4446 3254 4659
rect 3220 4350 3221 4449
rect 3235 4448 3236 4659
rect 3223 4450 3224 4659
rect 3244 4350 3245 4451
rect 3229 4350 3230 4453
rect 3409 4452 3410 4659
rect 3202 4350 3203 4455
rect 3229 4454 3230 4659
rect 3232 4350 3233 4455
rect 3241 4454 3242 4659
rect 3247 4454 3248 4659
rect 3316 4350 3317 4455
rect 3262 4456 3263 4659
rect 3334 4350 3335 4457
rect 3274 4350 3275 4459
rect 3292 4458 3293 4659
rect 3274 4460 3275 4659
rect 3280 4350 3281 4461
rect 3268 4350 3269 4463
rect 3280 4462 3281 4659
rect 3147 4350 3148 4465
rect 3268 4464 3269 4659
rect 3286 4464 3287 4659
rect 3286 4350 3287 4465
rect 3295 4464 3296 4659
rect 3430 4350 3431 4465
rect 3304 4350 3305 4467
rect 3316 4466 3317 4659
rect 3298 4350 3299 4469
rect 3304 4468 3305 4659
rect 3322 4468 3323 4659
rect 3403 4350 3404 4469
rect 3328 4468 3329 4659
rect 3328 4350 3329 4469
rect 3334 4470 3335 4659
rect 3343 4350 3344 4471
rect 3337 4350 3338 4473
rect 3346 4472 3347 4659
rect 3355 4350 3356 4473
rect 3370 4472 3371 4659
rect 3358 4474 3359 4659
rect 3361 4350 3362 4475
rect 3081 4350 3082 4477
rect 3361 4476 3362 4659
rect 3081 4478 3082 4659
rect 3352 4350 3353 4479
rect 3352 4480 3353 4659
rect 3367 4350 3368 4481
rect 3364 4482 3365 4659
rect 3433 4350 3434 4483
rect 3367 4484 3368 4659
rect 3466 4350 3467 4485
rect 2947 4486 2948 4659
rect 3466 4486 3467 4659
rect 3382 4488 3383 4659
rect 3391 4350 3392 4489
rect 3385 4490 3386 4659
rect 3394 4350 3395 4491
rect 3388 4492 3389 4659
rect 3397 4350 3398 4493
rect 3391 4494 3392 4659
rect 3400 4350 3401 4495
rect 3042 4350 3043 4497
rect 3400 4496 3401 4659
rect 3412 4496 3413 4659
rect 3520 4350 3521 4497
rect 3415 4350 3416 4499
rect 3418 4498 3419 4659
rect 3424 4350 3425 4499
rect 3469 4498 3470 4659
rect 3424 4500 3425 4659
rect 3508 4350 3509 4501
rect 3430 4502 3431 4659
rect 3439 4350 3440 4503
rect 3433 4504 3434 4659
rect 3442 4350 3443 4505
rect 3442 4506 3443 4659
rect 3457 4350 3458 4507
rect 3445 4508 3446 4659
rect 3460 4350 3461 4509
rect 3451 4350 3452 4511
rect 3454 4510 3455 4659
rect 3460 4510 3461 4659
rect 3761 4350 3762 4511
rect 3463 4350 3464 4513
rect 3739 4350 3740 4513
rect 3472 4514 3473 4659
rect 3475 4350 3476 4515
rect 3478 4514 3479 4659
rect 3505 4350 3506 4515
rect 3481 4516 3482 4659
rect 3751 4516 3752 4659
rect 3484 4518 3485 4659
rect 3499 4350 3500 4519
rect 3487 4350 3488 4521
rect 3743 4350 3744 4521
rect 3487 4522 3488 4659
rect 3529 4350 3530 4523
rect 3490 4524 3491 4659
rect 3532 4350 3533 4525
rect 3493 4526 3494 4659
rect 3511 4350 3512 4527
rect 3499 4528 3500 4659
rect 3517 4350 3518 4529
rect 3505 4530 3506 4659
rect 3523 4350 3524 4531
rect 3508 4532 3509 4659
rect 3526 4350 3527 4533
rect 3511 4534 3512 4659
rect 3547 4350 3548 4535
rect 3517 4536 3518 4659
rect 3535 4350 3536 4537
rect 3520 4538 3521 4659
rect 3538 4350 3539 4539
rect 3523 4540 3524 4659
rect 3804 4350 3805 4541
rect 3529 4542 3530 4659
rect 3770 4350 3771 4543
rect 3532 4544 3533 4659
rect 3709 4350 3710 4545
rect 3535 4546 3536 4659
rect 3562 4350 3563 4547
rect 3541 4548 3542 4659
rect 3568 4350 3569 4549
rect 3547 4550 3548 4659
rect 3574 4350 3575 4551
rect 3553 4350 3554 4553
rect 3821 4552 3822 4659
rect 3553 4554 3554 4659
rect 3885 4350 3886 4555
rect 3556 4556 3557 4659
rect 3577 4350 3578 4557
rect 3559 4350 3560 4559
rect 3797 4350 3798 4559
rect 3559 4560 3560 4659
rect 3871 4350 3872 4561
rect 3565 4562 3566 4659
rect 3580 4350 3581 4563
rect 3571 4564 3572 4659
rect 3586 4350 3587 4565
rect 3589 4564 3590 4659
rect 3598 4350 3599 4565
rect 3595 4566 3596 4659
rect 3622 4350 3623 4567
rect 3601 4568 3602 4659
rect 3604 4350 3605 4569
rect 3613 4568 3614 4659
rect 3628 4350 3629 4569
rect 3616 4350 3617 4571
rect 3917 4350 3918 4571
rect 3625 4572 3626 4659
rect 3664 4350 3665 4573
rect 3631 4574 3632 4659
rect 3935 4574 3936 4659
rect 3634 4350 3635 4577
rect 3832 4576 3833 4659
rect 3643 4578 3644 4659
rect 3646 4350 3647 4579
rect 3649 4578 3650 4659
rect 3652 4350 3653 4579
rect 3655 4578 3656 4659
rect 3658 4350 3659 4579
rect 3667 4578 3668 4659
rect 3688 4350 3689 4579
rect 3673 4580 3674 4659
rect 3961 4350 3962 4581
rect 3682 4350 3683 4583
rect 3953 4582 3954 4659
rect 3682 4584 3683 4659
rect 3938 4350 3939 4585
rect 3685 4350 3686 4587
rect 3941 4350 3942 4587
rect 3685 4588 3686 4659
rect 3694 4350 3695 4589
rect 3691 4590 3692 4659
rect 3886 4590 3887 4659
rect 3697 4592 3698 4659
rect 3712 4350 3713 4593
rect 3703 4594 3704 4659
rect 3718 4350 3719 4595
rect 3706 4350 3707 4597
rect 3773 4350 3774 4597
rect 3610 4350 3611 4599
rect 3706 4598 3707 4659
rect 3709 4598 3710 4659
rect 3924 4350 3925 4599
rect 3721 4350 3722 4601
rect 3826 4350 3827 4601
rect 3715 4602 3716 4659
rect 3825 4602 3826 4659
rect 3733 4604 3734 4659
rect 3749 4350 3750 4605
rect 3754 4604 3755 4659
rect 3758 4350 3759 4605
rect 3757 4606 3758 4659
rect 3878 4350 3879 4607
rect 3760 4608 3761 4659
rect 3776 4350 3777 4609
rect 3577 4610 3578 4659
rect 3775 4610 3776 4659
rect 3766 4612 3767 4659
rect 3782 4350 3783 4613
rect 3769 4614 3770 4659
rect 3920 4350 3921 4615
rect 3779 4350 3780 4617
rect 3874 4350 3875 4617
rect 3787 4618 3788 4659
rect 3788 4350 3789 4619
rect 3791 4350 3792 4619
rect 3889 4618 3890 4659
rect 3790 4620 3791 4659
rect 3927 4350 3928 4621
rect 3785 4350 3786 4623
rect 3928 4622 3929 4659
rect 3784 4624 3785 4659
rect 3794 4350 3795 4625
rect 3793 4626 3794 4659
rect 3823 4350 3824 4627
rect 3805 4628 3806 4659
rect 3974 4628 3975 4659
rect 3808 4630 3809 4659
rect 3942 4630 3943 4659
rect 3811 4632 3812 4659
rect 3828 4632 3829 4659
rect 3835 4350 3836 4633
rect 3844 4632 3845 4659
rect 3856 4350 3857 4633
rect 3859 4632 3860 4659
rect 3853 4350 3854 4635
rect 3856 4634 3857 4659
rect 3670 4350 3671 4637
rect 3853 4636 3854 4659
rect 3865 4350 3866 4637
rect 3880 4636 3881 4659
rect 3868 4350 3869 4639
rect 3883 4638 3884 4659
rect 3874 4640 3875 4659
rect 3948 4350 3949 4641
rect 3661 4642 3662 4659
rect 3949 4642 3950 4659
rect 3877 4644 3878 4659
rect 3945 4350 3946 4645
rect 3898 4350 3899 4647
rect 3913 4646 3914 4659
rect 3901 4350 3902 4649
rect 3916 4648 3917 4659
rect 3850 4350 3851 4651
rect 3900 4650 3901 4659
rect 3847 4350 3848 4653
rect 3850 4652 3851 4659
rect 3904 4350 3905 4653
rect 3919 4652 3920 4659
rect 3724 4350 3725 4655
rect 3903 4654 3904 4659
rect 3907 4350 3908 4655
rect 3922 4654 3923 4659
rect 3763 4656 3764 4659
rect 3907 4656 3908 4659
rect 3951 4350 3952 4657
rect 3977 4656 3978 4659
rect 2876 4663 2877 4666
rect 3009 4663 3010 4666
rect 2869 4663 2870 4668
rect 2876 4667 2877 5010
rect 2872 4663 2873 4670
rect 3009 4669 3010 5010
rect 2885 4663 2886 4672
rect 2994 4663 2995 4672
rect 2892 4663 2893 4674
rect 3346 4663 3347 4674
rect 2896 4675 2897 5010
rect 3196 4663 3197 4676
rect 2899 4663 2900 4678
rect 3316 4663 3317 4678
rect 2903 4663 2904 4680
rect 2918 4663 2919 4680
rect 2906 4663 2907 4682
rect 3278 4681 3279 5010
rect 2912 4683 2913 5010
rect 3260 4683 3261 5010
rect 2926 4685 2927 5010
rect 3048 4663 3049 4686
rect 2936 4663 2937 4688
rect 3235 4663 3236 4688
rect 2936 4689 2937 5010
rect 3081 4663 3082 4690
rect 2940 4663 2941 4692
rect 2950 4691 2951 5010
rect 2943 4663 2944 4694
rect 3331 4663 3332 4694
rect 2947 4663 2948 4696
rect 3166 4663 3167 4696
rect 2959 4697 2960 5010
rect 3385 4663 3386 4698
rect 2961 4663 2962 4700
rect 3541 4663 3542 4700
rect 2964 4663 2965 4702
rect 3643 4663 3644 4702
rect 2973 4663 2974 4704
rect 3045 4663 3046 4704
rect 2991 4663 2992 4706
rect 3012 4705 3013 5010
rect 2979 4663 2980 4708
rect 2991 4707 2992 5010
rect 2997 4707 2998 5010
rect 2997 4663 2998 4708
rect 3003 4663 3004 4708
rect 3221 4707 3222 5010
rect 3018 4663 3019 4710
rect 3021 4709 3022 5010
rect 3024 4663 3025 4710
rect 3299 4709 3300 5010
rect 3044 4711 3045 5010
rect 3164 4711 3165 5010
rect 3047 4713 3048 5010
rect 3054 4663 3055 4714
rect 3057 4663 3058 4714
rect 3149 4713 3150 5010
rect 3065 4715 3066 5010
rect 3361 4663 3362 4716
rect 3071 4717 3072 5010
rect 3508 4663 3509 4718
rect 3078 4663 3079 4720
rect 3080 4719 3081 5010
rect 3077 4721 3078 5010
rect 3145 4663 3146 4722
rect 2903 4723 2904 5010
rect 3146 4723 3147 5010
rect 3083 4725 3084 5010
rect 3108 4663 3109 4726
rect 3090 4663 3091 4728
rect 3107 4727 3108 5010
rect 3122 4727 3123 5010
rect 3181 4663 3182 4728
rect 2933 4663 2934 4730
rect 3182 4729 3183 5010
rect 3135 4663 3136 4732
rect 3217 4663 3218 4732
rect 3120 4663 3121 4734
rect 3134 4733 3135 5010
rect 3119 4735 3120 5010
rect 3178 4663 3179 4736
rect 3139 4663 3140 4738
rect 3520 4663 3521 4738
rect 3126 4663 3127 4740
rect 3140 4739 3141 5010
rect 3096 4663 3097 4742
rect 3125 4741 3126 5010
rect 3154 4663 3155 4742
rect 3490 4663 3491 4742
rect 3158 4743 3159 5010
rect 3205 4663 3206 4744
rect 3170 4745 3171 5010
rect 3433 4663 3434 4746
rect 3176 4747 3177 5010
rect 3241 4663 3242 4748
rect 3188 4749 3189 5010
rect 3229 4663 3230 4750
rect 3190 4663 3191 4752
rect 3197 4751 3198 5010
rect 3194 4753 3195 5010
rect 3265 4663 3266 4754
rect 3036 4663 3037 4756
rect 3266 4755 3267 5010
rect 3037 4757 3038 5010
rect 3344 4757 3345 5010
rect 3203 4759 3204 5010
rect 3280 4663 3281 4760
rect 3209 4761 3210 5010
rect 3253 4663 3254 4762
rect 3215 4763 3216 5010
rect 3292 4663 3293 4764
rect 3027 4663 3028 4766
rect 3293 4765 3294 5010
rect 3027 4767 3028 5010
rect 3286 4663 3287 4768
rect 3223 4663 3224 4770
rect 3458 4769 3459 5010
rect 3230 4771 3231 5010
rect 3502 4663 3503 4772
rect 3233 4773 3234 5010
rect 3304 4663 3305 4774
rect 2957 4663 2958 4776
rect 3305 4775 3306 5010
rect 3245 4777 3246 5010
rect 3340 4663 3341 4778
rect 3247 4663 3248 4780
rect 3380 4779 3381 5010
rect 3251 4781 3252 5010
rect 3334 4663 3335 4782
rect 3257 4783 3258 5010
rect 3358 4663 3359 4784
rect 3268 4663 3269 4786
rect 3772 4663 3773 4786
rect 3269 4787 3270 5010
rect 3352 4663 3353 4788
rect 3274 4663 3275 4790
rect 3750 4789 3751 5010
rect 3275 4791 3276 5010
rect 3382 4663 3383 4792
rect 3281 4793 3282 5010
rect 3370 4663 3371 4794
rect 3132 4663 3133 4796
rect 3371 4795 3372 5010
rect 2886 4797 2887 5010
rect 3131 4797 3132 5010
rect 3295 4663 3296 4798
rect 3308 4797 3309 5010
rect 3302 4799 3303 5010
rect 3391 4663 3392 4800
rect 3310 4663 3311 4802
rect 3398 4801 3399 5010
rect 3311 4803 3312 5010
rect 3442 4663 3443 4804
rect 3314 4805 3315 5010
rect 3445 4663 3446 4806
rect 3317 4807 3318 5010
rect 3406 4663 3407 4808
rect 3320 4809 3321 5010
rect 3409 4663 3410 4810
rect 3322 4663 3323 4812
rect 3599 4811 3600 5010
rect 3199 4663 3200 4814
rect 3323 4813 3324 5010
rect 3335 4813 3336 5010
rect 3466 4663 3467 4814
rect 3338 4815 3339 5010
rect 3469 4663 3470 4816
rect 3341 4817 3342 5010
rect 3430 4663 3431 4818
rect 3347 4819 3348 5010
rect 3412 4663 3413 4820
rect 3353 4821 3354 5010
rect 3484 4663 3485 4822
rect 3356 4823 3357 5010
rect 3418 4663 3419 4824
rect 3362 4825 3363 5010
rect 3493 4663 3494 4826
rect 3374 4827 3375 5010
rect 3505 4663 3506 4828
rect 3377 4829 3378 5010
rect 3772 4829 3773 5010
rect 3386 4831 3387 5010
rect 3517 4663 3518 4832
rect 3388 4663 3389 4834
rect 3739 4663 3740 4834
rect 3142 4663 3143 4836
rect 3389 4835 3390 5010
rect 3404 4835 3405 5010
rect 3671 4835 3672 5010
rect 3416 4837 3417 5010
rect 3424 4663 3425 4838
rect 3422 4839 3423 5010
rect 3553 4663 3554 4840
rect 3428 4841 3429 5010
rect 3472 4663 3473 4842
rect 3431 4843 3432 5010
rect 3481 4663 3482 4844
rect 3434 4845 3435 5010
rect 3535 4663 3536 4846
rect 3446 4847 3447 5010
rect 3454 4663 3455 4848
rect 3452 4849 3453 5010
rect 3896 4663 3897 4850
rect 3460 4663 3461 4852
rect 3699 4851 3700 5010
rect 3464 4853 3465 5010
rect 3583 4663 3584 4854
rect 3476 4855 3477 5010
rect 3939 4663 3940 4856
rect 3482 4857 3483 5010
rect 3571 4663 3572 4858
rect 3494 4859 3495 5010
rect 3589 4663 3590 4860
rect 3506 4861 3507 5010
rect 3595 4663 3596 4862
rect 3523 4663 3524 4864
rect 3775 4663 3776 4864
rect 3524 4865 3525 5010
rect 3631 4663 3632 4866
rect 3532 4663 3533 4868
rect 3659 4867 3660 5010
rect 3536 4869 3537 5010
rect 3649 4663 3650 4870
rect 3542 4871 3543 5010
rect 3655 4663 3656 4872
rect 3529 4663 3530 4874
rect 3656 4873 3657 5010
rect 3530 4875 3531 5010
rect 3625 4663 3626 4876
rect 3547 4663 3548 4878
rect 3596 4877 3597 5010
rect 3548 4879 3549 5010
rect 3661 4663 3662 4880
rect 3554 4881 3555 5010
rect 3673 4663 3674 4882
rect 3556 4663 3557 4884
rect 3593 4883 3594 5010
rect 3367 4663 3368 4886
rect 3557 4885 3558 5010
rect 3368 4887 3369 5010
rect 3499 4663 3500 4888
rect 3500 4889 3501 5010
rect 3559 4663 3560 4890
rect 3262 4663 3263 4892
rect 3560 4891 3561 5010
rect 3263 4893 3264 5010
rect 3328 4663 3329 4894
rect 3329 4895 3330 5010
rect 3400 4663 3401 4896
rect 3401 4897 3402 5010
rect 3487 4663 3488 4898
rect 3488 4899 3489 5010
rect 3601 4663 3602 4900
rect 3563 4901 3564 5010
rect 3667 4663 3668 4902
rect 3364 4663 3365 4904
rect 3668 4903 3669 5010
rect 3565 4663 3566 4906
rect 3782 4905 3783 5010
rect 3569 4907 3570 5010
rect 3853 4663 3854 4908
rect 3577 4663 3578 4910
rect 3893 4663 3894 4910
rect 3587 4911 3588 5010
rect 3685 4663 3686 4912
rect 3605 4913 3606 5010
rect 3709 4663 3710 4914
rect 3478 4663 3479 4916
rect 3708 4915 3709 5010
rect 3611 4917 3612 5010
rect 3775 4917 3776 5010
rect 3623 4919 3624 5010
rect 3960 4663 3961 4920
rect 3629 4921 3630 5010
rect 3733 4663 3734 4922
rect 3632 4923 3633 5010
rect 3769 4663 3770 4924
rect 3511 4663 3512 4926
rect 3768 4925 3769 5010
rect 3512 4927 3513 5010
rect 3613 4663 3614 4928
rect 3638 4927 3639 5010
rect 3697 4663 3698 4928
rect 3644 4929 3645 5010
rect 3900 4663 3901 4930
rect 3581 4931 3582 5010
rect 3899 4931 3900 5010
rect 3662 4933 3663 5010
rect 3703 4663 3704 4934
rect 3665 4935 3666 5010
rect 3706 4663 3707 4936
rect 3678 4937 3679 5010
rect 3846 4937 3847 5010
rect 3682 4663 3683 4940
rect 3932 4663 3933 4940
rect 3691 4663 3692 4942
rect 3839 4941 3840 5010
rect 3693 4943 3694 5010
rect 3983 4663 3984 4944
rect 3696 4945 3697 5010
rect 3754 4663 3755 4946
rect 3702 4947 3703 5010
rect 3928 4663 3929 4948
rect 3715 4663 3716 4950
rect 3832 4663 3833 4950
rect 3714 4951 3715 5010
rect 3760 4663 3761 4952
rect 3717 4953 3718 5010
rect 3903 4663 3904 4954
rect 3726 4955 3727 5010
rect 3766 4663 3767 4956
rect 3419 4957 3420 5010
rect 3765 4957 3766 5010
rect 3738 4959 3739 5010
rect 3787 4663 3788 4960
rect 3741 4961 3742 5010
rect 3790 4663 3791 4962
rect 3744 4963 3745 5010
rect 3863 4963 3864 5010
rect 3757 4663 3758 4966
rect 3828 4663 3829 4966
rect 3759 4967 3760 5010
rect 3922 4663 3923 4968
rect 3763 4663 3764 4970
rect 3835 4663 3836 4970
rect 3762 4971 3763 5010
rect 3793 4663 3794 4972
rect 3779 4973 3780 5010
rect 3886 4663 3887 4974
rect 3797 4975 3798 5010
rect 3893 4975 3894 5010
rect 3800 4977 3801 5010
rect 3902 4977 3903 5010
rect 3803 4979 3804 5010
rect 3844 4663 3845 4980
rect 3805 4663 3806 4982
rect 3909 4981 3910 5010
rect 3808 4663 3809 4984
rect 3970 4663 3971 4984
rect 3809 4985 3810 5010
rect 3856 4663 3857 4986
rect 3812 4987 3813 5010
rect 3859 4663 3860 4988
rect 3821 4989 3822 5010
rect 3874 4663 3875 4990
rect 3824 4991 3825 5010
rect 3877 4663 3878 4992
rect 3833 4993 3834 5010
rect 3880 4663 3881 4994
rect 3836 4995 3837 5010
rect 3883 4663 3884 4996
rect 3729 4997 3730 5010
rect 3882 4997 3883 5010
rect 3850 4663 3851 5000
rect 3896 4999 3897 5010
rect 3866 5001 3867 5010
rect 3913 4663 3914 5002
rect 3784 4663 3785 5004
rect 3912 5003 3913 5010
rect 3747 5005 3748 5010
rect 3785 5005 3786 5010
rect 3869 5005 3870 5010
rect 3916 4663 3917 5006
rect 3889 5007 3890 5010
rect 3919 4663 3920 5008
rect 3935 4663 3936 5008
rect 3967 4663 3968 5008
rect 2863 5014 2864 5017
rect 2876 5014 2877 5017
rect 2870 5014 2871 5019
rect 3009 5014 3010 5019
rect 2873 5014 2874 5021
rect 3047 5014 3048 5021
rect 2879 5014 2880 5023
rect 3194 5014 3195 5023
rect 2882 5014 2883 5025
rect 3012 5014 3013 5025
rect 2896 5014 2897 5027
rect 3131 5014 3132 5027
rect 2905 5028 2906 5319
rect 3275 5014 3276 5029
rect 2912 5030 2913 5319
rect 3146 5014 3147 5031
rect 2922 5014 2923 5033
rect 3149 5014 3150 5033
rect 2922 5034 2923 5319
rect 3278 5014 3279 5035
rect 2919 5014 2920 5037
rect 3279 5036 3280 5319
rect 2929 5014 2930 5039
rect 3335 5014 3336 5039
rect 2933 5014 2934 5041
rect 3069 5040 3070 5319
rect 2940 5014 2941 5043
rect 3311 5014 3312 5043
rect 2941 5044 2942 5319
rect 2950 5014 2951 5045
rect 2947 5014 2948 5047
rect 3263 5014 3264 5047
rect 2960 5048 2961 5319
rect 3386 5014 3387 5049
rect 2973 5014 2974 5051
rect 3221 5014 3222 5051
rect 2972 5052 2973 5319
rect 3192 5052 3193 5319
rect 2988 5054 2989 5319
rect 2991 5014 2992 5055
rect 2994 5054 2995 5319
rect 2997 5014 2998 5055
rect 3000 5054 3001 5319
rect 3308 5014 3309 5055
rect 3003 5014 3004 5057
rect 3317 5014 3318 5057
rect 3006 5014 3007 5059
rect 3027 5014 3028 5059
rect 3012 5060 3013 5319
rect 3021 5014 3022 5061
rect 3021 5062 3022 5319
rect 3125 5014 3126 5063
rect 3037 5014 3038 5065
rect 3164 5014 3165 5065
rect 3041 5014 3042 5067
rect 3140 5014 3141 5067
rect 2893 5014 2894 5069
rect 3141 5068 3142 5319
rect 3018 5070 3019 5319
rect 3042 5070 3043 5319
rect 3044 5014 3045 5071
rect 3071 5014 3072 5071
rect 3048 5072 3049 5319
rect 3107 5014 3108 5073
rect 3057 5074 3058 5319
rect 3269 5014 3270 5075
rect 2979 5076 2980 5319
rect 3270 5076 3271 5319
rect 3060 5078 3061 5319
rect 3065 5014 3066 5079
rect 3066 5080 3067 5319
rect 3080 5014 3081 5081
rect 3077 5014 3078 5083
rect 3114 5082 3115 5319
rect 3078 5084 3079 5319
rect 3083 5014 3084 5085
rect 3102 5084 3103 5319
rect 3134 5014 3135 5085
rect 3119 5014 3120 5087
rect 3129 5086 3130 5319
rect 3122 5014 3123 5089
rect 3132 5088 3133 5319
rect 3156 5088 3157 5319
rect 3170 5014 3171 5089
rect 3158 5014 3159 5091
rect 3162 5090 3163 5319
rect 3168 5090 3169 5319
rect 3197 5014 3198 5091
rect 3180 5092 3181 5319
rect 3182 5014 3183 5093
rect 3183 5094 3184 5319
rect 3266 5014 3267 5095
rect 3198 5096 3199 5319
rect 3458 5014 3459 5097
rect 3203 5014 3204 5099
rect 3240 5098 3241 5319
rect 3108 5100 3109 5319
rect 3204 5100 3205 5319
rect 3219 5100 3220 5319
rect 3320 5014 3321 5101
rect 3222 5102 3223 5319
rect 3371 5014 3372 5103
rect 3227 5014 3228 5105
rect 3372 5104 3373 5319
rect 3231 5106 3232 5319
rect 3560 5014 3561 5107
rect 3233 5014 3234 5109
rect 3273 5108 3274 5319
rect 3030 5014 3031 5111
rect 3234 5110 3235 5319
rect 3030 5112 3031 5319
rect 3096 5112 3097 5319
rect 3243 5112 3244 5319
rect 3314 5014 3315 5113
rect 3245 5014 3246 5115
rect 3675 5014 3676 5115
rect 3246 5116 3247 5319
rect 3380 5014 3381 5117
rect 3249 5118 3250 5319
rect 3389 5014 3390 5119
rect 3251 5014 3252 5121
rect 3291 5120 3292 5319
rect 3215 5014 3216 5123
rect 3252 5122 3253 5319
rect 3209 5014 3210 5125
rect 3216 5124 3217 5319
rect 3176 5014 3177 5127
rect 3210 5126 3211 5319
rect 3257 5014 3258 5127
rect 3309 5126 3310 5319
rect 3260 5014 3261 5129
rect 3312 5128 3313 5319
rect 3281 5014 3282 5131
rect 3321 5130 3322 5319
rect 2919 5132 2920 5319
rect 3282 5132 3283 5319
rect 3297 5132 3298 5319
rect 3404 5014 3405 5133
rect 3299 5014 3300 5135
rect 3315 5134 3316 5319
rect 3300 5136 3301 5319
rect 3557 5014 3558 5137
rect 3302 5014 3303 5139
rect 3318 5138 3319 5319
rect 3293 5014 3294 5141
rect 3303 5140 3304 5319
rect 3323 5014 3324 5141
rect 3722 5140 3723 5319
rect 3324 5142 3325 5319
rect 3338 5014 3339 5143
rect 3327 5144 3328 5319
rect 3599 5014 3600 5145
rect 3333 5146 3334 5319
rect 3446 5014 3447 5147
rect 3339 5148 3340 5319
rect 3347 5014 3348 5149
rect 3188 5014 3189 5151
rect 3348 5150 3349 5319
rect 3344 5014 3345 5153
rect 3360 5152 3361 5319
rect 3305 5014 3306 5155
rect 3345 5154 3346 5319
rect 3351 5154 3352 5319
rect 3356 5014 3357 5155
rect 3329 5014 3330 5157
rect 3357 5156 3358 5319
rect 3353 5014 3354 5159
rect 3393 5158 3394 5319
rect 3362 5014 3363 5161
rect 3408 5160 3409 5319
rect 3363 5162 3364 5319
rect 3659 5014 3660 5163
rect 3368 5014 3369 5165
rect 3678 5014 3679 5165
rect 3369 5166 3370 5319
rect 3431 5014 3432 5167
rect 3374 5014 3375 5169
rect 3414 5168 3415 5319
rect 3381 5170 3382 5319
rect 3611 5014 3612 5171
rect 3387 5172 3388 5319
rect 3782 5014 3783 5173
rect 3398 5014 3399 5175
rect 3432 5174 3433 5319
rect 3401 5014 3402 5177
rect 3429 5176 3430 5319
rect 3416 5014 3417 5179
rect 3636 5178 3637 5319
rect 3377 5014 3378 5181
rect 3417 5180 3418 5319
rect 3419 5014 3420 5181
rect 3426 5180 3427 5319
rect 3420 5182 3421 5319
rect 3817 5182 3818 5319
rect 3434 5014 3435 5185
rect 3459 5184 3460 5319
rect 3438 5186 3439 5319
rect 3775 5014 3776 5187
rect 3447 5188 3448 5319
rect 3708 5014 3709 5189
rect 3450 5190 3451 5319
rect 3656 5014 3657 5191
rect 3468 5192 3469 5319
rect 3842 5014 3843 5193
rect 3471 5194 3472 5319
rect 3665 5014 3666 5195
rect 3480 5196 3481 5319
rect 3662 5014 3663 5197
rect 3488 5014 3489 5199
rect 3519 5198 3520 5319
rect 3489 5200 3490 5319
rect 3711 5014 3712 5201
rect 3435 5202 3436 5319
rect 3711 5202 3712 5319
rect 3530 5014 3531 5205
rect 3779 5014 3780 5205
rect 3512 5014 3513 5207
rect 3531 5206 3532 5319
rect 3542 5014 3543 5207
rect 3561 5206 3562 5319
rect 3543 5208 3544 5319
rect 3838 5208 3839 5319
rect 3554 5014 3555 5211
rect 3585 5210 3586 5319
rect 3536 5014 3537 5213
rect 3555 5212 3556 5319
rect 3537 5214 3538 5319
rect 3638 5014 3639 5215
rect 3563 5014 3564 5217
rect 3579 5216 3580 5319
rect 3581 5014 3582 5217
rect 3768 5216 3769 5319
rect 3587 5014 3588 5219
rect 3687 5218 3688 5319
rect 3593 5014 3594 5221
rect 3671 5014 3672 5221
rect 3569 5014 3570 5223
rect 3594 5222 3595 5319
rect 3612 5222 3613 5319
rect 3747 5014 3748 5223
rect 3623 5014 3624 5225
rect 3902 5014 3903 5225
rect 3605 5014 3606 5227
rect 3624 5226 3625 5319
rect 3629 5014 3630 5227
rect 3648 5226 3649 5319
rect 3632 5014 3633 5229
rect 3875 5014 3876 5229
rect 3642 5230 3643 5319
rect 3702 5014 3703 5231
rect 3657 5232 3658 5319
rect 3714 5014 3715 5233
rect 3422 5014 3423 5235
rect 3715 5234 3716 5319
rect 3660 5236 3661 5319
rect 3831 5236 3832 5319
rect 3669 5238 3670 5319
rect 3726 5014 3727 5239
rect 3672 5240 3673 5319
rect 3729 5014 3730 5241
rect 3500 5014 3501 5243
rect 3729 5242 3730 5319
rect 3464 5014 3465 5245
rect 3501 5244 3502 5319
rect 3465 5246 3466 5319
rect 3596 5014 3597 5247
rect 3675 5246 3676 5319
rect 3696 5014 3697 5247
rect 3678 5248 3679 5319
rect 3732 5248 3733 5319
rect 3681 5250 3682 5319
rect 3744 5014 3745 5251
rect 3684 5252 3685 5319
rect 3741 5014 3742 5253
rect 3693 5014 3694 5255
rect 3912 5014 3913 5255
rect 3699 5014 3700 5257
rect 3772 5014 3773 5257
rect 3702 5258 3703 5319
rect 3759 5014 3760 5259
rect 3705 5260 3706 5319
rect 3762 5014 3763 5261
rect 3717 5014 3718 5263
rect 3863 5014 3864 5263
rect 3441 5264 3442 5319
rect 3718 5264 3719 5319
rect 3725 5264 3726 5319
rect 3806 5264 3807 5319
rect 3735 5266 3736 5319
rect 3785 5014 3786 5267
rect 3738 5014 3739 5269
rect 3853 5014 3854 5269
rect 3747 5270 3748 5319
rect 3797 5014 3798 5271
rect 3644 5014 3645 5273
rect 3796 5272 3797 5319
rect 3750 5274 3751 5319
rect 3800 5014 3801 5275
rect 3588 5276 3589 5319
rect 3799 5276 3800 5319
rect 3753 5278 3754 5319
rect 3869 5014 3870 5279
rect 3759 5280 3760 5319
rect 3803 5014 3804 5281
rect 3567 5282 3568 5319
rect 3803 5282 3804 5319
rect 3765 5284 3766 5319
rect 3821 5014 3822 5285
rect 3630 5286 3631 5319
rect 3820 5286 3821 5319
rect 3771 5288 3772 5319
rect 3809 5014 3810 5289
rect 3476 5014 3477 5291
rect 3810 5290 3811 5319
rect 3477 5292 3478 5319
rect 3482 5014 3483 5293
rect 3452 5014 3453 5295
rect 3483 5294 3484 5319
rect 3453 5296 3454 5319
rect 3494 5014 3495 5297
rect 3495 5298 3496 5319
rect 3506 5014 3507 5299
rect 3507 5300 3508 5319
rect 3856 5014 3857 5301
rect 3774 5302 3775 5319
rect 3846 5014 3847 5303
rect 3756 5304 3757 5319
rect 3845 5304 3846 5319
rect 3783 5306 3784 5319
rect 3833 5014 3834 5307
rect 3786 5308 3787 5319
rect 3836 5014 3837 5309
rect 3812 5014 3813 5311
rect 3849 5014 3850 5311
rect 3341 5014 3342 5313
rect 3813 5312 3814 5319
rect 3824 5014 3825 5313
rect 3896 5014 3897 5313
rect 3827 5314 3828 5319
rect 3866 5014 3867 5315
rect 3834 5316 3835 5319
rect 3889 5014 3890 5317
rect 2884 5325 2885 5618
rect 3270 5323 3271 5326
rect 2888 5327 2889 5618
rect 3141 5323 3142 5328
rect 2891 5329 2892 5618
rect 2895 5329 2896 5618
rect 2908 5323 2909 5330
rect 3210 5323 3211 5330
rect 2912 5323 2913 5332
rect 2922 5323 2923 5332
rect 2911 5333 2912 5618
rect 3129 5323 3130 5334
rect 2929 5323 2930 5336
rect 2934 5335 2935 5618
rect 2941 5335 2942 5618
rect 3211 5335 3212 5618
rect 2945 5323 2946 5338
rect 3180 5323 3181 5338
rect 2965 5339 2966 5618
rect 3229 5339 3230 5618
rect 2969 5323 2970 5342
rect 3042 5323 3043 5342
rect 2972 5323 2973 5344
rect 3348 5323 3349 5344
rect 2975 5345 2976 5618
rect 3102 5323 3103 5346
rect 2979 5323 2980 5348
rect 3765 5323 3766 5348
rect 2984 5349 2985 5618
rect 2988 5323 2989 5350
rect 2990 5349 2991 5618
rect 2994 5323 2995 5350
rect 2996 5349 2997 5618
rect 3048 5323 3049 5350
rect 2999 5351 3000 5618
rect 3042 5351 3043 5618
rect 3003 5323 3004 5354
rect 3381 5323 3382 5354
rect 3008 5355 3009 5618
rect 3012 5323 3013 5356
rect 3018 5323 3019 5356
rect 3318 5323 3319 5356
rect 3021 5323 3022 5358
rect 3268 5357 3269 5618
rect 3020 5359 3021 5618
rect 3114 5323 3115 5360
rect 3023 5361 3024 5618
rect 3096 5323 3097 5362
rect 3030 5323 3031 5364
rect 3360 5323 3361 5364
rect 3030 5365 3031 5618
rect 3187 5365 3188 5618
rect 3036 5367 3037 5618
rect 3060 5323 3061 5368
rect 3048 5369 3049 5618
rect 3066 5323 3067 5370
rect 3054 5323 3055 5372
rect 3385 5371 3386 5618
rect 3054 5373 3055 5618
rect 3078 5323 3079 5374
rect 3069 5323 3070 5376
rect 3208 5375 3209 5618
rect 3072 5377 3073 5618
rect 3286 5377 3287 5618
rect 3075 5379 3076 5618
rect 3417 5323 3418 5380
rect 3099 5381 3100 5618
rect 3400 5381 3401 5618
rect 3106 5383 3107 5618
rect 3175 5383 3176 5618
rect 3111 5323 3112 5386
rect 3369 5323 3370 5386
rect 3115 5387 3116 5618
rect 3204 5323 3205 5388
rect 2922 5389 2923 5618
rect 3205 5389 3206 5618
rect 3121 5391 3122 5618
rect 3162 5323 3163 5392
rect 3132 5323 3133 5394
rect 3178 5393 3179 5618
rect 3144 5323 3145 5396
rect 3357 5323 3358 5396
rect 3145 5397 3146 5618
rect 3168 5323 3169 5398
rect 3147 5323 3148 5400
rect 3781 5399 3782 5618
rect 3151 5401 3152 5618
rect 3240 5323 3241 5402
rect 2960 5323 2961 5404
rect 3241 5403 3242 5618
rect 3154 5405 3155 5618
rect 3243 5323 3244 5406
rect 3160 5407 3161 5618
rect 3219 5323 3220 5408
rect 3163 5409 3164 5618
rect 3252 5323 3253 5410
rect 3169 5411 3170 5618
rect 3279 5323 3280 5412
rect 3172 5413 3173 5618
rect 3282 5323 3283 5414
rect 3057 5323 3058 5416
rect 3283 5415 3284 5618
rect 3181 5417 3182 5618
rect 3309 5323 3310 5418
rect 3156 5323 3157 5420
rect 3310 5419 3311 5618
rect 3157 5421 3158 5618
rect 3216 5323 3217 5422
rect 3183 5323 3184 5424
rect 3214 5423 3215 5618
rect 3184 5425 3185 5618
rect 3312 5323 3313 5426
rect 3192 5323 3193 5428
rect 3244 5427 3245 5618
rect 3193 5429 3194 5618
rect 3234 5323 3235 5430
rect 3217 5431 3218 5618
rect 3321 5323 3322 5432
rect 3220 5433 3221 5618
rect 3324 5323 3325 5434
rect 3222 5323 3223 5436
rect 3223 5435 3224 5618
rect 3226 5435 3227 5618
rect 3514 5435 3515 5618
rect 3235 5437 3236 5618
rect 3345 5323 3346 5438
rect 3246 5323 3247 5440
rect 3319 5439 3320 5618
rect 3247 5441 3248 5618
rect 3393 5323 3394 5442
rect 3249 5323 3250 5444
rect 3397 5443 3398 5618
rect 3033 5445 3034 5618
rect 3250 5445 3251 5618
rect 3253 5445 3254 5618
rect 3291 5323 3292 5446
rect 3259 5447 3260 5618
rect 3303 5323 3304 5448
rect 3265 5449 3266 5618
rect 3315 5323 3316 5450
rect 3271 5451 3272 5618
rect 3414 5323 3415 5452
rect 3277 5453 3278 5618
rect 3408 5323 3409 5454
rect 3289 5455 3290 5618
rect 3333 5323 3334 5456
rect 3295 5457 3296 5618
rect 3429 5323 3430 5458
rect 3300 5323 3301 5460
rect 3610 5459 3611 5618
rect 3313 5461 3314 5618
rect 3690 5323 3691 5462
rect 3325 5463 3326 5618
rect 3351 5323 3352 5464
rect 3331 5465 3332 5618
rect 3447 5323 3448 5466
rect 3337 5467 3338 5618
rect 3426 5323 3427 5468
rect 3339 5323 3340 5470
rect 3349 5469 3350 5618
rect 3355 5469 3356 5618
rect 3489 5323 3490 5470
rect 3361 5471 3362 5618
rect 3459 5323 3460 5472
rect 3363 5323 3364 5474
rect 3622 5473 3623 5618
rect 3367 5475 3368 5618
rect 3483 5323 3484 5476
rect 3391 5477 3392 5618
rect 3501 5323 3502 5478
rect 3297 5323 3298 5480
rect 3502 5479 3503 5618
rect 3409 5481 3410 5618
rect 3519 5323 3520 5482
rect 3424 5483 3425 5618
rect 3432 5323 3433 5484
rect 3433 5485 3434 5618
rect 3507 5323 3508 5486
rect 3435 5323 3436 5488
rect 3655 5487 3656 5618
rect 3450 5323 3451 5490
rect 3743 5489 3744 5618
rect 3451 5491 3452 5618
rect 3531 5323 3532 5492
rect 3453 5323 3454 5494
rect 3553 5493 3554 5618
rect 3463 5495 3464 5618
rect 3549 5323 3550 5496
rect 3441 5323 3442 5498
rect 3550 5497 3551 5618
rect 3465 5323 3466 5500
rect 3634 5499 3635 5618
rect 3471 5323 3472 5502
rect 3732 5323 3733 5502
rect 3475 5503 3476 5618
rect 3555 5323 3556 5504
rect 3420 5323 3421 5506
rect 3556 5505 3557 5618
rect 3421 5507 3422 5618
rect 3718 5323 3719 5508
rect 3480 5323 3481 5510
rect 3799 5323 3800 5510
rect 3481 5511 3482 5618
rect 3874 5511 3875 5618
rect 3487 5513 3488 5618
rect 3585 5323 3586 5514
rect 3490 5515 3491 5618
rect 3561 5323 3562 5516
rect 3495 5323 3496 5518
rect 3792 5323 3793 5518
rect 3387 5323 3388 5520
rect 3496 5519 3497 5618
rect 3372 5323 3373 5522
rect 3388 5521 3389 5618
rect 3373 5523 3374 5618
rect 3715 5323 3716 5524
rect 3508 5525 3509 5618
rect 3525 5323 3526 5526
rect 3532 5525 3533 5618
rect 3750 5323 3751 5526
rect 3343 5527 3344 5618
rect 3750 5527 3751 5618
rect 3535 5529 3536 5618
rect 3594 5323 3595 5530
rect 3541 5531 3542 5618
rect 3852 5323 3853 5532
rect 3562 5533 3563 5618
rect 3789 5323 3790 5534
rect 3567 5323 3568 5536
rect 3871 5535 3872 5618
rect 3198 5323 3199 5538
rect 3568 5537 3569 5618
rect 3199 5539 3200 5618
rect 3273 5323 3274 5540
rect 3574 5539 3575 5618
rect 3834 5323 3835 5540
rect 3583 5541 3584 5618
rect 3636 5323 3637 5542
rect 3588 5323 3589 5544
rect 3598 5543 3599 5618
rect 3624 5323 3625 5544
rect 3853 5543 3854 5618
rect 3327 5323 3328 5546
rect 3625 5545 3626 5618
rect 3628 5545 3629 5618
rect 3884 5545 3885 5618
rect 3642 5323 3643 5548
rect 3878 5547 3879 5618
rect 3612 5323 3613 5550
rect 3643 5549 3644 5618
rect 3231 5323 3232 5552
rect 3613 5551 3614 5618
rect 3648 5323 3649 5552
rect 3841 5323 3842 5552
rect 3301 5553 3302 5618
rect 3649 5553 3650 5618
rect 3657 5323 3658 5554
rect 3692 5553 3693 5618
rect 3438 5323 3439 5556
rect 3658 5555 3659 5618
rect 3660 5323 3661 5556
rect 3835 5555 3836 5618
rect 3661 5557 3662 5618
rect 3820 5323 3821 5558
rect 3537 5323 3538 5560
rect 3821 5559 3822 5618
rect 3538 5561 3539 5618
rect 3768 5323 3769 5562
rect 3672 5323 3673 5564
rect 3689 5563 3690 5618
rect 3675 5323 3676 5566
rect 3737 5565 3738 5618
rect 3678 5323 3679 5568
rect 3707 5567 3708 5618
rect 3681 5323 3682 5570
rect 3698 5569 3699 5618
rect 3684 5323 3685 5572
rect 3713 5571 3714 5618
rect 3687 5323 3688 5574
rect 3716 5573 3717 5618
rect 3669 5323 3670 5576
rect 3686 5575 3687 5618
rect 3695 5575 3696 5618
rect 3832 5575 3833 5618
rect 3705 5323 3706 5578
rect 3725 5577 3726 5618
rect 3735 5323 3736 5578
rect 3857 5577 3858 5618
rect 3747 5323 3748 5580
rect 3845 5323 3846 5580
rect 3415 5581 3416 5618
rect 3746 5581 3747 5618
rect 3753 5323 3754 5582
rect 3769 5581 3770 5618
rect 3756 5323 3757 5584
rect 3763 5583 3764 5618
rect 3427 5585 3428 5618
rect 3757 5585 3758 5618
rect 3771 5323 3772 5586
rect 3793 5585 3794 5618
rect 3774 5323 3775 5588
rect 3796 5587 3797 5618
rect 3477 5323 3478 5590
rect 3775 5589 3776 5618
rect 3778 5589 3779 5618
rect 3811 5589 3812 5618
rect 3783 5323 3784 5592
rect 3805 5591 3806 5618
rect 3702 5323 3703 5594
rect 3784 5593 3785 5618
rect 3701 5595 3702 5618
rect 3861 5323 3862 5596
rect 3786 5323 3787 5598
rect 3808 5597 3809 5618
rect 3759 5323 3760 5600
rect 3787 5599 3788 5618
rect 3307 5601 3308 5618
rect 3760 5601 3761 5618
rect 3824 5323 3825 5602
rect 3847 5601 3848 5618
rect 3630 5323 3631 5604
rect 3825 5603 3826 5618
rect 3468 5323 3469 5606
rect 3631 5605 3632 5618
rect 3469 5607 3470 5618
rect 3677 5607 3678 5618
rect 3827 5323 3828 5608
rect 3844 5607 3845 5618
rect 3867 5323 3868 5608
rect 3887 5607 3888 5618
rect 3543 5323 3544 5610
rect 3867 5609 3868 5618
rect 3544 5611 3545 5618
rect 3579 5323 3580 5612
rect 3580 5613 3581 5618
rect 3817 5323 3818 5614
rect 3740 5615 3741 5618
rect 3818 5615 3819 5618
rect 2904 5622 2905 5625
rect 3358 5624 3359 5921
rect 2905 5626 2906 5921
rect 3778 5626 3779 5921
rect 2908 5622 2909 5629
rect 3178 5622 3179 5629
rect 2915 5622 2916 5631
rect 3214 5622 3215 5631
rect 2922 5632 2923 5921
rect 3184 5622 3185 5633
rect 2937 5622 2938 5635
rect 2951 5634 2952 5921
rect 2929 5636 2930 5921
rect 2938 5636 2939 5921
rect 2941 5622 2942 5637
rect 3295 5622 3296 5637
rect 2944 5638 2945 5921
rect 3172 5622 3173 5639
rect 2947 5640 2948 5921
rect 3418 5640 3419 5921
rect 2953 5622 2954 5643
rect 3217 5622 3218 5643
rect 2956 5622 2957 5645
rect 3127 5644 3128 5921
rect 2965 5622 2966 5647
rect 3298 5646 3299 5921
rect 2972 5648 2973 5921
rect 2996 5622 2997 5649
rect 2975 5622 2976 5651
rect 3442 5650 3443 5921
rect 2975 5652 2976 5921
rect 3205 5622 3206 5653
rect 2984 5622 2985 5655
rect 3148 5654 3149 5921
rect 2984 5656 2985 5921
rect 2990 5622 2991 5657
rect 2990 5658 2991 5921
rect 3133 5658 3134 5921
rect 3002 5660 3003 5921
rect 3008 5622 3009 5661
rect 3008 5662 3009 5921
rect 3262 5662 3263 5921
rect 3015 5664 3016 5921
rect 3346 5664 3347 5921
rect 3020 5622 3021 5667
rect 3094 5666 3095 5921
rect 3021 5668 3022 5921
rect 3042 5622 3043 5669
rect 3023 5622 3024 5671
rect 3193 5622 3194 5671
rect 3026 5622 3027 5673
rect 3217 5672 3218 5921
rect 3030 5622 3031 5675
rect 3283 5622 3284 5675
rect 3033 5622 3034 5677
rect 3472 5676 3473 5921
rect 3048 5622 3049 5679
rect 3070 5678 3071 5921
rect 3048 5680 3049 5921
rect 3490 5622 3491 5681
rect 3054 5622 3055 5683
rect 3082 5682 3083 5921
rect 3106 5622 3107 5683
rect 3220 5622 3221 5683
rect 3157 5622 3158 5685
rect 3193 5684 3194 5921
rect 3145 5622 3146 5687
rect 3157 5686 3158 5921
rect 3121 5622 3122 5689
rect 3145 5688 3146 5921
rect 3076 5690 3077 5921
rect 3121 5690 3122 5921
rect 3169 5622 3170 5691
rect 3295 5690 3296 5921
rect 3175 5622 3176 5693
rect 3340 5692 3341 5921
rect 3181 5622 3182 5695
rect 3370 5694 3371 5921
rect 3115 5622 3116 5697
rect 3181 5696 3182 5921
rect 3199 5622 3200 5697
rect 3256 5696 3257 5921
rect 3103 5622 3104 5699
rect 3199 5698 3200 5921
rect 3079 5700 3080 5921
rect 3103 5700 3104 5921
rect 3202 5700 3203 5921
rect 3421 5622 3422 5701
rect 3154 5622 3155 5703
rect 3421 5702 3422 5921
rect 3205 5704 3206 5921
rect 3568 5622 3569 5705
rect 3208 5622 3209 5707
rect 3403 5706 3404 5921
rect 3226 5622 3227 5709
rect 3670 5622 3671 5709
rect 3229 5622 3230 5711
rect 3430 5710 3431 5921
rect 3151 5622 3152 5713
rect 3229 5712 3230 5921
rect 3235 5622 3236 5713
rect 3406 5712 3407 5921
rect 3235 5714 3236 5921
rect 3385 5622 3386 5715
rect 3250 5622 3251 5717
rect 3499 5716 3500 5921
rect 3268 5622 3269 5719
rect 3316 5718 3317 5921
rect 2888 5622 2889 5721
rect 3268 5720 3269 5921
rect 3271 5622 3272 5721
rect 3520 5720 3521 5921
rect 3283 5722 3284 5921
rect 3307 5622 3308 5723
rect 3259 5622 3260 5725
rect 3307 5724 3308 5921
rect 3286 5622 3287 5727
rect 3523 5726 3524 5921
rect 3289 5622 3290 5729
rect 3334 5728 3335 5921
rect 3289 5730 3290 5921
rect 3502 5622 3503 5731
rect 3325 5622 3326 5733
rect 3364 5732 3365 5921
rect 3241 5622 3242 5735
rect 3325 5734 3326 5921
rect 2891 5622 2892 5737
rect 3241 5736 3242 5921
rect 3343 5622 3344 5737
rect 3586 5736 3587 5921
rect 2915 5738 2916 5921
rect 3343 5738 3344 5921
rect 3349 5622 3350 5739
rect 3352 5738 3353 5921
rect 3310 5622 3311 5741
rect 3349 5740 3350 5921
rect 3361 5622 3362 5741
rect 3890 5740 3891 5921
rect 3367 5622 3368 5743
rect 3604 5742 3605 5921
rect 3367 5744 3368 5921
rect 3388 5622 3389 5745
rect 3376 5746 3377 5921
rect 3469 5622 3470 5747
rect 3385 5748 3386 5921
rect 3613 5622 3614 5749
rect 3388 5750 3389 5921
rect 3625 5622 3626 5751
rect 3394 5752 3395 5921
rect 3574 5622 3575 5753
rect 3412 5754 3413 5921
rect 3957 5754 3958 5921
rect 3415 5622 3416 5757
rect 3448 5756 3449 5921
rect 3424 5622 3425 5759
rect 3674 5622 3675 5759
rect 3424 5760 3425 5921
rect 3790 5760 3791 5921
rect 3427 5622 3428 5763
rect 3574 5762 3575 5921
rect 3433 5622 3434 5765
rect 3616 5764 3617 5921
rect 3244 5622 3245 5767
rect 3433 5766 3434 5921
rect 3163 5622 3164 5769
rect 3244 5768 3245 5921
rect 3163 5770 3164 5921
rect 3187 5622 3188 5771
rect 3187 5772 3188 5921
rect 3397 5622 3398 5773
rect 3436 5772 3437 5921
rect 3496 5622 3497 5773
rect 3247 5622 3248 5775
rect 3496 5774 3497 5921
rect 3451 5622 3452 5777
rect 3640 5776 3641 5921
rect 3451 5778 3452 5921
rect 3658 5622 3659 5779
rect 3454 5780 3455 5921
rect 3825 5622 3826 5781
rect 3460 5782 3461 5921
rect 3649 5622 3650 5783
rect 3463 5622 3464 5785
rect 3664 5784 3665 5921
rect 3400 5622 3401 5787
rect 3463 5786 3464 5921
rect 2925 5622 2926 5789
rect 3400 5788 3401 5921
rect 3466 5788 3467 5921
rect 3514 5622 3515 5789
rect 3277 5622 3278 5791
rect 3514 5790 3515 5921
rect 3253 5622 3254 5793
rect 3277 5792 3278 5921
rect 3475 5622 3476 5793
rect 3658 5792 3659 5921
rect 3160 5622 3161 5795
rect 3475 5794 3476 5921
rect 3478 5794 3479 5921
rect 3911 5794 3912 5921
rect 3484 5796 3485 5921
rect 3908 5796 3909 5921
rect 3502 5798 3503 5921
rect 3556 5622 3557 5799
rect 3313 5622 3314 5801
rect 3556 5800 3557 5921
rect 3265 5622 3266 5803
rect 3313 5802 3314 5921
rect 3526 5802 3527 5921
rect 3893 5802 3894 5921
rect 3529 5804 3530 5921
rect 3580 5622 3581 5805
rect 3508 5622 3509 5807
rect 3580 5806 3581 5921
rect 3337 5622 3338 5809
rect 3508 5808 3509 5921
rect 3535 5622 3536 5809
rect 4013 5808 4014 5921
rect 3538 5622 3539 5811
rect 3864 5622 3865 5811
rect 3301 5622 3302 5813
rect 3538 5812 3539 5921
rect 3301 5814 3302 5921
rect 3850 5622 3851 5815
rect 3541 5622 3542 5817
rect 3670 5816 3671 5921
rect 3547 5818 3548 5921
rect 3610 5622 3611 5819
rect 3373 5622 3374 5821
rect 3610 5820 3611 5921
rect 3036 5622 3037 5823
rect 3373 5822 3374 5921
rect 3550 5622 3551 5823
rect 3589 5822 3590 5921
rect 3553 5822 3554 5921
rect 3553 5622 3554 5823
rect 3562 5622 3563 5825
rect 3568 5824 3569 5921
rect 3598 5622 3599 5825
rect 3730 5824 3731 5921
rect 3355 5622 3356 5827
rect 3598 5826 3599 5921
rect 3628 5622 3629 5827
rect 4030 5826 4031 5921
rect 3628 5828 3629 5921
rect 3695 5622 3696 5829
rect 3634 5622 3635 5831
rect 3745 5830 3746 5921
rect 3409 5622 3410 5833
rect 3634 5832 3635 5921
rect 3643 5622 3644 5833
rect 3748 5832 3749 5921
rect 3655 5622 3656 5835
rect 3743 5622 3744 5835
rect 3631 5622 3632 5837
rect 3742 5836 3743 5921
rect 3661 5622 3662 5839
rect 3766 5838 3767 5921
rect 3673 5840 3674 5921
rect 3960 5840 3961 5921
rect 3679 5842 3680 5921
rect 3874 5622 3875 5843
rect 3689 5622 3690 5845
rect 3799 5844 3800 5921
rect 3692 5622 3693 5847
rect 3823 5846 3824 5921
rect 3691 5848 3692 5921
rect 3871 5622 3872 5849
rect 3139 5850 3140 5921
rect 3871 5850 3872 5921
rect 3698 5622 3699 5853
rect 3820 5852 3821 5921
rect 3487 5622 3488 5855
rect 3697 5854 3698 5921
rect 3713 5622 3714 5855
rect 3862 5854 3863 5921
rect 3712 5856 3713 5921
rect 4010 5856 4011 5921
rect 3716 5622 3717 5859
rect 3811 5622 3812 5859
rect 3532 5622 3533 5861
rect 3715 5860 3716 5921
rect 3331 5622 3332 5863
rect 3532 5862 3533 5921
rect 3211 5622 3212 5865
rect 3331 5864 3332 5921
rect 3718 5864 3719 5921
rect 4017 5864 4018 5921
rect 3725 5622 3726 5867
rect 4003 5866 4004 5921
rect 3724 5868 3725 5921
rect 3814 5622 3815 5869
rect 3737 5622 3738 5871
rect 3865 5870 3866 5921
rect 3736 5872 3737 5921
rect 3935 5872 3936 5921
rect 3740 5622 3741 5875
rect 3868 5874 3869 5921
rect 3754 5876 3755 5921
rect 3828 5622 3829 5877
rect 3701 5622 3702 5879
rect 3829 5878 3830 5921
rect 3757 5622 3758 5881
rect 3884 5880 3885 5921
rect 3760 5622 3761 5883
rect 3808 5622 3809 5883
rect 3583 5622 3584 5885
rect 3760 5884 3761 5921
rect 3763 5622 3764 5885
rect 3860 5622 3861 5885
rect 3223 5622 3224 5887
rect 3859 5886 3860 5921
rect 3223 5888 3224 5921
rect 3319 5622 3320 5889
rect 3769 5622 3770 5889
rect 3914 5888 3915 5921
rect 3772 5890 3773 5921
rect 3996 5890 3997 5921
rect 3781 5622 3782 5893
rect 3926 5892 3927 5921
rect 3622 5622 3623 5895
rect 3781 5894 3782 5921
rect 3391 5622 3392 5897
rect 3622 5896 3623 5921
rect 3784 5622 3785 5897
rect 3929 5896 3930 5921
rect 3784 5898 3785 5921
rect 3887 5622 3888 5899
rect 3787 5622 3788 5901
rect 3947 5900 3948 5921
rect 3793 5622 3794 5903
rect 3938 5902 3939 5921
rect 3707 5622 3708 5905
rect 3793 5904 3794 5921
rect 3796 5622 3797 5905
rect 3941 5904 3942 5921
rect 3805 5622 3806 5907
rect 3944 5906 3945 5921
rect 3686 5622 3687 5909
rect 3805 5908 3806 5921
rect 3481 5622 3482 5911
rect 3685 5910 3686 5921
rect 3817 5910 3818 5921
rect 4020 5910 4021 5921
rect 3826 5912 3827 5921
rect 3932 5912 3933 5921
rect 3832 5622 3833 5915
rect 3841 5914 3842 5921
rect 3844 5622 3845 5915
rect 3983 5914 3984 5921
rect 3847 5622 3848 5917
rect 3986 5916 3987 5921
rect 3853 5622 3854 5919
rect 3902 5918 3903 5921
rect 3905 5918 3906 5921
rect 3989 5918 3990 5921
rect 2857 5925 2858 5928
rect 3150 5927 3151 6262
rect 2872 5929 2873 6262
rect 2879 5929 2880 6262
rect 2887 5925 2888 5930
rect 3053 5929 3054 6262
rect 2890 5925 2891 5932
rect 3277 5925 3278 5932
rect 2899 5933 2900 6262
rect 3241 5925 3242 5934
rect 2915 5925 2916 5936
rect 3117 5935 3118 6262
rect 2919 5925 2920 5938
rect 3295 5925 3296 5938
rect 2922 5925 2923 5940
rect 2926 5925 2927 5940
rect 2930 5939 2931 6262
rect 2990 5925 2991 5940
rect 2938 5925 2939 5942
rect 2939 5941 2940 6262
rect 2951 5925 2952 5942
rect 3207 5941 3208 6262
rect 2954 5925 2955 5944
rect 3331 5925 3332 5944
rect 2964 5945 2965 6262
rect 2984 5925 2985 5946
rect 2968 5925 2969 5948
rect 3279 5947 3280 6262
rect 2967 5949 2968 6262
rect 2990 5949 2991 6262
rect 2978 5951 2979 6262
rect 3499 5925 3500 5952
rect 2993 5925 2994 5954
rect 3313 5925 3314 5954
rect 2996 5955 2997 6262
rect 3127 5925 3128 5956
rect 3008 5925 3009 5958
rect 3256 5925 3257 5958
rect 3002 5925 3003 5960
rect 3008 5959 3009 6262
rect 3015 5925 3016 5960
rect 3334 5925 3335 5960
rect 3018 5925 3019 5962
rect 3264 5961 3265 6262
rect 3026 5963 3027 6262
rect 3094 5925 3095 5964
rect 3029 5965 3030 6262
rect 3070 5925 3071 5966
rect 3021 5925 3022 5968
rect 3071 5967 3072 6262
rect 3033 5925 3034 5970
rect 3163 5925 3164 5970
rect 3036 5925 3037 5972
rect 3126 5971 3127 6262
rect 3041 5973 3042 6262
rect 3082 5925 3083 5974
rect 3055 5925 3056 5976
rect 3223 5925 3224 5976
rect 3068 5977 3069 6262
rect 3273 5977 3274 6262
rect 3076 5925 3077 5980
rect 3202 5925 3203 5980
rect 3079 5925 3080 5982
rect 3385 5925 3386 5982
rect 2952 5983 2953 6262
rect 3080 5983 3081 6262
rect 3083 5983 3084 6262
rect 3139 5925 3140 5984
rect 3086 5985 3087 6262
rect 3133 5925 3134 5986
rect 2916 5987 2917 6262
rect 3132 5987 3133 6262
rect 3093 5989 3094 6262
rect 3349 5925 3350 5990
rect 3096 5991 3097 6262
rect 3145 5925 3146 5992
rect 3099 5993 3100 6262
rect 3148 5925 3149 5994
rect 3103 5925 3104 5996
rect 3540 5995 3541 6262
rect 2961 5925 2962 5998
rect 3102 5997 3103 6262
rect 3108 5997 3109 6262
rect 3298 5925 3299 5998
rect 3114 5999 3115 6262
rect 3181 5925 3182 6000
rect 3138 6001 3139 6262
rect 3343 5925 3344 6002
rect 3144 6003 3145 6262
rect 3433 5925 3434 6004
rect 3157 5925 3158 6006
rect 3787 5925 3788 6006
rect 3159 6007 3160 6262
rect 3268 5925 3269 6008
rect 3162 6009 3163 6262
rect 3229 5925 3230 6010
rect 3168 6011 3169 6262
rect 3217 5925 3218 6012
rect 3174 6013 3175 6262
rect 3193 5925 3194 6014
rect 3180 6015 3181 6262
rect 3244 5925 3245 6016
rect 3187 5925 3188 6018
rect 3935 5925 3936 6018
rect 2945 6019 2946 6262
rect 3186 6019 3187 6262
rect 3192 6019 3193 6262
rect 3463 5925 3464 6020
rect 3205 5925 3206 6022
rect 3642 6021 3643 6262
rect 3204 6023 3205 6262
rect 3340 5925 3341 6024
rect 3045 5925 3046 6026
rect 3339 6025 3340 6262
rect 3210 6027 3211 6262
rect 3262 5925 3263 6028
rect 3216 6029 3217 6262
rect 3370 5925 3371 6030
rect 3219 6031 3220 6262
rect 3373 5925 3374 6032
rect 3222 6033 3223 6262
rect 3283 5925 3284 6034
rect 3121 5925 3122 6036
rect 3282 6035 3283 6262
rect 2999 6037 3000 6262
rect 3120 6037 3121 6262
rect 3228 6037 3229 6262
rect 3358 5925 3359 6038
rect 3235 5925 3236 6040
rect 3348 6039 3349 6262
rect 3234 6041 3235 6262
rect 3325 5925 3326 6042
rect 3240 6043 3241 6262
rect 3307 5925 3308 6044
rect 3017 6045 3018 6262
rect 3306 6045 3307 6262
rect 3246 6047 3247 6262
rect 3400 5925 3401 6048
rect 3249 6049 3250 6262
rect 3403 5925 3404 6050
rect 3252 6051 3253 6262
rect 3406 5925 3407 6052
rect 3258 6053 3259 6262
rect 3418 5925 3419 6054
rect 3261 6055 3262 6262
rect 3421 5925 3422 6056
rect 3270 6057 3271 6262
rect 3346 5925 3347 6058
rect 3090 6059 3091 6262
rect 3345 6059 3346 6262
rect 3276 6061 3277 6262
rect 3430 5925 3431 6062
rect 3289 5925 3290 6064
rect 3480 6063 3481 6262
rect 3294 6065 3295 6262
rect 3472 5925 3473 6066
rect 3297 6067 3298 6262
rect 3475 5925 3476 6068
rect 3309 6069 3310 6262
rect 3316 5925 3317 6070
rect 3312 6071 3313 6262
rect 3496 5925 3497 6072
rect 3315 6073 3316 6262
rect 3442 5925 3443 6074
rect 3318 6075 3319 6262
rect 3364 5925 3365 6076
rect 3330 6077 3331 6262
rect 3514 5925 3515 6078
rect 3336 6079 3337 6262
rect 3520 5925 3521 6080
rect 3342 6081 3343 6262
rect 3460 5925 3461 6082
rect 3351 6083 3352 6262
rect 3352 5925 3353 6084
rect 3354 6083 3355 6262
rect 3702 6083 3703 6262
rect 3360 6085 3361 6262
rect 3544 5925 3545 6086
rect 3372 6087 3373 6262
rect 3556 5925 3557 6088
rect 3384 6089 3385 6262
rect 3508 5925 3509 6090
rect 3388 5925 3389 6092
rect 3699 6091 3700 6262
rect 3390 6093 3391 6262
rect 3526 5925 3527 6094
rect 3376 5925 3377 6096
rect 3525 6095 3526 6262
rect 3402 6097 3403 6262
rect 3630 6097 3631 6262
rect 3408 6099 3409 6262
rect 3610 5925 3611 6100
rect 3412 5925 3413 6102
rect 3606 6101 3607 6262
rect 3414 6103 3415 6262
rect 3598 5925 3599 6104
rect 3420 6105 3421 6262
rect 3604 5925 3605 6106
rect 3432 6107 3433 6262
rect 3484 5925 3485 6108
rect 3438 6109 3439 6262
rect 3622 5925 3623 6110
rect 3444 6111 3445 6262
rect 3932 5925 3933 6112
rect 3448 5925 3449 6114
rect 3636 6113 3637 6262
rect 3456 6115 3457 6262
rect 3634 5925 3635 6116
rect 3451 5925 3452 6118
rect 3633 6117 3634 6262
rect 3450 6119 3451 6262
rect 3616 5925 3617 6120
rect 3462 6121 3463 6262
rect 3574 5925 3575 6122
rect 3474 6123 3475 6262
rect 3960 5925 3961 6124
rect 3478 5925 3479 6126
rect 3957 5925 3958 6126
rect 3486 6127 3487 6262
rect 3658 5925 3659 6128
rect 3454 5925 3455 6130
rect 3657 6129 3658 6262
rect 3492 6131 3493 6262
rect 3670 5925 3671 6132
rect 3495 6133 3496 6262
rect 3664 5925 3665 6134
rect 3513 6135 3514 6262
rect 3685 5925 3686 6136
rect 3519 6137 3520 6262
rect 3691 5925 3692 6138
rect 3523 5925 3524 6140
rect 3705 6139 3706 6262
rect 3529 5925 3530 6142
rect 3603 6141 3604 6262
rect 3538 5925 3539 6144
rect 3760 5925 3761 6144
rect 3199 5925 3200 6146
rect 3537 6145 3538 6262
rect 3543 6145 3544 6262
rect 3652 5925 3653 6146
rect 3549 6147 3550 6262
rect 3580 5925 3581 6148
rect 3466 5925 3467 6150
rect 3579 6149 3580 6262
rect 3553 5925 3554 6152
rect 3576 6151 3577 6262
rect 3555 6153 3556 6262
rect 3712 5925 3713 6154
rect 3532 5925 3533 6156
rect 3712 6155 3713 6262
rect 3301 5925 3302 6158
rect 3531 6157 3532 6262
rect 3558 6157 3559 6262
rect 3679 5925 3680 6158
rect 3561 6159 3562 6262
rect 3673 5925 3674 6160
rect 3367 5925 3368 6162
rect 3672 6161 3673 6262
rect 3366 6163 3367 6262
rect 3424 5925 3425 6164
rect 3568 5925 3569 6164
rect 3591 6163 3592 6262
rect 3394 5925 3395 6166
rect 3567 6165 3568 6262
rect 3573 6165 3574 6262
rect 3589 5925 3590 6166
rect 3615 6165 3616 6262
rect 3724 5925 3725 6166
rect 3621 6167 3622 6262
rect 3730 5925 3731 6168
rect 3628 5925 3629 6170
rect 3874 5925 3875 6170
rect 3396 6171 3397 6262
rect 3627 6171 3628 6262
rect 3640 5925 3641 6172
rect 3893 5925 3894 6172
rect 3547 5925 3548 6174
rect 3639 6173 3640 6262
rect 3651 6173 3652 6262
rect 3748 5925 3749 6174
rect 3663 6175 3664 6262
rect 3999 5925 4000 6176
rect 3687 6177 3688 6262
rect 3754 5925 3755 6178
rect 3693 6179 3694 6262
rect 3742 5925 3743 6180
rect 3697 5925 3698 6182
rect 4037 5925 4038 6182
rect 3696 6183 3697 6262
rect 3778 5925 3779 6184
rect 3715 5925 3716 6186
rect 4013 5925 4014 6186
rect 3718 5925 3719 6188
rect 4027 5925 4028 6188
rect 3727 6189 3728 6262
rect 3805 5925 3806 6190
rect 3730 6191 3731 6262
rect 3799 5925 3800 6192
rect 3733 6193 3734 6262
rect 3817 5925 3818 6194
rect 3736 5925 3737 6196
rect 3950 5925 3951 6196
rect 3736 6197 3737 6262
rect 3823 5925 3824 6198
rect 3739 6199 3740 6262
rect 3826 5925 3827 6200
rect 3745 5925 3746 6202
rect 3890 5925 3891 6202
rect 3748 6203 3749 6262
rect 3823 6203 3824 6262
rect 3760 6205 3761 6262
rect 3859 5925 3860 6206
rect 3763 6207 3764 6262
rect 3862 5925 3863 6208
rect 3766 5925 3767 6210
rect 3996 5925 3997 6210
rect 3766 6211 3767 6262
rect 3868 5925 3869 6212
rect 3769 6213 3770 6262
rect 3793 5925 3794 6214
rect 3586 5925 3587 6216
rect 3793 6215 3794 6262
rect 3502 5925 3503 6218
rect 3585 6217 3586 6262
rect 3048 5925 3049 6220
rect 3501 6219 3502 6262
rect 3772 5925 3773 6220
rect 3814 6219 3815 6262
rect 3436 5925 3437 6222
rect 3772 6221 3773 6262
rect 3779 6221 3780 6262
rect 3790 5925 3791 6222
rect 3784 5925 3785 6224
rect 4040 5925 4041 6224
rect 3786 6225 3787 6262
rect 3865 5925 3866 6226
rect 3796 6227 3797 6262
rect 3844 6227 3845 6262
rect 3805 6229 3806 6262
rect 3938 5925 3939 6230
rect 3808 6231 3809 6262
rect 3941 5925 3942 6232
rect 3811 6233 3812 6262
rect 3926 5925 3927 6234
rect 3817 6235 3818 6262
rect 3944 5925 3945 6236
rect 3826 6237 3827 6262
rect 3841 5925 3842 6238
rect 3781 5925 3782 6240
rect 3840 6239 3841 6262
rect 3829 5925 3830 6242
rect 3853 6241 3854 6262
rect 3789 6243 3790 6262
rect 3830 6243 3831 6262
rect 3847 6243 3848 6262
rect 3905 5925 3906 6244
rect 3850 6245 3851 6262
rect 3986 5925 3987 6246
rect 3859 6247 3860 6262
rect 3884 5925 3885 6248
rect 3820 5925 3821 6250
rect 3884 6249 3885 6262
rect 3820 6251 3821 6262
rect 3947 5925 3948 6252
rect 3866 6253 3867 6262
rect 3914 5925 3915 6254
rect 3902 5925 3903 6256
rect 3992 5925 3993 6256
rect 3929 5925 3930 6258
rect 4003 5925 4004 6258
rect 3953 5925 3954 6260
rect 3983 5925 3984 6260
rect 2872 6266 2873 6269
rect 3150 6266 3151 6269
rect 2875 6270 2876 6555
rect 3064 6270 3065 6555
rect 2879 6266 2880 6273
rect 2913 6266 2914 6273
rect 2878 6274 2879 6555
rect 3053 6266 3054 6275
rect 2897 6276 2898 6555
rect 3159 6266 3160 6277
rect 2902 6266 2903 6279
rect 3096 6266 3097 6279
rect 2903 6280 2904 6555
rect 3080 6266 3081 6281
rect 2906 6266 2907 6283
rect 3219 6266 3220 6283
rect 2909 6266 2910 6285
rect 3699 6266 3700 6285
rect 2910 6286 2911 6555
rect 3190 6286 3191 6555
rect 2914 6288 2915 6555
rect 3246 6266 3247 6289
rect 2927 6266 2928 6291
rect 3132 6266 3133 6291
rect 2930 6266 2931 6293
rect 3138 6266 3139 6293
rect 2933 6294 2934 6555
rect 2939 6266 2940 6295
rect 2945 6294 2946 6555
rect 3220 6294 3221 6555
rect 2948 6266 2949 6297
rect 3162 6266 3163 6297
rect 2948 6298 2949 6555
rect 3154 6298 3155 6555
rect 2964 6300 2965 6555
rect 3258 6266 3259 6301
rect 2967 6266 2968 6303
rect 3099 6266 3100 6303
rect 2967 6304 2968 6555
rect 3238 6304 3239 6555
rect 2971 6266 2972 6307
rect 3014 6266 3015 6307
rect 2971 6308 2972 6555
rect 3256 6308 3257 6555
rect 2978 6266 2979 6311
rect 3106 6310 3107 6555
rect 2955 6266 2956 6313
rect 2978 6312 2979 6555
rect 2955 6314 2956 6555
rect 2981 6266 2982 6315
rect 2990 6266 2991 6315
rect 2991 6314 2992 6555
rect 2999 6266 3000 6315
rect 3102 6266 3103 6315
rect 3016 6316 3017 6555
rect 3304 6316 3305 6555
rect 3026 6266 3027 6319
rect 3031 6318 3032 6555
rect 3029 6266 3030 6321
rect 3058 6320 3059 6555
rect 3046 6322 3047 6555
rect 3117 6266 3118 6323
rect 3061 6324 3062 6555
rect 3249 6266 3250 6325
rect 3086 6266 3087 6327
rect 3136 6326 3137 6555
rect 3067 6328 3068 6555
rect 3085 6328 3086 6555
rect 3090 6266 3091 6329
rect 3318 6266 3319 6329
rect 2952 6266 2953 6331
rect 3091 6330 3092 6555
rect 2907 6332 2908 6555
rect 2952 6332 2953 6555
rect 3093 6266 3094 6333
rect 3351 6266 3352 6333
rect 3100 6334 3101 6555
rect 3192 6266 3193 6335
rect 3103 6336 3104 6555
rect 3345 6266 3346 6337
rect 3108 6266 3109 6339
rect 3112 6338 3113 6555
rect 3114 6266 3115 6339
rect 3118 6338 3119 6555
rect 3126 6266 3127 6339
rect 3342 6266 3343 6339
rect 3070 6340 3071 6555
rect 3343 6340 3344 6555
rect 3129 6266 3130 6343
rect 3396 6266 3397 6343
rect 3120 6266 3121 6345
rect 3130 6344 3131 6555
rect 2923 6266 2924 6347
rect 3121 6346 3122 6555
rect 3142 6346 3143 6555
rect 3144 6266 3145 6347
rect 3148 6346 3149 6555
rect 3168 6266 3169 6347
rect 3166 6348 3167 6555
rect 3180 6266 3181 6349
rect 3172 6350 3173 6555
rect 3174 6266 3175 6351
rect 3178 6350 3179 6555
rect 3282 6266 3283 6351
rect 3184 6352 3185 6555
rect 3186 6266 3187 6353
rect 3196 6352 3197 6555
rect 3204 6266 3205 6353
rect 3199 6354 3200 6555
rect 3207 6266 3208 6355
rect 3202 6356 3203 6555
rect 3210 6266 3211 6357
rect 3041 6266 3042 6359
rect 3211 6358 3212 6555
rect 3208 6360 3209 6555
rect 3216 6266 3217 6361
rect 3214 6362 3215 6555
rect 3228 6266 3229 6363
rect 3222 6266 3223 6365
rect 3232 6364 3233 6555
rect 3226 6366 3227 6555
rect 3537 6266 3538 6367
rect 3234 6266 3235 6369
rect 3244 6368 3245 6555
rect 3250 6368 3251 6555
rect 3252 6266 3253 6369
rect 3264 6266 3265 6369
rect 3286 6368 3287 6555
rect 3268 6370 3269 6555
rect 3315 6266 3316 6371
rect 3270 6266 3271 6373
rect 3316 6372 3317 6555
rect 3273 6266 3274 6375
rect 3319 6374 3320 6555
rect 3274 6376 3275 6555
rect 3276 6266 3277 6377
rect 3277 6378 3278 6555
rect 3279 6266 3280 6379
rect 3292 6378 3293 6555
rect 3294 6266 3295 6379
rect 3295 6380 3296 6555
rect 3297 6266 3298 6381
rect 3298 6382 3299 6555
rect 3306 6266 3307 6383
rect 3307 6384 3308 6555
rect 3309 6266 3310 6385
rect 3310 6386 3311 6555
rect 3312 6266 3313 6387
rect 2981 6388 2982 6555
rect 3313 6388 3314 6555
rect 3328 6388 3329 6555
rect 3330 6266 3331 6389
rect 3334 6388 3335 6555
rect 3336 6266 3337 6389
rect 3337 6390 3338 6555
rect 3339 6266 3340 6391
rect 3340 6392 3341 6555
rect 3348 6266 3349 6393
rect 3346 6394 3347 6555
rect 3402 6266 3403 6395
rect 3349 6396 3350 6555
rect 3540 6266 3541 6397
rect 3352 6398 3353 6555
rect 3674 6398 3675 6555
rect 3354 6266 3355 6401
rect 3394 6400 3395 6555
rect 3358 6402 3359 6555
rect 3360 6266 3361 6403
rect 3364 6402 3365 6555
rect 3480 6266 3481 6403
rect 3366 6266 3367 6405
rect 3388 6404 3389 6555
rect 3367 6406 3368 6555
rect 3642 6266 3643 6407
rect 3370 6408 3371 6555
rect 3372 6266 3373 6409
rect 3376 6408 3377 6555
rect 3384 6266 3385 6409
rect 3382 6410 3383 6555
rect 3390 6266 3391 6411
rect 3400 6410 3401 6555
rect 3712 6266 3713 6411
rect 3406 6412 3407 6555
rect 3752 6412 3753 6555
rect 3408 6266 3409 6415
rect 3778 6414 3779 6555
rect 3412 6416 3413 6555
rect 3414 6266 3415 6417
rect 3418 6416 3419 6555
rect 3420 6266 3421 6417
rect 3424 6416 3425 6555
rect 3772 6266 3773 6417
rect 3430 6418 3431 6555
rect 3432 6266 3433 6419
rect 3436 6418 3437 6555
rect 3462 6266 3463 6419
rect 3442 6420 3443 6555
rect 3456 6266 3457 6421
rect 3444 6266 3445 6423
rect 3448 6422 3449 6555
rect 3454 6422 3455 6555
rect 3525 6266 3526 6423
rect 3466 6424 3467 6555
rect 3782 6266 3783 6425
rect 3472 6426 3473 6555
rect 3495 6266 3496 6427
rect 3474 6266 3475 6429
rect 3830 6266 3831 6429
rect 3478 6430 3479 6555
rect 3492 6266 3493 6431
rect 3486 6266 3487 6433
rect 3487 6432 3488 6555
rect 3493 6432 3494 6555
rect 3513 6266 3514 6433
rect 3501 6266 3502 6435
rect 3627 6266 3628 6435
rect 3505 6436 3506 6555
rect 3579 6266 3580 6437
rect 3511 6438 3512 6555
rect 3591 6266 3592 6439
rect 3517 6440 3518 6555
rect 3543 6266 3544 6441
rect 3519 6266 3520 6443
rect 3526 6442 3527 6555
rect 3523 6444 3524 6555
rect 3555 6266 3556 6445
rect 3529 6446 3530 6555
rect 3585 6266 3586 6447
rect 3531 6266 3532 6449
rect 3583 6448 3584 6555
rect 3535 6450 3536 6555
rect 3549 6266 3550 6451
rect 3553 6450 3554 6555
rect 3802 6450 3803 6555
rect 3556 6452 3557 6555
rect 3576 6266 3577 6453
rect 3558 6266 3559 6455
rect 3880 6266 3881 6455
rect 3561 6266 3562 6457
rect 3845 6456 3846 6555
rect 3565 6458 3566 6555
rect 3615 6266 3616 6459
rect 3567 6266 3568 6461
rect 3571 6460 3572 6555
rect 3589 6460 3590 6555
rect 3603 6266 3604 6461
rect 3592 6462 3593 6555
rect 3608 6462 3609 6555
rect 3595 6464 3596 6555
rect 3633 6266 3634 6465
rect 3598 6466 3599 6555
rect 3639 6266 3640 6467
rect 3606 6266 3607 6469
rect 3702 6266 3703 6469
rect 3611 6470 3612 6555
rect 3657 6266 3658 6471
rect 3617 6472 3618 6555
rect 3840 6266 3841 6473
rect 3630 6266 3631 6475
rect 3793 6266 3794 6475
rect 3621 6266 3622 6477
rect 3793 6476 3794 6555
rect 3636 6266 3637 6479
rect 3755 6478 3756 6555
rect 3635 6480 3636 6555
rect 3651 6266 3652 6481
rect 3641 6482 3642 6555
rect 3663 6266 3664 6483
rect 3647 6484 3648 6555
rect 3687 6266 3688 6485
rect 3653 6486 3654 6555
rect 3814 6266 3815 6487
rect 3659 6488 3660 6555
rect 3696 6266 3697 6489
rect 3662 6490 3663 6555
rect 3665 6490 3666 6555
rect 3669 6266 3670 6491
rect 3705 6266 3706 6491
rect 3000 6492 3001 6555
rect 3668 6492 3669 6555
rect 3672 6266 3673 6493
rect 3775 6492 3776 6555
rect 3677 6494 3678 6555
rect 3693 6266 3694 6495
rect 3698 6494 3699 6555
rect 3727 6266 3728 6495
rect 3701 6496 3702 6555
rect 3823 6496 3824 6555
rect 3704 6498 3705 6555
rect 3736 6266 3737 6499
rect 3707 6500 3708 6555
rect 3739 6266 3740 6501
rect 3716 6502 3717 6555
rect 3760 6266 3761 6503
rect 3541 6504 3542 6555
rect 3759 6504 3760 6555
rect 3719 6506 3720 6555
rect 3748 6266 3749 6507
rect 3728 6508 3729 6555
rect 3769 6266 3770 6509
rect 3573 6266 3574 6511
rect 3769 6510 3770 6555
rect 3733 6266 3734 6513
rect 3887 6266 3888 6513
rect 3734 6514 3735 6555
rect 3766 6266 3767 6515
rect 3746 6516 3747 6555
rect 3789 6266 3790 6517
rect 3749 6518 3750 6555
rect 3786 6266 3787 6519
rect 3763 6266 3764 6521
rect 3826 6266 3827 6521
rect 3559 6522 3560 6555
rect 3762 6522 3763 6555
rect 3730 6266 3731 6525
rect 3826 6524 3827 6555
rect 3772 6526 3773 6555
rect 3811 6266 3812 6527
rect 3790 6528 3791 6555
rect 3805 6266 3806 6529
rect 3450 6266 3451 6531
rect 3805 6530 3806 6555
rect 3796 6266 3797 6533
rect 3837 6266 3838 6533
rect 3796 6534 3797 6555
rect 3817 6266 3818 6535
rect 3799 6536 3800 6555
rect 3820 6266 3821 6537
rect 3671 6538 3672 6555
rect 3819 6538 3820 6555
rect 3808 6266 3809 6541
rect 3842 6540 3843 6555
rect 3438 6266 3439 6543
rect 3809 6542 3810 6555
rect 3829 6542 3830 6555
rect 3850 6266 3851 6543
rect 3832 6544 3833 6555
rect 3853 6266 3854 6545
rect 3847 6266 3848 6547
rect 3866 6266 3867 6547
rect 3859 6548 3860 6555
rect 3870 6266 3871 6549
rect 3008 6266 3009 6551
rect 3869 6550 3870 6555
rect 3863 6266 3864 6553
rect 3873 6266 3874 6553
rect 2887 6559 2888 6562
rect 2896 6561 2897 6822
rect 2890 6559 2891 6564
rect 3064 6559 3065 6564
rect 2900 6565 2901 6822
rect 3268 6559 3269 6566
rect 2903 6567 2904 6822
rect 3144 6567 3145 6822
rect 2907 6559 2908 6570
rect 2921 6559 2922 6570
rect 2907 6571 2908 6822
rect 3154 6559 3155 6572
rect 2914 6571 2915 6822
rect 2914 6559 2915 6572
rect 2924 6559 2925 6574
rect 3202 6559 3203 6574
rect 2924 6575 2925 6822
rect 3046 6559 3047 6576
rect 2928 6577 2929 6822
rect 3045 6577 3046 6822
rect 2933 6559 2934 6580
rect 2940 6579 2941 6822
rect 2945 6559 2946 6580
rect 3214 6559 3215 6580
rect 2952 6559 2953 6582
rect 3081 6581 3082 6822
rect 2962 6583 2963 6822
rect 2991 6559 2992 6584
rect 2964 6559 2965 6586
rect 3258 6585 3259 6822
rect 2974 6559 2975 6588
rect 3250 6559 3251 6588
rect 2974 6589 2975 6822
rect 3246 6589 3247 6822
rect 2981 6559 2982 6592
rect 3241 6559 3242 6592
rect 2985 6593 2986 6822
rect 3190 6559 3191 6594
rect 2995 6595 2996 6822
rect 3292 6559 3293 6596
rect 3004 6597 3005 6822
rect 3031 6559 3032 6598
rect 3006 6559 3007 6600
rect 3106 6559 3107 6600
rect 2917 6601 2918 6822
rect 3105 6601 3106 6822
rect 3000 6559 3001 6604
rect 3007 6603 3008 6822
rect 3013 6603 3014 6822
rect 3605 6559 3606 6604
rect 3016 6605 3017 6822
rect 3252 6605 3253 6822
rect 3030 6607 3031 6822
rect 3334 6559 3335 6608
rect 3034 6559 3035 6610
rect 3337 6559 3338 6610
rect 3033 6611 3034 6822
rect 3058 6559 3059 6612
rect 3037 6559 3038 6614
rect 3321 6613 3322 6822
rect 3036 6615 3037 6822
rect 3061 6559 3062 6616
rect 3063 6615 3064 6822
rect 3330 6615 3331 6822
rect 3070 6559 3071 6618
rect 3333 6617 3334 6822
rect 3085 6559 3086 6620
rect 3349 6559 3350 6620
rect 3084 6621 3085 6822
rect 3091 6559 3092 6622
rect 3100 6559 3101 6622
rect 3189 6621 3190 6822
rect 3099 6623 3100 6822
rect 3112 6559 3113 6624
rect 3108 6625 3109 6822
rect 3118 6559 3119 6626
rect 3111 6627 3112 6822
rect 3121 6559 3122 6628
rect 3126 6627 3127 6822
rect 3130 6559 3131 6628
rect 3132 6627 3133 6822
rect 3142 6559 3143 6628
rect 3136 6559 3137 6630
rect 3234 6629 3235 6822
rect 3138 6631 3139 6822
rect 3148 6559 3149 6632
rect 3150 6631 3151 6822
rect 3166 6559 3167 6632
rect 3156 6633 3157 6822
rect 3343 6559 3344 6634
rect 3162 6635 3163 6822
rect 3172 6559 3173 6636
rect 3165 6637 3166 6822
rect 3295 6559 3296 6638
rect 3020 6639 3021 6822
rect 3294 6639 3295 6822
rect 3174 6641 3175 6822
rect 3184 6559 3185 6642
rect 3178 6559 3179 6644
rect 3438 6643 3439 6822
rect 3180 6645 3181 6822
rect 3196 6559 3197 6646
rect 3183 6647 3184 6822
rect 3199 6559 3200 6648
rect 3192 6649 3193 6822
rect 3208 6559 3209 6650
rect 3195 6651 3196 6822
rect 3211 6559 3212 6652
rect 3204 6653 3205 6822
rect 3220 6559 3221 6654
rect 3210 6655 3211 6822
rect 3232 6559 3233 6656
rect 3216 6657 3217 6822
rect 3244 6559 3245 6658
rect 3222 6659 3223 6822
rect 3238 6559 3239 6660
rect 3226 6559 3227 6662
rect 3355 6559 3356 6662
rect 2952 6663 2953 6822
rect 3225 6663 3226 6822
rect 3228 6663 3229 6822
rect 3262 6559 3263 6664
rect 3240 6665 3241 6822
rect 3256 6559 3257 6666
rect 3264 6665 3265 6822
rect 3274 6559 3275 6666
rect 3267 6667 3268 6822
rect 3277 6559 3278 6668
rect 3270 6669 3271 6822
rect 3286 6559 3287 6670
rect 3276 6671 3277 6822
rect 3316 6559 3317 6672
rect 3282 6673 3283 6822
rect 3298 6559 3299 6674
rect 3288 6675 3289 6822
rect 3304 6559 3305 6676
rect 3291 6677 3292 6822
rect 3307 6559 3308 6678
rect 3300 6679 3301 6822
rect 3310 6559 3311 6680
rect 3303 6681 3304 6822
rect 3313 6559 3314 6682
rect 3088 6559 3089 6684
rect 3312 6683 3313 6822
rect 2971 6559 2972 6686
rect 3087 6685 3088 6822
rect 2971 6687 2972 6822
rect 3261 6687 3262 6822
rect 3315 6687 3316 6822
rect 3319 6559 3320 6688
rect 3318 6689 3319 6822
rect 3328 6559 3329 6690
rect 3324 6691 3325 6822
rect 3340 6559 3341 6692
rect 3339 6693 3340 6822
rect 3352 6559 3353 6694
rect 3348 6695 3349 6822
rect 3358 6559 3359 6696
rect 3364 6559 3365 6696
rect 3390 6695 3391 6822
rect 3367 6559 3368 6698
rect 3597 6697 3598 6822
rect 3366 6699 3367 6822
rect 3370 6559 3371 6700
rect 3372 6699 3373 6822
rect 3863 6559 3864 6700
rect 3376 6559 3377 6702
rect 3378 6701 3379 6822
rect 3382 6559 3383 6702
rect 3384 6701 3385 6822
rect 3388 6559 3389 6702
rect 3396 6701 3397 6822
rect 3394 6559 3395 6704
rect 3420 6703 3421 6822
rect 3402 6705 3403 6822
rect 3412 6559 3413 6706
rect 3406 6559 3407 6708
rect 3426 6707 3427 6822
rect 3418 6559 3419 6710
rect 3585 6709 3586 6822
rect 3430 6559 3431 6712
rect 3456 6711 3457 6822
rect 3432 6713 3433 6822
rect 3744 6713 3745 6822
rect 3436 6559 3437 6716
rect 3450 6715 3451 6822
rect 3448 6559 3449 6718
rect 3462 6717 3463 6822
rect 3468 6717 3469 6822
rect 3807 6717 3808 6822
rect 3472 6559 3473 6720
rect 3489 6719 3490 6822
rect 3478 6559 3479 6722
rect 3480 6721 3481 6822
rect 3487 6559 3488 6722
rect 3501 6721 3502 6822
rect 3493 6559 3494 6724
rect 3507 6723 3508 6822
rect 3511 6559 3512 6724
rect 3810 6723 3811 6822
rect 3523 6559 3524 6726
rect 3816 6559 3817 6726
rect 3517 6559 3518 6728
rect 3522 6727 3523 6822
rect 3526 6559 3527 6728
rect 3852 6559 3853 6728
rect 3535 6559 3536 6730
rect 3546 6729 3547 6822
rect 3529 6559 3530 6732
rect 3534 6731 3535 6822
rect 3505 6559 3506 6734
rect 3528 6733 3529 6822
rect 3540 6733 3541 6822
rect 3541 6559 3542 6734
rect 3552 6733 3553 6822
rect 3553 6559 3554 6734
rect 3555 6733 3556 6822
rect 3556 6559 3557 6734
rect 3571 6559 3572 6734
rect 3759 6559 3760 6734
rect 3565 6559 3566 6736
rect 3570 6735 3571 6822
rect 3559 6559 3560 6738
rect 3564 6737 3565 6822
rect 3576 6737 3577 6822
rect 3583 6559 3584 6738
rect 3582 6739 3583 6822
rect 3793 6559 3794 6740
rect 3589 6559 3590 6742
rect 3608 6559 3609 6742
rect 3342 6743 3343 6822
rect 3609 6743 3610 6822
rect 3588 6745 3589 6822
rect 3592 6559 3593 6746
rect 3400 6559 3401 6748
rect 3591 6747 3592 6822
rect 3603 6747 3604 6822
rect 3617 6559 3618 6748
rect 3611 6559 3612 6750
rect 3621 6749 3622 6822
rect 3360 6751 3361 6822
rect 3612 6751 3613 6822
rect 3627 6751 3628 6822
rect 3659 6559 3660 6752
rect 3630 6753 3631 6822
rect 3668 6559 3669 6754
rect 3466 6559 3467 6756
rect 3669 6755 3670 6822
rect 3633 6757 3634 6822
rect 3641 6559 3642 6758
rect 3635 6559 3636 6760
rect 3639 6759 3640 6822
rect 3645 6759 3646 6822
rect 3653 6559 3654 6760
rect 3474 6761 3475 6822
rect 3654 6761 3655 6822
rect 3651 6763 3652 6822
rect 3768 6763 3769 6822
rect 3662 6559 3663 6766
rect 3840 6765 3841 6822
rect 3663 6767 3664 6822
rect 3671 6559 3672 6768
rect 3424 6559 3425 6770
rect 3672 6769 3673 6822
rect 3666 6771 3667 6822
rect 3674 6559 3675 6772
rect 3454 6559 3455 6774
rect 3675 6773 3676 6822
rect 3677 6559 3678 6774
rect 3777 6773 3778 6822
rect 3678 6775 3679 6822
rect 3775 6559 3776 6776
rect 3690 6777 3691 6822
rect 3716 6559 3717 6778
rect 3693 6779 3694 6822
rect 3719 6559 3720 6780
rect 3696 6781 3697 6822
rect 3701 6559 3702 6782
rect 3698 6559 3699 6784
rect 3826 6559 3827 6784
rect 3442 6559 3443 6786
rect 3699 6785 3700 6822
rect 3346 6559 3347 6788
rect 3441 6787 3442 6822
rect 3103 6559 3104 6790
rect 3345 6789 3346 6822
rect 3702 6789 3703 6822
rect 3704 6559 3705 6790
rect 3705 6791 3706 6822
rect 3707 6559 3708 6792
rect 3714 6791 3715 6822
rect 3784 6791 3785 6822
rect 3720 6793 3721 6822
rect 3728 6559 3729 6794
rect 3726 6795 3727 6822
rect 3734 6559 3735 6796
rect 3732 6797 3733 6822
rect 3749 6559 3750 6798
rect 3746 6559 3747 6800
rect 3753 6799 3754 6822
rect 3750 6801 3751 6822
rect 3805 6559 3806 6802
rect 3756 6803 3757 6822
rect 3772 6559 3773 6804
rect 3771 6805 3772 6822
rect 3819 6559 3820 6806
rect 3794 6807 3795 6822
rect 3796 6559 3797 6808
rect 3647 6559 3648 6810
rect 3797 6809 3798 6822
rect 3799 6559 3800 6810
rect 3845 6559 3846 6810
rect 3827 6811 3828 6822
rect 3829 6559 3830 6812
rect 3830 6813 3831 6822
rect 3835 6559 3836 6814
rect 3832 6559 3833 6816
rect 3838 6559 3839 6816
rect 3849 6559 3850 6816
rect 3864 6815 3865 6822
rect 3790 6559 3791 6818
rect 3850 6817 3851 6822
rect 3408 6819 3409 6822
rect 3791 6819 3792 6822
rect 2896 6826 2897 6829
rect 3105 6826 3106 6829
rect 2907 6826 2908 6831
rect 3144 6826 3145 6831
rect 2912 6832 2913 7097
rect 3180 6826 3181 6833
rect 2914 6826 2915 6835
rect 3242 6834 3243 7097
rect 2922 6836 2923 7097
rect 3264 6826 3265 6837
rect 2924 6826 2925 6839
rect 3045 6826 3046 6839
rect 2940 6826 2941 6841
rect 2971 6826 2972 6841
rect 2952 6826 2953 6843
rect 3113 6842 3114 7097
rect 2959 6826 2960 6845
rect 2966 6844 2967 7097
rect 2963 6846 2964 7097
rect 3183 6826 3184 6847
rect 2978 6826 2979 6849
rect 3258 6826 3259 6849
rect 2979 6850 2980 7097
rect 3138 6826 3139 6851
rect 2981 6826 2982 6853
rect 3027 6826 3028 6853
rect 2982 6854 2983 7097
rect 3004 6826 3005 6855
rect 2917 6826 2918 6857
rect 3004 6856 3005 7097
rect 2985 6826 2986 6859
rect 3252 6826 3253 6859
rect 2988 6826 2989 6861
rect 3013 6826 3014 6861
rect 2995 6862 2996 7097
rect 3284 6862 3285 7097
rect 3007 6826 3008 6865
rect 3010 6864 3011 7097
rect 3022 6864 3023 7097
rect 3033 6826 3034 6865
rect 3034 6866 3035 7097
rect 3315 6826 3316 6867
rect 3036 6826 3037 6869
rect 3251 6868 3252 7097
rect 3037 6870 3038 7097
rect 3254 6870 3255 7097
rect 3044 6872 3045 7097
rect 3278 6872 3279 7097
rect 3059 6874 3060 7097
rect 3081 6826 3082 6875
rect 3066 6826 3067 6877
rect 3291 6826 3292 6877
rect 3065 6878 3066 7097
rect 3087 6826 3088 6879
rect 3071 6880 3072 7097
rect 3290 6880 3291 7097
rect 3077 6882 3078 7097
rect 3099 6826 3100 6883
rect 3086 6884 3087 7097
rect 3111 6826 3112 6885
rect 3092 6886 3093 7097
rect 3324 6826 3325 6887
rect 3101 6888 3102 7097
rect 3132 6826 3133 6889
rect 3119 6890 3120 7097
rect 3150 6826 3151 6891
rect 3143 6892 3144 7097
rect 3174 6826 3175 6893
rect 3149 6894 3150 7097
rect 3156 6826 3157 6895
rect 3167 6894 3168 7097
rect 3210 6826 3211 6895
rect 3173 6896 3174 7097
rect 3216 6826 3217 6897
rect 3179 6898 3180 7097
rect 3192 6826 3193 6899
rect 2928 6826 2929 6901
rect 3191 6900 3192 7097
rect 2929 6902 2930 7097
rect 3248 6902 3249 7097
rect 3182 6904 3183 7097
rect 3195 6826 3196 6905
rect 3084 6826 3085 6907
rect 3194 6906 3195 7097
rect 3083 6908 3084 7097
rect 3108 6826 3109 6909
rect 3107 6910 3108 7097
rect 3126 6826 3127 6911
rect 3125 6912 3126 7097
rect 3162 6826 3163 6913
rect 3161 6914 3162 7097
rect 3204 6826 3205 6915
rect 2903 6826 2904 6917
rect 3203 6916 3204 7097
rect 3189 6826 3190 6919
rect 3345 6826 3346 6919
rect 3206 6920 3207 7097
rect 3270 6826 3271 6921
rect 3212 6922 3213 7097
rect 3222 6826 3223 6923
rect 3215 6924 3216 7097
rect 3225 6826 3226 6925
rect 2974 6826 2975 6927
rect 3224 6926 3225 7097
rect 3218 6928 3219 7097
rect 3276 6826 3277 6929
rect 3230 6930 3231 7097
rect 3240 6826 3241 6931
rect 3234 6826 3235 6933
rect 3314 6932 3315 7097
rect 3233 6934 3234 7097
rect 3267 6826 3268 6935
rect 3236 6936 3237 7097
rect 3246 6826 3247 6937
rect 3266 6936 3267 7097
rect 3282 6826 3283 6937
rect 3272 6938 3273 7097
rect 3288 6826 3289 6939
rect 3165 6826 3166 6941
rect 3287 6940 3288 7097
rect 3300 6826 3301 6941
rect 3308 6940 3309 7097
rect 3228 6826 3229 6943
rect 3299 6942 3300 7097
rect 3227 6944 3228 7097
rect 3261 6826 3262 6945
rect 3318 6826 3319 6945
rect 3326 6944 3327 7097
rect 3323 6946 3324 7097
rect 3675 6826 3676 6947
rect 3330 6826 3331 6949
rect 3338 6948 3339 7097
rect 3321 6826 3322 6951
rect 3329 6950 3330 7097
rect 3312 6826 3313 6953
rect 3320 6952 3321 7097
rect 3303 6826 3304 6955
rect 3311 6954 3312 7097
rect 3294 6826 3295 6957
rect 3302 6956 3303 7097
rect 3342 6826 3343 6957
rect 3344 6956 3345 7097
rect 3333 6826 3334 6959
rect 3341 6958 3342 7097
rect 3296 6960 3297 7097
rect 3332 6960 3333 7097
rect 3348 6826 3349 6961
rect 3353 6960 3354 7097
rect 3063 6826 3064 6963
rect 3347 6962 3348 7097
rect 3402 6826 3403 6963
rect 3834 6962 3835 7097
rect 3372 6826 3373 6965
rect 3401 6964 3402 7097
rect 3366 6826 3367 6967
rect 3371 6966 3372 7097
rect 3360 6826 3361 6969
rect 3365 6968 3366 7097
rect 3408 6826 3409 6969
rect 3413 6968 3414 7097
rect 3426 6826 3427 6969
rect 3788 6826 3789 6969
rect 3390 6826 3391 6971
rect 3425 6970 3426 7097
rect 3378 6826 3379 6973
rect 3389 6972 3390 7097
rect 3336 6826 3337 6975
rect 3377 6974 3378 7097
rect 3335 6976 3336 7097
rect 3474 6826 3475 6977
rect 3441 6826 3442 6979
rect 3464 6978 3465 7097
rect 3456 6826 3457 6981
rect 3810 6826 3811 6981
rect 3450 6826 3451 6983
rect 3455 6982 3456 7097
rect 3473 6982 3474 7097
rect 3862 6982 3863 7097
rect 3480 6826 3481 6985
rect 3485 6984 3486 7097
rect 3468 6826 3469 6987
rect 3479 6986 3480 7097
rect 3462 6826 3463 6989
rect 3467 6988 3468 7097
rect 3438 6826 3439 6991
rect 3461 6990 3462 7097
rect 3432 6826 3433 6993
rect 3437 6992 3438 7097
rect 3396 6826 3397 6995
rect 3431 6994 3432 7097
rect 3384 6826 3385 6997
rect 3395 6996 3396 7097
rect 3383 6998 3384 7097
rect 3614 6998 3615 7097
rect 3489 6826 3490 7001
rect 3840 6826 3841 7001
rect 3494 7002 3495 7097
rect 3672 6826 3673 7003
rect 3501 6826 3502 7005
rect 3512 7004 3513 7097
rect 3522 6826 3523 7005
rect 3530 7004 3531 7097
rect 3524 7006 3525 7097
rect 3669 6826 3670 7007
rect 3528 6826 3529 7009
rect 3542 7008 3543 7097
rect 3534 6826 3535 7011
rect 3548 7010 3549 7097
rect 3536 7012 3537 7097
rect 3576 6826 3577 7013
rect 3546 6826 3547 7015
rect 3560 7014 3561 7097
rect 3552 6826 3553 7017
rect 3566 7016 3567 7097
rect 3564 6826 3565 7019
rect 3575 7018 3576 7097
rect 3572 7020 3573 7097
rect 3705 6826 3706 7021
rect 3587 7022 3588 7097
rect 3588 6826 3589 7023
rect 3591 6826 3592 7023
rect 3654 6826 3655 7023
rect 3420 6826 3421 7025
rect 3590 7024 3591 7097
rect 3419 7026 3420 7097
rect 3585 6826 3586 7027
rect 3600 6826 3601 7027
rect 3728 7026 3729 7097
rect 3594 6826 3595 7029
rect 3599 7028 3600 7097
rect 3603 6826 3604 7029
rect 3623 7028 3624 7097
rect 3597 6826 3598 7031
rect 3602 7030 3603 7097
rect 3627 6826 3628 7031
rect 3653 7030 3654 7097
rect 3630 6826 3631 7033
rect 3656 7032 3657 7097
rect 3633 6826 3634 7035
rect 3873 7034 3874 7097
rect 3639 6826 3640 7037
rect 3647 7036 3648 7097
rect 3666 6826 3667 7037
rect 3683 7036 3684 7097
rect 3645 6826 3646 7039
rect 3665 7038 3666 7097
rect 3686 7038 3687 7097
rect 3777 6826 3778 7039
rect 3507 6826 3508 7041
rect 3778 7040 3779 7097
rect 3506 7042 3507 7097
rect 3817 6826 3818 7043
rect 3693 6826 3694 7045
rect 3716 7044 3717 7097
rect 2951 7046 2952 7097
rect 3692 7046 3693 7097
rect 3696 6826 3697 7047
rect 3707 7046 3708 7097
rect 3678 6826 3679 7049
rect 3695 7048 3696 7097
rect 3699 6826 3700 7049
rect 3710 7048 3711 7097
rect 3702 6826 3703 7051
rect 3843 6826 3844 7051
rect 3720 6826 3721 7053
rect 3781 6826 3782 7053
rect 3719 7054 3720 7097
rect 3830 6826 3831 7055
rect 3407 7056 3408 7097
rect 3831 7056 3832 7097
rect 3722 7058 3723 7097
rect 3836 6826 3837 7059
rect 3726 6826 3727 7061
rect 3784 6826 3785 7061
rect 3609 6826 3610 7063
rect 3725 7062 3726 7097
rect 3747 6826 3748 7063
rect 3824 7062 3825 7097
rect 3749 7064 3750 7097
rect 3750 6826 3751 7065
rect 3756 6826 3757 7065
rect 3781 7064 3782 7097
rect 3617 7066 3618 7097
rect 3755 7066 3756 7097
rect 3765 7066 3766 7097
rect 3807 6826 3808 7067
rect 3753 6826 3754 7069
rect 3808 7068 3809 7097
rect 3732 6826 3733 7071
rect 3752 7070 3753 7097
rect 3714 6826 3715 7073
rect 3731 7072 3732 7097
rect 3690 6826 3691 7075
rect 3713 7074 3714 7097
rect 3663 6826 3664 7077
rect 3689 7076 3690 7097
rect 3775 7076 3776 7097
rect 3866 7076 3867 7097
rect 3794 6826 3795 7079
rect 3799 7078 3800 7097
rect 3768 6826 3769 7081
rect 3793 7080 3794 7097
rect 3797 6826 3798 7081
rect 3802 7080 3803 7097
rect 3771 6826 3772 7083
rect 3796 7082 3797 7097
rect 3621 6826 3622 7085
rect 3772 7084 3773 7097
rect 3811 7084 3812 7097
rect 3850 6826 3851 7085
rect 3814 6826 3815 7087
rect 3827 6826 3828 7087
rect 3582 6826 3583 7089
rect 3814 7088 3815 7097
rect 3570 6826 3571 7091
rect 3581 7090 3582 7097
rect 3555 6826 3556 7093
rect 3569 7092 3570 7097
rect 3540 6826 3541 7095
rect 3554 7094 3555 7097
rect 3854 6826 3855 7095
rect 3864 6826 3865 7095
rect 2893 7101 2894 7104
rect 3203 7101 3204 7104
rect 2908 7101 2909 7106
rect 3204 7105 3205 7390
rect 2911 7107 2912 7390
rect 2963 7101 2964 7108
rect 2915 7101 2916 7110
rect 3101 7101 3102 7110
rect 2919 7101 2920 7112
rect 3194 7101 3195 7112
rect 2918 7113 2919 7390
rect 3083 7101 3084 7114
rect 2921 7115 2922 7390
rect 3077 7101 3078 7116
rect 2926 7101 2927 7118
rect 3251 7101 3252 7118
rect 2925 7119 2926 7390
rect 3248 7101 3249 7120
rect 2928 7121 2929 7390
rect 3105 7121 3106 7390
rect 2950 7123 2951 7390
rect 3189 7123 3190 7390
rect 2954 7101 2955 7126
rect 3191 7101 3192 7126
rect 2956 7127 2957 7390
rect 2966 7101 2967 7128
rect 2959 7129 2960 7390
rect 3081 7129 3082 7390
rect 2969 7101 2970 7132
rect 3096 7131 3097 7390
rect 2969 7133 2970 7390
rect 3461 7101 3462 7134
rect 2972 7101 2973 7136
rect 3227 7101 3228 7136
rect 2973 7137 2974 7390
rect 3236 7101 3237 7138
rect 2966 7139 2967 7390
rect 3237 7139 3238 7390
rect 2976 7101 2977 7142
rect 3113 7101 3114 7142
rect 2985 7101 2986 7144
rect 3306 7143 3307 7390
rect 2995 7101 2996 7146
rect 3093 7145 3094 7390
rect 2994 7147 2995 7390
rect 3010 7101 3011 7148
rect 3000 7149 3001 7390
rect 3004 7101 3005 7150
rect 3006 7149 3007 7390
rect 3063 7149 3064 7390
rect 3009 7151 3010 7390
rect 3254 7101 3255 7152
rect 3022 7101 3023 7154
rect 3258 7153 3259 7390
rect 3030 7155 3031 7390
rect 3065 7101 3066 7156
rect 3037 7101 3038 7158
rect 3272 7101 3273 7158
rect 2979 7101 2980 7160
rect 3036 7159 3037 7390
rect 2979 7161 2980 7390
rect 2982 7101 2983 7162
rect 3041 7101 3042 7162
rect 3161 7101 3162 7162
rect 3042 7163 3043 7390
rect 3320 7101 3321 7164
rect 3048 7165 3049 7390
rect 3059 7101 3060 7166
rect 3060 7167 3061 7390
rect 3165 7167 3166 7390
rect 3074 7101 3075 7170
rect 3338 7101 3339 7170
rect 3075 7171 3076 7390
rect 3311 7101 3312 7172
rect 3086 7101 3087 7174
rect 3240 7173 3241 7390
rect 3087 7175 3088 7390
rect 3314 7101 3315 7176
rect 3107 7101 3108 7178
rect 3677 7101 3678 7178
rect 3111 7179 3112 7390
rect 3119 7101 3120 7180
rect 3117 7181 3118 7390
rect 3125 7101 3126 7182
rect 3123 7183 3124 7390
rect 3149 7101 3150 7184
rect 3129 7185 3130 7390
rect 3278 7101 3279 7186
rect 3143 7101 3144 7188
rect 3153 7187 3154 7390
rect 3147 7189 3148 7390
rect 3215 7101 3216 7190
rect 3167 7101 3168 7192
rect 3177 7191 3178 7390
rect 3171 7193 3172 7390
rect 3179 7101 3180 7194
rect 3173 7101 3174 7196
rect 3195 7195 3196 7390
rect 3174 7197 3175 7390
rect 3182 7101 3183 7198
rect 3197 7101 3198 7198
rect 3261 7197 3262 7390
rect 3200 7101 3201 7200
rect 3425 7101 3426 7200
rect 3201 7201 3202 7390
rect 3212 7101 3213 7202
rect 3206 7101 3207 7204
rect 3213 7203 3214 7390
rect 3057 7205 3058 7390
rect 3207 7205 3208 7390
rect 3222 7205 3223 7390
rect 3233 7101 3234 7206
rect 3224 7101 3225 7208
rect 3743 7101 3744 7208
rect 3218 7101 3219 7210
rect 3225 7209 3226 7390
rect 3219 7211 3220 7390
rect 3230 7101 3231 7212
rect 3231 7213 3232 7390
rect 3329 7101 3330 7214
rect 3071 7101 3072 7216
rect 3330 7215 3331 7390
rect 3242 7101 3243 7218
rect 3255 7217 3256 7390
rect 3089 7101 3090 7220
rect 3243 7219 3244 7390
rect 3246 7219 3247 7390
rect 3341 7101 3342 7220
rect 3144 7221 3145 7390
rect 3342 7221 3343 7390
rect 3266 7101 3267 7224
rect 3267 7223 3268 7390
rect 3287 7101 3288 7224
rect 3294 7223 3295 7390
rect 3288 7225 3289 7390
rect 3344 7101 3345 7226
rect 3299 7101 3300 7228
rect 3312 7227 3313 7390
rect 3302 7101 3303 7230
rect 3315 7229 3316 7390
rect 3303 7231 3304 7390
rect 3308 7101 3309 7232
rect 3296 7101 3297 7234
rect 3309 7233 3310 7390
rect 3290 7101 3291 7236
rect 3297 7235 3298 7390
rect 3284 7101 3285 7238
rect 3291 7237 3292 7390
rect 3132 7239 3133 7390
rect 3285 7239 3286 7390
rect 3318 7239 3319 7390
rect 3323 7101 3324 7240
rect 3321 7241 3322 7390
rect 3335 7101 3336 7242
rect 3326 7101 3327 7244
rect 3327 7243 3328 7390
rect 3333 7243 3334 7390
rect 3602 7101 3603 7244
rect 3339 7245 3340 7390
rect 3347 7101 3348 7246
rect 3345 7247 3346 7390
rect 3383 7101 3384 7248
rect 3348 7249 3349 7390
rect 3599 7101 3600 7250
rect 3351 7251 3352 7390
rect 3389 7101 3390 7252
rect 3353 7101 3354 7254
rect 3736 7253 3737 7390
rect 3357 7255 3358 7390
rect 3377 7101 3378 7256
rect 3363 7257 3364 7390
rect 3365 7101 3366 7258
rect 3369 7257 3370 7390
rect 3371 7101 3372 7258
rect 3381 7257 3382 7390
rect 3590 7101 3591 7258
rect 3393 7259 3394 7390
rect 3494 7101 3495 7260
rect 3399 7261 3400 7390
rect 3413 7101 3414 7262
rect 3401 7101 3402 7264
rect 3611 7101 3612 7264
rect 3405 7265 3406 7390
rect 3407 7101 3408 7266
rect 3411 7265 3412 7390
rect 3762 7101 3763 7266
rect 3423 7267 3424 7390
rect 3536 7101 3537 7268
rect 3429 7269 3430 7390
rect 3455 7101 3456 7270
rect 3431 7101 3432 7272
rect 3746 7101 3747 7272
rect 3435 7273 3436 7390
rect 3817 7101 3818 7274
rect 3437 7101 3438 7276
rect 3765 7101 3766 7276
rect 3441 7277 3442 7390
rect 3710 7101 3711 7278
rect 3450 7279 3451 7390
rect 3467 7101 3468 7280
rect 3456 7281 3457 7390
rect 3569 7101 3570 7282
rect 3462 7283 3463 7390
rect 3772 7101 3773 7284
rect 3464 7101 3465 7286
rect 3703 7285 3704 7390
rect 3395 7101 3396 7288
rect 3465 7287 3466 7390
rect 3468 7287 3469 7390
rect 3542 7101 3543 7288
rect 3473 7101 3474 7290
rect 3866 7101 3867 7290
rect 3474 7291 3475 7390
rect 3485 7101 3486 7292
rect 3477 7293 3478 7390
rect 3512 7101 3513 7294
rect 3479 7101 3480 7296
rect 3862 7101 3863 7296
rect 3483 7297 3484 7390
rect 3778 7101 3779 7298
rect 3489 7299 3490 7390
rect 3575 7101 3576 7300
rect 3501 7301 3502 7390
rect 3530 7101 3531 7302
rect 3513 7303 3514 7390
rect 3728 7101 3729 7304
rect 3506 7101 3507 7306
rect 3729 7305 3730 7390
rect 3507 7307 3508 7390
rect 3560 7101 3561 7308
rect 3519 7309 3520 7390
rect 3572 7101 3573 7310
rect 3522 7311 3523 7390
rect 3581 7101 3582 7312
rect 3528 7313 3529 7390
rect 3617 7101 3618 7314
rect 3534 7315 3535 7390
rect 3805 7101 3806 7316
rect 3537 7317 3538 7390
rect 3566 7101 3567 7318
rect 3546 7319 3547 7390
rect 3686 7101 3687 7320
rect 3552 7321 3553 7390
rect 3653 7101 3654 7322
rect 3554 7101 3555 7324
rect 3651 7323 3652 7390
rect 3555 7325 3556 7390
rect 3656 7101 3657 7326
rect 3564 7327 3565 7390
rect 3722 7101 3723 7328
rect 3582 7329 3583 7390
rect 3658 7329 3659 7390
rect 3587 7101 3588 7332
rect 3758 7101 3759 7332
rect 3600 7333 3601 7390
rect 3713 7101 3714 7334
rect 3603 7335 3604 7390
rect 3716 7101 3717 7336
rect 3606 7337 3607 7390
rect 3689 7101 3690 7338
rect 3609 7339 3610 7390
rect 3692 7101 3693 7340
rect 3618 7341 3619 7390
rect 3695 7101 3696 7342
rect 3623 7101 3624 7344
rect 3859 7101 3860 7344
rect 3624 7345 3625 7390
rect 3719 7101 3720 7346
rect 3419 7101 3420 7348
rect 3719 7347 3720 7390
rect 3627 7349 3628 7390
rect 3852 7101 3853 7350
rect 3636 7351 3637 7390
rect 3749 7101 3750 7352
rect 3639 7353 3640 7390
rect 3731 7101 3732 7354
rect 3642 7355 3643 7390
rect 3655 7355 3656 7390
rect 3645 7357 3646 7390
rect 3725 7101 3726 7358
rect 3661 7359 3662 7390
rect 3799 7101 3800 7360
rect 3665 7101 3666 7362
rect 3764 7361 3765 7390
rect 3647 7101 3648 7364
rect 3664 7363 3665 7390
rect 3387 7365 3388 7390
rect 3648 7365 3649 7390
rect 3667 7365 3668 7390
rect 3683 7101 3684 7366
rect 3680 7101 3681 7368
rect 3802 7101 3803 7368
rect 3679 7369 3680 7390
rect 3775 7101 3776 7370
rect 3682 7371 3683 7390
rect 3771 7371 3772 7390
rect 3685 7373 3686 7390
rect 3781 7101 3782 7374
rect 3697 7375 3698 7390
rect 3793 7101 3794 7376
rect 3700 7377 3701 7390
rect 3796 7101 3797 7378
rect 3707 7101 3708 7380
rect 3841 7101 3842 7380
rect 3548 7101 3549 7382
rect 3706 7381 3707 7390
rect 3524 7101 3525 7384
rect 3549 7383 3550 7390
rect 3716 7383 3717 7390
rect 3811 7101 3812 7384
rect 3752 7101 3753 7386
rect 3755 7101 3756 7386
rect 3757 7385 3758 7390
rect 3838 7101 3839 7386
rect 3814 7101 3815 7388
rect 3820 7101 3821 7388
rect 2911 7394 2912 7397
rect 2956 7394 2957 7397
rect 2918 7398 2919 7633
rect 3000 7394 3001 7399
rect 2928 7394 2929 7401
rect 3255 7394 3256 7401
rect 2935 7394 2936 7403
rect 3189 7394 3190 7403
rect 2962 7394 2963 7405
rect 3345 7394 3346 7405
rect 2962 7406 2963 7633
rect 3333 7394 3334 7407
rect 2966 7394 2967 7409
rect 3291 7394 3292 7409
rect 2969 7394 2970 7411
rect 3315 7394 3316 7411
rect 2969 7412 2970 7633
rect 3036 7394 3037 7413
rect 2925 7414 2926 7633
rect 3035 7414 3036 7633
rect 2973 7394 2974 7417
rect 3004 7416 3005 7633
rect 2979 7394 2980 7419
rect 2989 7418 2990 7633
rect 2985 7394 2986 7421
rect 3294 7394 3295 7421
rect 2979 7422 2980 7633
rect 2986 7422 2987 7633
rect 2994 7394 2995 7423
rect 3135 7422 3136 7633
rect 3006 7394 3007 7425
rect 3252 7424 3253 7633
rect 3007 7426 3008 7633
rect 3050 7426 3051 7633
rect 3009 7394 3010 7429
rect 3231 7394 3232 7429
rect 3017 7430 3018 7633
rect 3045 7394 3046 7431
rect 3038 7432 3039 7633
rect 3258 7394 3259 7433
rect 3042 7394 3043 7435
rect 3411 7394 3412 7435
rect 3030 7394 3031 7437
rect 3041 7436 3042 7633
rect 3054 7436 3055 7633
rect 3090 7394 3091 7437
rect 2953 7394 2954 7439
rect 3090 7438 3091 7633
rect 3057 7394 3058 7441
rect 3330 7394 3331 7441
rect 3057 7442 3058 7633
rect 3168 7442 3169 7633
rect 3063 7394 3064 7445
rect 3078 7444 3079 7633
rect 3075 7394 3076 7447
rect 3102 7446 3103 7633
rect 3093 7394 3094 7449
rect 3108 7448 3109 7633
rect 3105 7394 3106 7451
rect 3120 7450 3121 7633
rect 3111 7394 3112 7453
rect 3126 7452 3127 7633
rect 3096 7394 3097 7455
rect 3111 7454 3112 7633
rect 3081 7394 3082 7457
rect 3096 7456 3097 7633
rect 3114 7456 3115 7633
rect 3417 7456 3418 7633
rect 3123 7394 3124 7459
rect 3138 7458 3139 7633
rect 3129 7394 3130 7461
rect 3243 7394 3244 7461
rect 3132 7394 3133 7463
rect 3399 7394 3400 7463
rect 3117 7394 3118 7465
rect 3132 7464 3133 7633
rect 3147 7394 3148 7465
rect 3150 7464 3151 7633
rect 3153 7394 3154 7465
rect 3156 7464 3157 7633
rect 3165 7394 3166 7465
rect 3315 7464 3316 7633
rect 3171 7394 3172 7467
rect 3186 7466 3187 7633
rect 3171 7468 3172 7633
rect 3246 7394 3247 7469
rect 3174 7394 3175 7471
rect 3189 7470 3190 7633
rect 2958 7472 2959 7633
rect 3174 7472 3175 7633
rect 3177 7394 3178 7473
rect 3210 7472 3211 7633
rect 3048 7394 3049 7475
rect 3177 7474 3178 7633
rect 3047 7476 3048 7633
rect 3300 7476 3301 7633
rect 3192 7478 3193 7633
rect 3195 7394 3196 7479
rect 3207 7394 3208 7479
rect 3258 7478 3259 7633
rect 3213 7394 3214 7481
rect 3228 7480 3229 7633
rect 3219 7394 3220 7483
rect 3246 7482 3247 7633
rect 2914 7394 2915 7485
rect 3219 7484 3220 7633
rect 2914 7486 2915 7633
rect 3216 7486 3217 7633
rect 3222 7394 3223 7487
rect 3249 7486 3250 7633
rect 3201 7394 3202 7489
rect 3222 7488 3223 7633
rect 3234 7488 3235 7633
rect 3237 7394 3238 7489
rect 3237 7490 3238 7633
rect 3240 7394 3241 7491
rect 3225 7394 3226 7493
rect 3240 7492 3241 7633
rect 3204 7394 3205 7495
rect 3225 7494 3226 7633
rect 2932 7394 2933 7497
rect 3204 7496 3205 7633
rect 3243 7496 3244 7633
rect 3318 7394 3319 7497
rect 3261 7394 3262 7499
rect 3276 7498 3277 7633
rect 3267 7394 3268 7501
rect 3270 7500 3271 7633
rect 3144 7502 3145 7633
rect 3267 7502 3268 7633
rect 3282 7502 3283 7633
rect 3297 7394 3298 7503
rect 3285 7394 3286 7505
rect 3345 7504 3346 7633
rect 3291 7506 3292 7633
rect 3306 7394 3307 7507
rect 3294 7508 3295 7633
rect 3309 7394 3310 7509
rect 3297 7510 3298 7633
rect 3312 7394 3313 7511
rect 3306 7512 3307 7633
rect 3321 7394 3322 7513
rect 3312 7514 3313 7633
rect 3327 7394 3328 7515
rect 3318 7516 3319 7633
rect 3330 7516 3331 7633
rect 3342 7394 3343 7517
rect 3360 7516 3361 7633
rect 3288 7394 3289 7519
rect 3342 7518 3343 7633
rect 3288 7520 3289 7633
rect 3303 7394 3304 7521
rect 3348 7394 3349 7521
rect 3384 7520 3385 7633
rect 3348 7522 3349 7633
rect 3363 7394 3364 7523
rect 3339 7394 3340 7525
rect 3363 7524 3364 7633
rect 3351 7394 3352 7527
rect 3372 7526 3373 7633
rect 3354 7528 3355 7633
rect 3357 7394 3358 7529
rect 3369 7394 3370 7529
rect 3736 7394 3737 7529
rect 3387 7394 3388 7531
rect 3414 7530 3415 7633
rect 3381 7394 3382 7533
rect 3387 7532 3388 7633
rect 3390 7532 3391 7633
rect 3405 7394 3406 7533
rect 3393 7394 3394 7535
rect 3408 7534 3409 7633
rect 3396 7536 3397 7633
rect 3558 7536 3559 7633
rect 3399 7538 3400 7633
rect 3465 7394 3466 7539
rect 3402 7540 3403 7633
rect 3719 7394 3720 7541
rect 3420 7542 3421 7633
rect 3549 7394 3550 7543
rect 3426 7544 3427 7633
rect 3441 7394 3442 7545
rect 3435 7394 3436 7547
rect 3441 7546 3442 7633
rect 3429 7394 3430 7549
rect 3435 7548 3436 7633
rect 3423 7394 3424 7551
rect 3429 7550 3430 7633
rect 3447 7550 3448 7633
rect 3456 7394 3457 7551
rect 3453 7552 3454 7633
rect 3468 7394 3469 7553
rect 3459 7554 3460 7633
rect 3474 7394 3475 7555
rect 3462 7394 3463 7557
rect 3561 7394 3562 7557
rect 3462 7558 3463 7633
rect 3710 7394 3711 7559
rect 3468 7560 3469 7633
rect 3528 7394 3529 7561
rect 3477 7394 3478 7563
rect 3480 7562 3481 7633
rect 3483 7394 3484 7563
rect 3486 7562 3487 7633
rect 3489 7394 3490 7563
rect 3648 7394 3649 7563
rect 3501 7562 3502 7633
rect 3501 7394 3502 7563
rect 3510 7564 3511 7633
rect 3704 7564 3705 7633
rect 3513 7394 3514 7567
rect 3622 7566 3623 7633
rect 3525 7568 3526 7633
rect 3534 7394 3535 7569
rect 3528 7570 3529 7633
rect 3537 7394 3538 7571
rect 3537 7572 3538 7633
rect 3629 7572 3630 7633
rect 3540 7574 3541 7633
rect 3546 7394 3547 7575
rect 3543 7576 3544 7633
rect 3552 7394 3553 7577
rect 3546 7578 3547 7633
rect 3555 7394 3556 7579
rect 3561 7578 3562 7633
rect 3664 7394 3665 7579
rect 3573 7580 3574 7633
rect 3582 7394 3583 7581
rect 3579 7582 3580 7633
rect 3600 7394 3601 7583
rect 3582 7584 3583 7633
rect 3603 7394 3604 7585
rect 3564 7394 3565 7587
rect 3603 7586 3604 7633
rect 3507 7394 3508 7589
rect 3564 7588 3565 7633
rect 3507 7590 3508 7633
rect 3519 7394 3520 7591
rect 3585 7590 3586 7633
rect 3609 7394 3610 7591
rect 3594 7592 3595 7633
rect 3618 7394 3619 7593
rect 3576 7594 3577 7633
rect 3619 7594 3620 7633
rect 3600 7596 3601 7633
rect 3624 7394 3625 7597
rect 3606 7394 3607 7599
rect 3781 7394 3782 7599
rect 3606 7600 3607 7633
rect 3639 7394 3640 7601
rect 3450 7394 3451 7603
rect 3640 7602 3641 7633
rect 3609 7604 3610 7633
rect 3729 7394 3730 7605
rect 3612 7606 3613 7633
rect 3661 7394 3662 7607
rect 3627 7394 3628 7609
rect 3725 7394 3726 7609
rect 3633 7610 3634 7633
rect 3636 7394 3637 7611
rect 3642 7394 3643 7611
rect 3658 7394 3659 7611
rect 3645 7394 3646 7613
rect 3655 7394 3656 7613
rect 3643 7614 3644 7633
rect 3655 7614 3656 7633
rect 3652 7616 3653 7633
rect 3716 7394 3717 7617
rect 3658 7618 3659 7633
rect 3685 7394 3686 7619
rect 3670 7394 3671 7621
rect 3722 7394 3723 7621
rect 3522 7394 3523 7623
rect 3721 7622 3722 7633
rect 3670 7624 3671 7633
rect 3697 7394 3698 7625
rect 3673 7626 3674 7633
rect 3700 7394 3701 7627
rect 3679 7394 3680 7629
rect 3774 7394 3775 7629
rect 3321 7630 3322 7633
rect 3679 7630 3680 7633
rect 3682 7394 3683 7631
rect 3727 7630 3728 7633
rect 3743 7394 3744 7631
rect 3760 7394 3761 7631
rect 2809 7637 2810 7640
rect 3447 7637 3448 7640
rect 2888 7641 2889 7850
rect 2894 7641 2895 7850
rect 2924 7641 2925 7850
rect 3060 7641 3061 7850
rect 2928 7637 2929 7644
rect 3038 7637 3039 7644
rect 2931 7645 2932 7850
rect 3219 7637 3220 7646
rect 2964 7647 2965 7850
rect 3273 7647 3274 7850
rect 2967 7649 2968 7850
rect 3246 7637 3247 7650
rect 2969 7637 2970 7652
rect 3041 7637 3042 7652
rect 2972 7637 2973 7654
rect 3017 7637 3018 7654
rect 2986 7637 2987 7656
rect 3321 7655 3322 7850
rect 2989 7637 2990 7658
rect 3013 7657 3014 7850
rect 3035 7637 3036 7658
rect 3063 7657 3064 7850
rect 3039 7659 3040 7850
rect 3405 7659 3406 7850
rect 3050 7637 3051 7662
rect 3276 7637 3277 7662
rect 3057 7637 3058 7664
rect 3144 7637 3145 7664
rect 2960 7665 2961 7850
rect 3144 7665 3145 7850
rect 3072 7667 3073 7850
rect 3078 7637 3079 7668
rect 3078 7669 3079 7850
rect 3114 7637 3115 7670
rect 3084 7671 3085 7850
rect 3102 7637 3103 7672
rect 3090 7671 3091 7850
rect 3090 7637 3091 7672
rect 3096 7671 3097 7850
rect 3096 7637 3097 7672
rect 3102 7673 3103 7850
rect 3108 7637 3109 7674
rect 3105 7675 3106 7850
rect 3111 7637 3112 7676
rect 3108 7677 3109 7850
rect 3138 7637 3139 7678
rect 3114 7679 3115 7850
rect 3132 7637 3133 7680
rect 3117 7681 3118 7850
rect 3135 7637 3136 7682
rect 3120 7637 3121 7684
rect 3138 7683 3139 7850
rect 3123 7685 3124 7850
rect 3351 7685 3352 7850
rect 3129 7687 3130 7850
rect 3171 7637 3172 7688
rect 3156 7637 3157 7690
rect 3180 7689 3181 7850
rect 2957 7691 2958 7850
rect 3156 7691 3157 7850
rect 3165 7691 3166 7850
rect 3363 7637 3364 7692
rect 3174 7637 3175 7694
rect 3198 7693 3199 7850
rect 3177 7637 3178 7696
rect 3201 7695 3202 7850
rect 3189 7637 3190 7698
rect 3213 7697 3214 7850
rect 3204 7637 3205 7700
rect 3318 7637 3319 7700
rect 3216 7637 3217 7702
rect 3264 7701 3265 7850
rect 3192 7637 3193 7704
rect 3216 7703 3217 7850
rect 3219 7703 3220 7850
rect 3249 7637 3250 7704
rect 3222 7637 3223 7706
rect 3246 7705 3247 7850
rect 3210 7637 3211 7708
rect 3222 7707 3223 7850
rect 3186 7637 3187 7710
rect 3210 7709 3211 7850
rect 3225 7637 3226 7710
rect 3249 7709 3250 7850
rect 3228 7709 3229 7850
rect 3228 7637 3229 7710
rect 3234 7637 3235 7712
rect 3285 7711 3286 7850
rect 3234 7713 3235 7850
rect 3240 7637 3241 7714
rect 3029 7715 3030 7850
rect 3240 7715 3241 7850
rect 3252 7637 3253 7716
rect 3267 7715 3268 7850
rect 3252 7717 3253 7850
rect 3258 7637 3259 7718
rect 3270 7637 3271 7718
rect 3309 7717 3310 7850
rect 3282 7637 3283 7720
rect 3333 7719 3334 7850
rect 3288 7637 3289 7722
rect 3357 7721 3358 7850
rect 2921 7637 2922 7724
rect 3288 7723 3289 7850
rect 2920 7725 2921 7850
rect 3016 7725 3017 7850
rect 3294 7637 3295 7726
rect 3339 7725 3340 7850
rect 3300 7637 3301 7728
rect 3303 7727 3304 7850
rect 3312 7637 3313 7728
rect 3363 7727 3364 7850
rect 3327 7729 3328 7850
rect 3345 7637 3346 7730
rect 3306 7637 3307 7732
rect 3345 7731 3346 7850
rect 3330 7637 3331 7734
rect 3381 7733 3382 7850
rect 3348 7637 3349 7736
rect 3423 7735 3424 7850
rect 3369 7737 3370 7850
rect 3468 7637 3469 7738
rect 3372 7637 3373 7740
rect 3393 7739 3394 7850
rect 3375 7741 3376 7850
rect 3387 7637 3388 7742
rect 3032 7743 3033 7850
rect 3387 7743 3388 7850
rect 3390 7637 3391 7744
rect 3465 7743 3466 7850
rect 3315 7637 3316 7746
rect 3390 7745 3391 7850
rect 3399 7637 3400 7746
rect 3417 7745 3418 7850
rect 3354 7637 3355 7748
rect 3399 7747 3400 7850
rect 3342 7637 3343 7750
rect 3354 7749 3355 7850
rect 3297 7637 3298 7752
rect 3342 7751 3343 7850
rect 3297 7753 3298 7850
rect 3429 7637 3430 7754
rect 3402 7637 3403 7756
rect 3471 7755 3472 7850
rect 3411 7757 3412 7850
rect 3414 7637 3415 7758
rect 3384 7637 3385 7760
rect 3414 7759 3415 7850
rect 3420 7637 3421 7760
rect 3721 7637 3722 7760
rect 3396 7637 3397 7762
rect 3420 7761 3421 7850
rect 3426 7637 3427 7762
rect 3495 7761 3496 7850
rect 3426 7763 3427 7850
rect 3546 7637 3547 7764
rect 3429 7765 3430 7850
rect 3462 7637 3463 7766
rect 3435 7637 3436 7768
rect 3665 7767 3666 7850
rect 3435 7769 3436 7850
rect 3453 7637 3454 7770
rect 3441 7637 3442 7772
rect 3477 7771 3478 7850
rect 3162 7773 3163 7850
rect 3441 7773 3442 7850
rect 3447 7773 3448 7850
rect 3650 7773 3651 7850
rect 3459 7637 3460 7776
rect 3522 7775 3523 7850
rect 3459 7777 3460 7850
rect 3640 7637 3641 7778
rect 3453 7779 3454 7850
rect 3639 7779 3640 7850
rect 3486 7637 3487 7782
rect 3633 7781 3634 7850
rect 3504 7783 3505 7850
rect 3712 7783 3713 7850
rect 3510 7637 3511 7786
rect 3700 7637 3701 7786
rect 3150 7637 3151 7788
rect 3510 7787 3511 7850
rect 3126 7637 3127 7790
rect 3150 7789 3151 7850
rect 3126 7791 3127 7850
rect 3168 7637 3169 7792
rect 3516 7791 3517 7850
rect 3707 7637 3708 7792
rect 3525 7637 3526 7794
rect 3552 7793 3553 7850
rect 3480 7637 3481 7796
rect 3525 7795 3526 7850
rect 3528 7637 3529 7796
rect 3555 7795 3556 7850
rect 3537 7637 3538 7798
rect 3567 7797 3568 7850
rect 3507 7637 3508 7800
rect 3537 7799 3538 7850
rect 3540 7637 3541 7800
rect 3619 7637 3620 7800
rect 3501 7637 3502 7802
rect 3540 7801 3541 7850
rect 3543 7637 3544 7802
rect 3597 7801 3598 7850
rect 3561 7637 3562 7804
rect 3588 7803 3589 7850
rect 3564 7637 3565 7806
rect 3591 7805 3592 7850
rect 3564 7807 3565 7850
rect 3629 7637 3630 7808
rect 3570 7809 3571 7850
rect 3573 7637 3574 7810
rect 3573 7811 3574 7850
rect 3576 7637 3577 7812
rect 3579 7637 3580 7812
rect 3695 7811 3696 7850
rect 3582 7637 3583 7814
rect 3662 7813 3663 7850
rect 3585 7637 3586 7816
rect 3727 7637 3728 7816
rect 3594 7637 3595 7818
rect 3618 7817 3619 7850
rect 3237 7637 3238 7820
rect 3594 7819 3595 7850
rect 3237 7821 3238 7850
rect 3243 7637 3244 7822
rect 3600 7637 3601 7822
rect 3624 7821 3625 7850
rect 3600 7823 3601 7850
rect 3609 7637 3610 7824
rect 3603 7637 3604 7826
rect 3627 7825 3628 7850
rect 3606 7637 3607 7828
rect 3615 7827 3616 7850
rect 3612 7829 3613 7850
rect 3636 7637 3637 7830
rect 3630 7831 3631 7850
rect 3730 7831 3731 7850
rect 3655 7637 3656 7834
rect 3702 7833 3703 7850
rect 3656 7835 3657 7850
rect 3733 7835 3734 7850
rect 3670 7637 3671 7838
rect 3689 7837 3690 7850
rect 3652 7637 3653 7840
rect 3671 7839 3672 7850
rect 3673 7637 3674 7840
rect 3692 7839 3693 7850
rect 3674 7841 3675 7850
rect 3686 7637 3687 7842
rect 3676 7637 3677 7844
rect 3705 7843 3706 7850
rect 3658 7637 3659 7846
rect 3677 7845 3678 7850
rect 3659 7847 3660 7850
rect 3679 7637 3680 7848
rect 2884 7854 2885 7857
rect 2894 7854 2895 7857
rect 2888 7854 2889 7859
rect 2917 7854 2918 7859
rect 2914 7860 2915 8097
rect 3063 7854 3064 7861
rect 2918 7862 2919 8097
rect 3285 7854 3286 7863
rect 2921 7864 2922 8097
rect 3198 7854 3199 7865
rect 2931 7854 2932 7867
rect 3006 7866 3007 8097
rect 2946 7854 2947 7869
rect 3288 7854 3289 7869
rect 2960 7854 2961 7871
rect 3138 7854 3139 7871
rect 2961 7872 2962 8097
rect 3108 7854 3109 7873
rect 2965 7874 2966 8097
rect 3267 7854 3268 7875
rect 2967 7854 2968 7877
rect 3234 7854 3235 7877
rect 2968 7878 2969 8097
rect 3129 7854 3130 7879
rect 2975 7880 2976 8097
rect 3136 7880 3137 8097
rect 2995 7854 2996 7883
rect 3213 7854 3214 7883
rect 2943 7854 2944 7885
rect 2994 7884 2995 8097
rect 2997 7884 2998 8097
rect 3013 7854 3014 7885
rect 3003 7886 3004 8097
rect 3345 7854 3346 7887
rect 3018 7888 3019 8097
rect 3390 7854 3391 7889
rect 3022 7854 3023 7891
rect 3156 7854 3157 7891
rect 3025 7892 3026 8097
rect 3268 7892 3269 8097
rect 3029 7854 3030 7895
rect 3385 7894 3386 8097
rect 3032 7854 3033 7897
rect 3331 7896 3332 8097
rect 3016 7854 3017 7899
rect 3031 7898 3032 8097
rect 3037 7898 3038 8097
rect 3540 7854 3541 7899
rect 3046 7900 3047 8097
rect 3391 7900 3392 8097
rect 3049 7902 3050 8097
rect 3235 7902 3236 8097
rect 3058 7904 3059 8097
rect 3078 7854 3079 7905
rect 3060 7854 3061 7907
rect 3064 7906 3065 8097
rect 3072 7854 3073 7907
rect 3073 7906 3074 8097
rect 3102 7854 3103 7907
rect 3103 7906 3104 8097
rect 3105 7854 3106 7907
rect 3106 7906 3107 8097
rect 3112 7906 3113 8097
rect 3399 7854 3400 7907
rect 3114 7854 3115 7909
rect 3115 7908 3116 8097
rect 3117 7854 3118 7909
rect 3118 7908 3119 8097
rect 3120 7854 3121 7909
rect 3327 7854 3328 7909
rect 3121 7910 3122 8097
rect 3144 7854 3145 7911
rect 3126 7854 3127 7913
rect 3133 7912 3134 8097
rect 3127 7914 3128 8097
rect 3150 7854 3151 7915
rect 3139 7916 3140 8097
rect 3643 7854 3644 7917
rect 3145 7918 3146 8097
rect 3180 7854 3181 7919
rect 3157 7920 3158 8097
rect 3210 7854 3211 7921
rect 3165 7854 3166 7923
rect 3303 7854 3304 7923
rect 3172 7924 3173 8097
rect 3216 7854 3217 7925
rect 3175 7926 3176 8097
rect 3219 7854 3220 7927
rect 3184 7928 3185 8097
rect 3240 7854 3241 7929
rect 3186 7854 3187 7931
rect 3367 7930 3368 8097
rect 3189 7854 3190 7933
rect 3375 7854 3376 7933
rect 3190 7934 3191 8097
rect 3246 7854 3247 7935
rect 3193 7936 3194 8097
rect 3249 7854 3250 7937
rect 3196 7938 3197 8097
rect 3222 7854 3223 7939
rect 3201 7854 3202 7941
rect 3484 7940 3485 8097
rect 3202 7942 3203 8097
rect 3228 7854 3229 7943
rect 3205 7944 3206 8097
rect 3237 7854 3238 7945
rect 3208 7946 3209 8097
rect 3264 7854 3265 7947
rect 3211 7948 3212 8097
rect 3273 7854 3274 7949
rect 3241 7950 3242 8097
rect 3426 7854 3427 7951
rect 3247 7952 3248 8097
rect 3309 7854 3310 7953
rect 3259 7954 3260 8097
rect 3420 7854 3421 7955
rect 3265 7956 3266 8097
rect 3351 7854 3352 7957
rect 3271 7958 3272 8097
rect 3333 7854 3334 7959
rect 3277 7960 3278 8097
rect 3297 7854 3298 7961
rect 3283 7962 3284 8097
rect 3339 7854 3340 7963
rect 3252 7854 3253 7965
rect 3340 7964 3341 8097
rect 3253 7966 3254 8097
rect 3354 7854 3355 7967
rect 3286 7968 3287 8097
rect 3342 7854 3343 7969
rect 3289 7970 3290 8097
rect 3321 7854 3322 7971
rect 3291 7854 3292 7973
rect 3646 7854 3647 7973
rect 3295 7974 3296 8097
rect 3393 7854 3394 7975
rect 3301 7976 3302 8097
rect 3357 7854 3358 7977
rect 3304 7978 3305 8097
rect 3360 7854 3361 7979
rect 3307 7980 3308 8097
rect 3363 7854 3364 7981
rect 3313 7982 3314 8097
rect 3417 7854 3418 7983
rect 3319 7984 3320 8097
rect 3381 7854 3382 7985
rect 3325 7986 3326 8097
rect 3487 7986 3488 8097
rect 3337 7988 3338 8097
rect 3387 7854 3388 7989
rect 3343 7990 3344 8097
rect 3369 7854 3370 7991
rect 3349 7992 3350 8097
rect 3535 7992 3536 8097
rect 3355 7994 3356 8097
rect 3405 7854 3406 7995
rect 3358 7996 3359 8097
rect 3408 7854 3409 7997
rect 3361 7998 3362 8097
rect 3411 7854 3412 7999
rect 3364 8000 3365 8097
rect 3414 7854 3415 8001
rect 3373 8002 3374 8097
rect 3423 7854 3424 8003
rect 3388 8004 3389 8097
rect 3441 7854 3442 8005
rect 3397 8006 3398 8097
rect 3453 7854 3454 8007
rect 3403 8008 3404 8097
rect 3459 7854 3460 8009
rect 3415 8010 3416 8097
rect 3465 7854 3466 8011
rect 3429 7854 3430 8013
rect 3653 7854 3654 8013
rect 3433 8014 3434 8097
rect 3552 7854 3553 8015
rect 3316 8016 3317 8097
rect 3552 8016 3553 8097
rect 3435 7854 3436 8019
rect 3650 7854 3651 8019
rect 3436 8020 3437 8097
rect 3555 7854 3556 8021
rect 3439 8022 3440 8097
rect 3504 7854 3505 8023
rect 3447 7854 3448 8025
rect 3639 7854 3640 8025
rect 3451 8026 3452 8097
rect 3537 7854 3538 8027
rect 3454 8028 3455 8097
rect 3674 7854 3675 8029
rect 3457 8030 3458 8097
rect 3471 7854 3472 8031
rect 3460 8032 3461 8097
rect 3594 7854 3595 8033
rect 3463 8034 3464 8097
rect 3597 7854 3598 8035
rect 3466 8036 3467 8097
rect 3525 7854 3526 8037
rect 3472 8038 3473 8097
rect 3522 7854 3523 8039
rect 3475 8040 3476 8097
rect 3633 7854 3634 8041
rect 3477 7854 3478 8043
rect 3668 7854 3669 8043
rect 3478 8044 3479 8097
rect 3570 7854 3571 8045
rect 3481 8046 3482 8097
rect 3573 7854 3574 8047
rect 3490 8048 3491 8097
rect 3642 8048 3643 8097
rect 3493 8050 3494 8097
rect 3600 7854 3601 8051
rect 3495 7854 3496 8053
rect 3572 8052 3573 8097
rect 3499 8054 3500 8097
rect 3627 7854 3628 8055
rect 3502 8056 3503 8097
rect 3603 8056 3604 8097
rect 3514 8058 3515 8097
rect 3665 7854 3666 8059
rect 3516 7854 3517 8061
rect 3733 7854 3734 8061
rect 3517 8062 3518 8097
rect 3588 7854 3589 8063
rect 3520 8064 3521 8097
rect 3662 7854 3663 8065
rect 3529 8066 3530 8097
rect 3612 7854 3613 8067
rect 3532 8068 3533 8097
rect 3615 7854 3616 8069
rect 3545 8070 3546 8097
rect 3567 7854 3568 8071
rect 3549 8072 3550 8097
rect 3659 7854 3660 8073
rect 3564 7854 3565 8075
rect 3600 8074 3601 8097
rect 3575 8076 3576 8097
rect 3677 7854 3678 8077
rect 3587 8078 3588 8097
rect 3689 7854 3690 8079
rect 3591 7854 3592 8081
rect 3712 7854 3713 8081
rect 3590 8082 3591 8097
rect 3692 7854 3693 8083
rect 3618 7854 3619 8085
rect 3740 7854 3741 8085
rect 3569 8086 3570 8097
rect 3617 8086 3618 8097
rect 3624 7854 3625 8087
rect 3716 7854 3717 8087
rect 3630 7854 3631 8089
rect 3747 7854 3748 8089
rect 3645 8090 3646 8097
rect 3666 8090 3667 8097
rect 3656 7854 3657 8093
rect 3754 7854 3755 8093
rect 3671 7854 3672 8095
rect 3705 7854 3706 8095
rect 3760 7854 3761 8095
rect 3764 7854 3765 8095
rect 2921 8101 2922 8104
rect 3208 8101 3209 8104
rect 2918 8101 2919 8106
rect 2920 8105 2921 8316
rect 2927 8105 2928 8316
rect 3304 8101 3305 8106
rect 2932 8101 2933 8108
rect 3085 8101 3086 8108
rect 2931 8109 2932 8316
rect 3145 8101 3146 8110
rect 2935 8101 2936 8112
rect 3091 8101 3092 8112
rect 2954 8101 2955 8114
rect 3103 8101 3104 8114
rect 2965 8101 2966 8116
rect 3227 8115 3228 8316
rect 2975 8101 2976 8118
rect 3106 8101 3107 8118
rect 2975 8119 2976 8316
rect 2997 8101 2998 8120
rect 2987 8101 2988 8122
rect 3271 8101 3272 8122
rect 2991 8101 2992 8124
rect 3046 8101 3047 8124
rect 2990 8125 2991 8316
rect 3283 8101 3284 8126
rect 2993 8127 2994 8316
rect 3340 8101 3341 8128
rect 3003 8129 3004 8316
rect 3006 8101 3007 8130
rect 3018 8101 3019 8130
rect 3319 8101 3320 8130
rect 3018 8131 3019 8316
rect 3307 8101 3308 8132
rect 3025 8101 3026 8134
rect 3263 8133 3264 8316
rect 3027 8135 3028 8316
rect 3188 8135 3189 8316
rect 3034 8137 3035 8316
rect 3235 8101 3236 8138
rect 3041 8139 3042 8316
rect 3218 8139 3219 8316
rect 3049 8101 3050 8142
rect 3200 8141 3201 8316
rect 3056 8143 3057 8316
rect 3058 8101 3059 8144
rect 3062 8143 3063 8316
rect 3064 8101 3065 8144
rect 2925 8101 2926 8146
rect 3065 8145 3066 8316
rect 3068 8145 3069 8316
rect 3139 8101 3140 8146
rect 2961 8101 2962 8148
rect 3140 8147 3141 8316
rect 3073 8101 3074 8150
rect 3074 8149 3075 8316
rect 3077 8149 3078 8316
rect 3133 8101 3134 8150
rect 3080 8151 3081 8316
rect 3136 8101 3137 8152
rect 3095 8153 3096 8316
rect 3115 8101 3116 8154
rect 3097 8101 3098 8156
rect 3245 8155 3246 8316
rect 3098 8157 3099 8316
rect 3118 8101 3119 8158
rect 3101 8159 3102 8316
rect 3121 8101 3122 8160
rect 3119 8161 3120 8316
rect 3205 8101 3206 8162
rect 3127 8101 3128 8164
rect 3538 8101 3539 8164
rect 3131 8165 3132 8316
rect 3157 8101 3158 8166
rect 3134 8167 3135 8316
rect 3172 8101 3173 8168
rect 3021 8101 3022 8170
rect 3173 8169 3174 8316
rect 3021 8171 3022 8316
rect 3031 8101 3032 8172
rect 3031 8173 3032 8316
rect 3265 8101 3266 8174
rect 3143 8175 3144 8316
rect 3175 8101 3176 8176
rect 3152 8177 3153 8316
rect 3196 8101 3197 8178
rect 3158 8179 3159 8316
rect 3184 8101 3185 8180
rect 3164 8181 3165 8316
rect 3190 8101 3191 8182
rect 3167 8183 3168 8316
rect 3193 8101 3194 8184
rect 3170 8185 3171 8316
rect 3202 8101 3203 8186
rect 3182 8187 3183 8316
rect 3211 8101 3212 8188
rect 3194 8189 3195 8316
rect 3268 8101 3269 8190
rect 3212 8191 3213 8316
rect 3247 8101 3248 8192
rect 3215 8193 3216 8316
rect 3286 8101 3287 8194
rect 3224 8195 3225 8316
rect 3253 8101 3254 8196
rect 3230 8197 3231 8316
rect 3259 8101 3260 8198
rect 3236 8199 3237 8316
rect 3277 8101 3278 8200
rect 3241 8101 3242 8202
rect 3413 8201 3414 8316
rect 3242 8203 3243 8316
rect 3301 8101 3302 8204
rect 3248 8205 3249 8316
rect 3289 8101 3290 8206
rect 3254 8207 3255 8316
rect 3295 8101 3296 8208
rect 3260 8209 3261 8316
rect 3313 8101 3314 8210
rect 3266 8211 3267 8316
rect 3325 8101 3326 8212
rect 3272 8213 3273 8316
rect 3337 8101 3338 8214
rect 3275 8215 3276 8316
rect 3535 8101 3536 8216
rect 3281 8217 3282 8316
rect 3367 8101 3368 8218
rect 3287 8219 3288 8316
rect 3355 8101 3356 8220
rect 3290 8221 3291 8316
rect 3358 8101 3359 8222
rect 3293 8223 3294 8316
rect 3361 8101 3362 8224
rect 3296 8225 3297 8316
rect 3364 8101 3365 8226
rect 3299 8227 3300 8316
rect 3373 8101 3374 8228
rect 3311 8229 3312 8316
rect 3391 8101 3392 8230
rect 3316 8101 3317 8232
rect 3419 8231 3420 8316
rect 3317 8233 3318 8316
rect 3385 8101 3386 8234
rect 3320 8235 3321 8316
rect 3388 8101 3389 8236
rect 3323 8237 3324 8316
rect 3397 8101 3398 8238
rect 3329 8239 3330 8316
rect 3403 8101 3404 8240
rect 3089 8241 3090 8316
rect 3404 8241 3405 8316
rect 3341 8243 3342 8316
rect 3470 8243 3471 8316
rect 3349 8101 3350 8246
rect 3559 8101 3560 8246
rect 3359 8247 3360 8316
rect 3433 8101 3434 8248
rect 3362 8249 3363 8316
rect 3436 8101 3437 8250
rect 3365 8251 3366 8316
rect 3439 8101 3440 8252
rect 3377 8253 3378 8316
rect 3451 8101 3452 8254
rect 3386 8255 3387 8316
rect 3454 8101 3455 8256
rect 3389 8257 3390 8316
rect 3457 8101 3458 8258
rect 3343 8101 3344 8260
rect 3458 8259 3459 8316
rect 3392 8261 3393 8316
rect 3466 8101 3467 8262
rect 3331 8101 3332 8264
rect 3467 8263 3468 8316
rect 3398 8265 3399 8316
rect 3472 8101 3473 8266
rect 3401 8267 3402 8316
rect 3475 8101 3476 8268
rect 3410 8269 3411 8316
rect 3460 8101 3461 8270
rect 3415 8101 3416 8272
rect 3522 8271 3523 8316
rect 3422 8273 3423 8316
rect 3532 8101 3533 8274
rect 3425 8275 3426 8316
rect 3499 8101 3500 8276
rect 3428 8277 3429 8316
rect 3555 8277 3556 8316
rect 3437 8279 3438 8316
rect 3514 8101 3515 8280
rect 3440 8281 3441 8316
rect 3502 8101 3503 8282
rect 3449 8283 3450 8316
rect 3478 8101 3479 8284
rect 3452 8285 3453 8316
rect 3481 8101 3482 8286
rect 3455 8287 3456 8316
rect 3481 8287 3482 8316
rect 3461 8289 3462 8316
rect 3515 8289 3516 8316
rect 3463 8101 3464 8292
rect 3531 8291 3532 8316
rect 3464 8293 3465 8316
rect 3520 8101 3521 8294
rect 3474 8295 3475 8316
rect 3529 8101 3530 8296
rect 3490 8101 3491 8298
rect 3635 8101 3636 8298
rect 3493 8101 3494 8300
rect 3552 8101 3553 8300
rect 3494 8301 3495 8316
rect 3575 8101 3576 8302
rect 3506 8303 3507 8316
rect 3587 8101 3588 8304
rect 3509 8305 3510 8316
rect 3590 8101 3591 8306
rect 3517 8101 3518 8308
rect 3603 8101 3604 8308
rect 3525 8309 3526 8316
rect 3569 8101 3570 8310
rect 3528 8311 3529 8316
rect 3572 8101 3573 8312
rect 3642 8101 3643 8312
rect 3649 8101 3650 8312
rect 3645 8101 3646 8314
rect 3659 8101 3660 8314
rect 2821 8322 2822 8511
rect 2975 8320 2976 8323
rect 2917 8320 2918 8325
rect 3021 8320 3022 8325
rect 2917 8326 2918 8511
rect 3170 8320 3171 8327
rect 2924 8320 2925 8329
rect 3065 8320 3066 8329
rect 2927 8320 2928 8331
rect 3017 8330 3018 8511
rect 2931 8332 2932 8511
rect 3167 8320 3168 8333
rect 2934 8320 2935 8335
rect 3086 8334 3087 8511
rect 2953 8320 2954 8337
rect 3074 8320 3075 8337
rect 2953 8338 2954 8511
rect 3140 8320 3141 8339
rect 2969 8320 2970 8341
rect 3131 8320 3132 8341
rect 2972 8320 2973 8343
rect 2976 8342 2977 8511
rect 2979 8342 2980 8511
rect 3098 8320 3099 8343
rect 2981 8320 2982 8345
rect 3056 8320 3057 8345
rect 2988 8346 2989 8511
rect 3062 8320 3063 8347
rect 2991 8348 2992 8511
rect 3098 8348 3099 8511
rect 2997 8320 2998 8351
rect 3077 8320 3078 8351
rect 2950 8320 2951 8353
rect 3077 8352 3078 8511
rect 2950 8354 2951 8511
rect 3074 8354 3075 8511
rect 3003 8320 3004 8357
rect 3053 8356 3054 8511
rect 3002 8358 3003 8511
rect 3413 8320 3414 8359
rect 3005 8360 3006 8511
rect 3245 8320 3246 8361
rect 3008 8362 3009 8511
rect 3101 8320 3102 8363
rect 3014 8364 3015 8511
rect 3095 8320 3096 8365
rect 3024 8320 3025 8367
rect 3080 8320 3081 8367
rect 3023 8368 3024 8511
rect 3031 8320 3032 8369
rect 3032 8370 3033 8511
rect 3134 8320 3135 8371
rect 3038 8320 3039 8373
rect 3410 8320 3411 8373
rect 2960 8374 2961 8511
rect 3038 8374 3039 8511
rect 3041 8374 3042 8511
rect 3143 8320 3144 8375
rect 3044 8376 3045 8511
rect 3158 8320 3159 8377
rect 3050 8378 3051 8511
rect 3164 8320 3165 8379
rect 3056 8380 3057 8511
rect 3119 8320 3120 8381
rect 3062 8382 3063 8511
rect 3152 8320 3153 8383
rect 3068 8320 3069 8385
rect 3404 8320 3405 8385
rect 3092 8386 3093 8511
rect 3242 8320 3243 8387
rect 3095 8388 3096 8511
rect 3182 8320 3183 8389
rect 3104 8390 3105 8511
rect 3212 8320 3213 8391
rect 3107 8392 3108 8511
rect 3215 8320 3216 8393
rect 3110 8394 3111 8511
rect 3227 8320 3228 8395
rect 3089 8320 3090 8397
rect 3228 8396 3229 8511
rect 3089 8398 3090 8511
rect 3173 8320 3174 8399
rect 3113 8400 3114 8511
rect 3150 8400 3151 8511
rect 3120 8402 3121 8511
rect 3287 8320 3288 8403
rect 3123 8404 3124 8511
rect 3272 8320 3273 8405
rect 3132 8406 3133 8511
rect 3218 8320 3219 8407
rect 3138 8408 3139 8511
rect 3224 8320 3225 8409
rect 3144 8410 3145 8511
rect 3293 8320 3294 8411
rect 3153 8412 3154 8511
rect 3194 8320 3195 8413
rect 3156 8414 3157 8511
rect 3254 8320 3255 8415
rect 3162 8416 3163 8511
rect 3299 8320 3300 8417
rect 3174 8418 3175 8511
rect 3290 8320 3291 8419
rect 3183 8420 3184 8511
rect 3230 8320 3231 8421
rect 3186 8422 3187 8511
rect 3260 8320 3261 8423
rect 3188 8320 3189 8425
rect 3416 8320 3417 8425
rect 3195 8426 3196 8511
rect 3320 8320 3321 8427
rect 3200 8320 3201 8429
rect 3522 8320 3523 8429
rect 3210 8430 3211 8511
rect 3292 8430 3293 8511
rect 3213 8432 3214 8511
rect 3236 8320 3237 8433
rect 3216 8434 3217 8511
rect 3323 8320 3324 8435
rect 3234 8436 3235 8511
rect 3365 8320 3366 8437
rect 3246 8438 3247 8511
rect 3377 8320 3378 8439
rect 3189 8440 3190 8511
rect 3376 8440 3377 8511
rect 3248 8320 3249 8443
rect 3325 8442 3326 8511
rect 3249 8444 3250 8511
rect 3398 8320 3399 8445
rect 3252 8446 3253 8511
rect 3401 8320 3402 8447
rect 3255 8448 3256 8511
rect 3359 8320 3360 8449
rect 3258 8450 3259 8511
rect 3362 8320 3363 8451
rect 3263 8320 3264 8453
rect 3419 8320 3420 8453
rect 3266 8320 3267 8455
rect 3477 8320 3478 8455
rect 3267 8456 3268 8511
rect 3344 8456 3345 8511
rect 3270 8458 3271 8511
rect 3389 8320 3390 8459
rect 3273 8460 3274 8511
rect 3296 8320 3297 8461
rect 3275 8320 3276 8463
rect 3455 8320 3456 8463
rect 3276 8464 3277 8511
rect 3407 8320 3408 8465
rect 3279 8466 3280 8511
rect 3425 8320 3426 8467
rect 3281 8320 3282 8469
rect 3337 8468 3338 8511
rect 3177 8470 3178 8511
rect 3282 8470 3283 8511
rect 3295 8470 3296 8511
rect 3422 8320 3423 8471
rect 3304 8472 3305 8511
rect 3437 8320 3438 8473
rect 3307 8474 3308 8511
rect 3440 8320 3441 8475
rect 3311 8320 3312 8477
rect 3319 8476 3320 8511
rect 3317 8320 3318 8479
rect 3474 8320 3475 8479
rect 3316 8480 3317 8511
rect 3449 8320 3450 8481
rect 3329 8320 3330 8483
rect 3481 8320 3482 8483
rect 3328 8484 3329 8511
rect 3461 8320 3462 8485
rect 3331 8486 3332 8511
rect 3464 8320 3465 8487
rect 3341 8320 3342 8489
rect 3383 8488 3384 8511
rect 3358 8490 3359 8511
rect 3515 8320 3516 8491
rect 3367 8492 3368 8511
rect 3506 8320 3507 8493
rect 3370 8494 3371 8511
rect 3509 8320 3510 8495
rect 3386 8320 3387 8497
rect 3491 8320 3492 8497
rect 3386 8498 3387 8511
rect 3525 8320 3526 8499
rect 3392 8320 3393 8501
rect 3559 8320 3560 8501
rect 3406 8502 3407 8511
rect 3528 8320 3529 8503
rect 3417 8504 3418 8511
rect 3494 8320 3495 8505
rect 3428 8320 3429 8507
rect 3562 8320 3563 8507
rect 3452 8320 3453 8509
rect 3470 8320 3471 8509
rect 3548 8320 3549 8509
rect 3552 8320 3553 8509
rect 2815 8515 2816 8518
rect 2821 8515 2822 8518
rect 2881 8517 2882 8654
rect 2891 8517 2892 8654
rect 2917 8515 2918 8518
rect 3123 8515 3124 8518
rect 2920 8515 2921 8520
rect 3041 8515 3042 8520
rect 2933 8521 2934 8654
rect 3142 8521 3143 8654
rect 2941 8515 2942 8524
rect 3107 8515 3108 8524
rect 2945 8525 2946 8654
rect 3174 8515 3175 8526
rect 2952 8527 2953 8654
rect 3074 8515 3075 8528
rect 2960 8515 2961 8530
rect 3032 8515 3033 8530
rect 2962 8531 2963 8654
rect 3077 8515 3078 8532
rect 2968 8533 2969 8654
rect 3092 8515 3093 8534
rect 2972 8515 2973 8536
rect 2993 8535 2994 8654
rect 2991 8515 2992 8538
rect 3053 8515 3054 8538
rect 2990 8539 2991 8654
rect 3014 8515 3015 8540
rect 2995 8515 2996 8542
rect 3089 8515 3090 8542
rect 3002 8543 3003 8654
rect 3017 8515 3018 8544
rect 2931 8515 2932 8546
rect 3017 8545 3018 8654
rect 3005 8515 3006 8548
rect 3153 8515 3154 8548
rect 3005 8549 3006 8654
rect 3038 8515 3039 8550
rect 3008 8515 3009 8552
rect 3023 8515 3024 8552
rect 3008 8553 3009 8654
rect 3044 8515 3045 8554
rect 2998 8515 2999 8556
rect 3044 8555 3045 8654
rect 2924 8515 2925 8558
rect 2999 8557 3000 8654
rect 3014 8557 3015 8654
rect 3050 8515 3051 8558
rect 3026 8559 3027 8654
rect 3056 8515 3057 8560
rect 3032 8561 3033 8654
rect 3062 8515 3063 8562
rect 3038 8563 3039 8654
rect 3095 8515 3096 8564
rect 3041 8565 3042 8654
rect 3086 8515 3087 8566
rect 3053 8567 3054 8654
rect 3104 8515 3105 8568
rect 3056 8569 3057 8654
rect 3098 8515 3099 8570
rect 3059 8571 3060 8654
rect 3132 8515 3133 8572
rect 3062 8573 3063 8654
rect 3183 8515 3184 8574
rect 3065 8575 3066 8654
rect 3138 8515 3139 8576
rect 3068 8577 3069 8654
rect 3270 8515 3271 8578
rect 3071 8579 3072 8654
rect 3252 8515 3253 8580
rect 3074 8581 3075 8654
rect 3144 8515 3145 8582
rect 3080 8583 3081 8654
rect 3348 8515 3349 8584
rect 3086 8585 3087 8654
rect 3156 8515 3157 8586
rect 3092 8587 3093 8654
rect 3162 8515 3163 8588
rect 3101 8589 3102 8654
rect 3334 8515 3335 8590
rect 3104 8591 3105 8654
rect 3292 8515 3293 8592
rect 3107 8593 3108 8654
rect 3186 8515 3187 8594
rect 3117 8515 3118 8596
rect 3125 8595 3126 8654
rect 3116 8597 3117 8654
rect 3276 8515 3277 8598
rect 3119 8599 3120 8654
rect 3189 8515 3190 8600
rect 3122 8601 3123 8654
rect 3341 8515 3342 8602
rect 3128 8603 3129 8654
rect 3150 8515 3151 8604
rect 3132 8605 3133 8654
rect 3177 8515 3178 8606
rect 3145 8607 3146 8654
rect 3258 8515 3259 8608
rect 3151 8609 3152 8654
rect 3319 8515 3320 8610
rect 3161 8611 3162 8654
rect 3267 8515 3268 8612
rect 3167 8613 3168 8654
rect 3328 8515 3329 8614
rect 3171 8615 3172 8654
rect 3331 8515 3332 8616
rect 3174 8617 3175 8654
rect 3216 8515 3217 8618
rect 3178 8619 3179 8654
rect 3273 8515 3274 8620
rect 3184 8621 3185 8654
rect 3279 8515 3280 8622
rect 3187 8623 3188 8654
rect 3295 8515 3296 8624
rect 3190 8625 3191 8654
rect 3316 8515 3317 8626
rect 3193 8627 3194 8654
rect 3386 8515 3387 8628
rect 3195 8515 3196 8630
rect 3344 8515 3345 8630
rect 3210 8515 3211 8632
rect 3325 8515 3326 8632
rect 3213 8515 3214 8634
rect 3322 8515 3323 8634
rect 3228 8515 3229 8636
rect 3285 8515 3286 8636
rect 3234 8515 3235 8638
rect 3383 8515 3384 8638
rect 3246 8515 3247 8640
rect 3399 8515 3400 8640
rect 3249 8515 3250 8642
rect 3380 8515 3381 8642
rect 3255 8515 3256 8644
rect 3376 8515 3377 8644
rect 3304 8515 3305 8646
rect 3389 8515 3390 8646
rect 3307 8515 3308 8648
rect 3413 8515 3414 8648
rect 3367 8515 3368 8650
rect 3420 8515 3421 8650
rect 3370 8515 3371 8652
rect 3417 8515 3418 8652
rect 2884 8658 2885 8661
rect 2891 8658 2892 8661
rect 2881 8658 2882 8663
rect 2891 8662 2892 8735
rect 2882 8664 2883 8735
rect 2888 8664 2889 8735
rect 2923 8658 2924 8665
rect 3002 8658 3003 8665
rect 2930 8658 2931 8667
rect 3014 8658 3015 8667
rect 2933 8658 2934 8669
rect 3008 8658 3009 8669
rect 2942 8658 2943 8671
rect 2999 8658 3000 8671
rect 2949 8658 2950 8673
rect 2962 8658 2963 8673
rect 2956 8658 2957 8675
rect 3038 8658 3039 8675
rect 2959 8658 2960 8677
rect 3005 8658 3006 8677
rect 2965 8678 2966 8735
rect 2990 8658 2991 8679
rect 2968 8658 2969 8681
rect 3000 8680 3001 8735
rect 2972 8658 2973 8683
rect 3044 8658 3045 8683
rect 2981 8684 2982 8735
rect 3056 8658 3057 8685
rect 2993 8658 2994 8687
rect 3041 8658 3042 8687
rect 2984 8658 2985 8689
rect 2993 8688 2994 8735
rect 2984 8690 2985 8735
rect 3026 8658 3027 8691
rect 2996 8658 2997 8693
rect 3032 8658 3033 8693
rect 2987 8694 2988 8735
rect 2997 8694 2998 8735
rect 3003 8694 3004 8735
rect 3015 8694 3016 8735
rect 3006 8696 3007 8735
rect 3074 8658 3075 8697
rect 3017 8658 3018 8699
rect 3142 8658 3143 8699
rect 3018 8700 3019 8735
rect 3128 8658 3129 8701
rect 3030 8702 3031 8735
rect 3051 8702 3052 8735
rect 3042 8704 3043 8735
rect 3119 8658 3120 8705
rect 3045 8706 3046 8735
rect 3080 8658 3081 8707
rect 3053 8658 3054 8709
rect 3071 8658 3072 8709
rect 3055 8710 3056 8735
rect 3086 8658 3087 8711
rect 3059 8658 3060 8713
rect 3065 8658 3066 8713
rect 3058 8714 3059 8735
rect 3107 8658 3108 8715
rect 3092 8658 3093 8717
rect 3139 8658 3140 8717
rect 3101 8658 3102 8719
rect 3167 8658 3168 8719
rect 3104 8658 3105 8721
rect 3125 8658 3126 8721
rect 3116 8658 3117 8723
rect 3158 8658 3159 8723
rect 3122 8658 3123 8725
rect 3164 8658 3165 8725
rect 3145 8658 3146 8727
rect 3171 8658 3172 8727
rect 3161 8658 3162 8729
rect 3187 8658 3188 8729
rect 3184 8658 3185 8731
rect 3206 8658 3207 8731
rect 3193 8658 3194 8733
rect 3199 8658 3200 8733
rect 2875 8739 2876 8742
rect 2888 8739 2889 8742
rect 2882 8739 2883 8744
rect 2891 8739 2892 8744
rect 2917 8739 2918 8744
rect 2924 8739 2925 8744
rect 2962 8739 2963 8744
rect 2965 8739 2966 8744
rect 2968 8739 2969 8744
rect 3006 8739 3007 8744
rect 2971 8739 2972 8746
rect 2981 8739 2982 8746
rect 2975 8739 2976 8748
rect 2984 8739 2985 8748
rect 2987 8739 2988 8748
rect 2993 8739 2994 8748
rect 2997 8739 2998 8748
rect 3003 8739 3004 8748
rect 3012 8739 3013 8748
rect 3030 8739 3031 8748
rect 3015 8739 3016 8750
rect 3027 8739 3028 8750
rect 3018 8739 3019 8752
rect 3055 8739 3056 8752
rect 3042 8739 3043 8754
rect 3051 8739 3052 8754
rect 3045 8739 3046 8756
rect 3048 8739 3049 8756
<< via >>
rect 2941 1415 2942 1416
rect 2963 1415 2964 1416
rect 2944 1417 2945 1418
rect 3035 1417 3036 1418
rect 2947 1419 2948 1420
rect 2953 1419 2954 1420
rect 2957 1419 2958 1420
rect 2978 1419 2979 1420
rect 2960 1421 2961 1422
rect 2999 1421 3000 1422
rect 2966 1423 2967 1424
rect 3005 1423 3006 1424
rect 2984 1425 2985 1426
rect 3002 1425 3003 1426
rect 2987 1427 2988 1428
rect 2996 1427 2997 1428
rect 3011 1427 3012 1428
rect 3014 1427 3015 1428
rect 3017 1427 3018 1428
rect 3020 1427 3021 1428
rect 3026 1427 3027 1428
rect 3032 1427 3033 1428
rect 3044 1427 3045 1428
rect 3050 1427 3051 1428
rect 3047 1429 3048 1430
rect 3059 1429 3060 1430
rect 3056 1431 3057 1432
rect 3068 1431 3069 1432
rect 2809 1441 2810 1442
rect 3242 1441 3243 1442
rect 2938 1443 2939 1444
rect 2990 1443 2991 1444
rect 2944 1445 2945 1446
rect 3114 1445 3115 1446
rect 2947 1447 2948 1448
rect 2967 1447 2968 1448
rect 2953 1449 2954 1450
rect 2980 1449 2981 1450
rect 2973 1451 2974 1452
rect 3084 1451 3085 1452
rect 2978 1453 2979 1454
rect 3030 1453 3031 1454
rect 2984 1455 2985 1456
rect 3017 1455 3018 1456
rect 2987 1457 2988 1458
rect 3102 1457 3103 1458
rect 2987 1459 2988 1460
rect 3054 1459 3055 1460
rect 2993 1461 2994 1462
rect 3174 1461 3175 1462
rect 2996 1463 2997 1464
rect 3060 1463 3061 1464
rect 2999 1465 3000 1466
rect 3063 1465 3064 1466
rect 3000 1467 3001 1468
rect 3014 1467 3015 1468
rect 2950 1469 2951 1470
rect 3015 1469 3016 1470
rect 3002 1471 3003 1472
rect 3066 1471 3067 1472
rect 3005 1473 3006 1474
rect 3069 1473 3070 1474
rect 3011 1475 3012 1476
rect 3018 1475 3019 1476
rect 2963 1477 2964 1478
rect 3012 1477 3013 1478
rect 2952 1479 2953 1480
rect 2964 1479 2965 1480
rect 3023 1479 3024 1480
rect 3087 1479 3088 1480
rect 3026 1481 3027 1482
rect 3093 1481 3094 1482
rect 2931 1483 2932 1484
rect 3027 1483 3028 1484
rect 3035 1483 3036 1484
rect 3120 1483 3121 1484
rect 3036 1485 3037 1486
rect 3129 1485 3130 1486
rect 3039 1487 3040 1488
rect 3090 1487 3091 1488
rect 3044 1489 3045 1490
rect 3111 1489 3112 1490
rect 3047 1491 3048 1492
rect 3126 1491 3127 1492
rect 3056 1493 3057 1494
rect 3144 1493 3145 1494
rect 3150 1493 3151 1494
rect 3236 1493 3237 1494
rect 3153 1495 3154 1496
rect 3183 1495 3184 1496
rect 3156 1497 3157 1498
rect 3211 1497 3212 1498
rect 3165 1499 3166 1500
rect 3225 1499 3226 1500
rect 3177 1501 3178 1502
rect 3229 1501 3230 1502
rect 3190 1503 3191 1504
rect 3197 1503 3198 1504
rect 3204 1503 3205 1504
rect 3251 1503 3252 1504
rect 2920 1512 2921 1513
rect 2986 1512 2987 1513
rect 2920 1514 2921 1515
rect 2993 1514 2994 1515
rect 2936 1516 2937 1517
rect 3124 1516 3125 1517
rect 2938 1518 2939 1519
rect 3256 1518 3257 1519
rect 2934 1520 2935 1521
rect 2939 1520 2940 1521
rect 2933 1522 2934 1523
rect 2948 1522 2949 1523
rect 2917 1524 2918 1525
rect 2948 1524 2949 1525
rect 2941 1526 2942 1527
rect 3253 1526 3254 1527
rect 2955 1528 2956 1529
rect 3001 1528 3002 1529
rect 2809 1530 2810 1531
rect 2954 1530 2955 1531
rect 2957 1530 2958 1531
rect 3063 1530 3064 1531
rect 2924 1532 2925 1533
rect 3064 1532 3065 1533
rect 2960 1534 2961 1535
rect 3076 1534 3077 1535
rect 2964 1536 2965 1537
rect 2973 1536 2974 1537
rect 2970 1538 2971 1539
rect 3007 1538 3008 1539
rect 2971 1540 2972 1541
rect 3331 1540 3332 1541
rect 2990 1542 2991 1543
rect 3058 1542 3059 1543
rect 3015 1544 3016 1545
rect 3079 1544 3080 1545
rect 2967 1546 2968 1547
rect 3016 1546 3017 1547
rect 3018 1546 3019 1547
rect 3042 1546 3043 1547
rect 3025 1548 3026 1549
rect 3030 1548 3031 1549
rect 3035 1548 3036 1549
rect 3343 1548 3344 1549
rect 3046 1550 3047 1551
rect 3160 1550 3161 1551
rect 3069 1552 3070 1553
rect 3133 1552 3134 1553
rect 3072 1554 3073 1555
rect 3093 1554 3094 1555
rect 2984 1556 2985 1557
rect 3094 1556 3095 1557
rect 2917 1558 2918 1559
rect 2983 1558 2984 1559
rect 3084 1558 3085 1559
rect 3169 1558 3170 1559
rect 3087 1560 3088 1561
rect 3181 1560 3182 1561
rect 3102 1562 3103 1563
rect 3196 1562 3197 1563
rect 3111 1564 3112 1565
rect 3277 1564 3278 1565
rect 3114 1566 3115 1567
rect 3205 1566 3206 1567
rect 2931 1568 2932 1569
rect 3115 1568 3116 1569
rect 2930 1570 2931 1571
rect 3215 1570 3216 1571
rect 3120 1572 3121 1573
rect 3211 1572 3212 1573
rect 3027 1574 3028 1575
rect 3121 1574 3122 1575
rect 3126 1574 3127 1575
rect 3229 1574 3230 1575
rect 3032 1576 3033 1577
rect 3127 1576 3128 1577
rect 3129 1576 3130 1577
rect 3346 1576 3347 1577
rect 2977 1578 2978 1579
rect 3130 1578 3131 1579
rect 3141 1578 3142 1579
rect 3202 1578 3203 1579
rect 3142 1580 3143 1581
rect 3361 1580 3362 1581
rect 3144 1582 3145 1583
rect 3399 1582 3400 1583
rect 3054 1584 3055 1585
rect 3145 1584 3146 1585
rect 3150 1584 3151 1585
rect 3355 1584 3356 1585
rect 3066 1586 3067 1587
rect 3151 1586 3152 1587
rect 3153 1586 3154 1587
rect 3358 1586 3359 1587
rect 2998 1588 2999 1589
rect 3154 1588 3155 1589
rect 3156 1588 3157 1589
rect 3283 1588 3284 1589
rect 3060 1590 3061 1591
rect 3157 1590 3158 1591
rect 2902 1592 2903 1593
rect 3061 1592 3062 1593
rect 3162 1592 3163 1593
rect 3217 1592 3218 1593
rect 3165 1594 3166 1595
rect 3271 1594 3272 1595
rect 3174 1596 3175 1597
rect 3310 1596 3311 1597
rect 3175 1598 3176 1599
rect 3378 1598 3379 1599
rect 3177 1600 3178 1601
rect 3313 1600 3314 1601
rect 3178 1602 3179 1603
rect 3193 1602 3194 1603
rect 3183 1604 3184 1605
rect 3247 1604 3248 1605
rect 3090 1606 3091 1607
rect 3184 1606 3185 1607
rect 3012 1608 3013 1609
rect 3091 1608 3092 1609
rect 2974 1610 2975 1611
rect 3013 1610 3014 1611
rect 3187 1610 3188 1611
rect 3375 1610 3376 1611
rect 3222 1612 3223 1613
rect 3325 1612 3326 1613
rect 3225 1614 3226 1615
rect 3316 1614 3317 1615
rect 3236 1616 3237 1617
rect 3328 1616 3329 1617
rect 3241 1618 3242 1619
rect 3385 1618 3386 1619
rect 3259 1620 3260 1621
rect 3417 1620 3418 1621
rect 3274 1622 3275 1623
rect 3406 1622 3407 1623
rect 3295 1624 3296 1625
rect 3434 1624 3435 1625
rect 3319 1626 3320 1627
rect 3382 1626 3383 1627
rect 3322 1628 3323 1629
rect 3403 1628 3404 1629
rect 2894 1637 2895 1638
rect 3450 1637 3451 1638
rect 2917 1639 2918 1640
rect 2941 1639 2942 1640
rect 2933 1641 2934 1642
rect 2977 1641 2978 1642
rect 2932 1643 2933 1644
rect 3145 1643 3146 1644
rect 2944 1645 2945 1646
rect 2971 1645 2972 1646
rect 2930 1647 2931 1648
rect 2971 1647 2972 1648
rect 2954 1649 2955 1650
rect 3005 1649 3006 1650
rect 2948 1651 2949 1652
rect 2953 1651 2954 1652
rect 2974 1651 2975 1652
rect 3053 1651 3054 1652
rect 2881 1653 2882 1654
rect 2974 1653 2975 1654
rect 2983 1653 2984 1654
rect 3032 1653 3033 1654
rect 2990 1655 2991 1656
rect 3138 1655 3139 1656
rect 3010 1657 3011 1658
rect 3207 1657 3208 1658
rect 3011 1659 3012 1660
rect 3160 1659 3161 1660
rect 3035 1661 3036 1662
rect 3501 1661 3502 1662
rect 2986 1663 2987 1664
rect 3035 1663 3036 1664
rect 2987 1665 2988 1666
rect 3079 1665 3080 1666
rect 2929 1667 2930 1668
rect 3080 1667 3081 1668
rect 3039 1669 3040 1670
rect 3225 1669 3226 1670
rect 2922 1671 2923 1672
rect 3038 1671 3039 1672
rect 3041 1671 3042 1672
rect 3070 1671 3071 1672
rect 3007 1673 3008 1674
rect 3071 1673 3072 1674
rect 3046 1675 3047 1676
rect 3178 1675 3179 1676
rect 3049 1677 3050 1678
rect 3144 1677 3145 1678
rect 2902 1679 2903 1680
rect 3050 1679 3051 1680
rect 3058 1679 3059 1680
rect 3105 1679 3106 1680
rect 3013 1681 3014 1682
rect 3059 1681 3060 1682
rect 3001 1683 3002 1684
rect 3014 1683 3015 1684
rect 3061 1683 3062 1684
rect 3147 1683 3148 1684
rect 3016 1685 3017 1686
rect 3062 1685 3063 1686
rect 3064 1685 3065 1686
rect 3117 1685 3118 1686
rect 3083 1687 3084 1688
rect 3448 1687 3449 1688
rect 3124 1689 3125 1690
rect 3171 1689 3172 1690
rect 3076 1691 3077 1692
rect 3123 1691 3124 1692
rect 2915 1693 2916 1694
rect 3077 1693 3078 1694
rect 3130 1693 3131 1694
rect 3213 1693 3214 1694
rect 3151 1695 3152 1696
rect 3198 1695 3199 1696
rect 3089 1697 3090 1698
rect 3150 1697 3151 1698
rect 3175 1697 3176 1698
rect 3222 1697 3223 1698
rect 3127 1699 3128 1700
rect 3174 1699 3175 1700
rect 3184 1699 3185 1700
rect 3234 1699 3235 1700
rect 3190 1701 3191 1702
rect 3352 1701 3353 1702
rect 3142 1703 3143 1704
rect 3351 1703 3352 1704
rect 3094 1705 3095 1706
rect 3141 1705 3142 1706
rect 3093 1707 3094 1708
rect 3121 1707 3122 1708
rect 3193 1707 3194 1708
rect 3358 1707 3359 1708
rect 3202 1709 3203 1710
rect 3357 1709 3358 1710
rect 3154 1711 3155 1712
rect 3201 1711 3202 1712
rect 3205 1711 3206 1712
rect 3306 1711 3307 1712
rect 3157 1713 3158 1714
rect 3204 1713 3205 1714
rect 3211 1713 3212 1714
rect 3264 1713 3265 1714
rect 2998 1715 2999 1716
rect 3210 1715 3211 1716
rect 3229 1715 3230 1716
rect 3349 1715 3350 1716
rect 3181 1717 3182 1718
rect 3228 1717 3229 1718
rect 3133 1719 3134 1720
rect 3180 1719 3181 1720
rect 3091 1721 3092 1722
rect 3132 1721 3133 1722
rect 3187 1721 3188 1722
rect 3348 1721 3349 1722
rect 3025 1723 3026 1724
rect 3186 1723 3187 1724
rect 2925 1725 2926 1726
rect 3026 1725 3027 1726
rect 3231 1725 3232 1726
rect 3360 1725 3361 1726
rect 3247 1727 3248 1728
rect 3465 1727 3466 1728
rect 3196 1729 3197 1730
rect 3246 1729 3247 1730
rect 3253 1729 3254 1730
rect 3336 1729 3337 1730
rect 3256 1731 3257 1732
rect 3339 1731 3340 1732
rect 3271 1733 3272 1734
rect 3406 1733 3407 1734
rect 3270 1735 3271 1736
rect 3371 1735 3372 1736
rect 3274 1737 3275 1738
rect 3514 1737 3515 1738
rect 3283 1739 3284 1740
rect 3384 1739 3385 1740
rect 3295 1741 3296 1742
rect 3375 1741 3376 1742
rect 3217 1743 3218 1744
rect 3294 1743 3295 1744
rect 3028 1745 3029 1746
rect 3216 1745 3217 1746
rect 3300 1745 3301 1746
rect 3417 1745 3418 1746
rect 3310 1747 3311 1748
rect 3402 1747 3403 1748
rect 3313 1749 3314 1750
rect 3405 1749 3406 1750
rect 3312 1751 3313 1752
rect 3525 1751 3526 1752
rect 3316 1753 3317 1754
rect 3471 1753 3472 1754
rect 3315 1755 3316 1756
rect 3389 1755 3390 1756
rect 3319 1757 3320 1758
rect 3420 1757 3421 1758
rect 3255 1759 3256 1760
rect 3318 1759 3319 1760
rect 3322 1759 3323 1760
rect 3423 1759 3424 1760
rect 3325 1761 3326 1762
rect 3408 1761 3409 1762
rect 3241 1763 3242 1764
rect 3324 1763 3325 1764
rect 3073 1765 3074 1766
rect 3240 1765 3241 1766
rect 3331 1765 3332 1766
rect 3432 1765 3433 1766
rect 3343 1767 3344 1768
rect 3453 1767 3454 1768
rect 3259 1769 3260 1770
rect 3342 1769 3343 1770
rect 3346 1769 3347 1770
rect 3438 1769 3439 1770
rect 3355 1771 3356 1772
rect 3456 1771 3457 1772
rect 3354 1773 3355 1774
rect 3363 1773 3364 1774
rect 3372 1773 3373 1774
rect 3410 1773 3411 1774
rect 3328 1775 3329 1776
rect 3411 1775 3412 1776
rect 3378 1777 3379 1778
rect 3459 1777 3460 1778
rect 3277 1779 3278 1780
rect 3378 1779 3379 1780
rect 3276 1781 3277 1782
rect 3392 1781 3393 1782
rect 3468 1781 3469 1782
rect 3477 1781 3478 1782
rect 3552 1781 3553 1782
rect 3572 1781 3573 1782
rect 2863 1790 2864 1791
rect 2974 1790 2975 1791
rect 2866 1792 2867 1793
rect 2870 1792 2871 1793
rect 2884 1792 2885 1793
rect 2888 1792 2889 1793
rect 2894 1792 2895 1793
rect 2932 1792 2933 1793
rect 2901 1794 2902 1795
rect 3067 1794 3068 1795
rect 2904 1796 2905 1797
rect 3050 1796 3051 1797
rect 2914 1798 2915 1799
rect 3077 1798 3078 1799
rect 2918 1800 2919 1801
rect 3123 1800 3124 1801
rect 2922 1802 2923 1803
rect 3043 1802 3044 1803
rect 2925 1804 2926 1805
rect 3041 1804 3042 1805
rect 2928 1806 2929 1807
rect 3064 1806 3065 1807
rect 2953 1808 2954 1809
rect 2998 1808 2999 1809
rect 2959 1810 2960 1811
rect 3196 1810 3197 1811
rect 2962 1812 2963 1813
rect 2987 1812 2988 1813
rect 2968 1814 2969 1815
rect 3168 1814 3169 1815
rect 2971 1816 2972 1817
rect 2995 1816 2996 1817
rect 2983 1818 2984 1819
rect 3062 1818 3063 1819
rect 2990 1820 2991 1821
rect 3132 1820 3133 1821
rect 2989 1822 2990 1823
rect 3035 1822 3036 1823
rect 3007 1824 3008 1825
rect 3038 1824 3039 1825
rect 3014 1826 3015 1827
rect 3073 1826 3074 1827
rect 3026 1828 3027 1829
rect 3055 1828 3056 1829
rect 3032 1830 3033 1831
rect 3049 1830 3050 1831
rect 3005 1832 3006 1833
rect 3031 1832 3032 1833
rect 3004 1834 3005 1835
rect 3178 1834 3179 1835
rect 3034 1836 3035 1837
rect 3171 1836 3172 1837
rect 3053 1838 3054 1839
rect 3085 1838 3086 1839
rect 2941 1840 2942 1841
rect 3052 1840 3053 1841
rect 2940 1842 2941 1843
rect 3011 1842 3012 1843
rect 2977 1844 2978 1845
rect 3010 1844 3011 1845
rect 2977 1846 2978 1847
rect 3130 1846 3131 1847
rect 3059 1848 3060 1849
rect 3091 1848 3092 1849
rect 3061 1850 3062 1851
rect 3577 1850 3578 1851
rect 3080 1852 3081 1853
rect 3100 1852 3101 1853
rect 3079 1854 3080 1855
rect 3511 1854 3512 1855
rect 3089 1856 3090 1857
rect 3213 1856 3214 1857
rect 3096 1858 3097 1859
rect 3334 1858 3335 1859
rect 2917 1860 2918 1861
rect 3097 1860 3098 1861
rect 3111 1860 3112 1861
rect 3274 1860 3275 1861
rect 3136 1862 3137 1863
rect 3225 1862 3226 1863
rect 2911 1864 2912 1865
rect 3226 1864 3227 1865
rect 2910 1866 2911 1867
rect 3070 1866 3071 1867
rect 3138 1866 3139 1867
rect 3160 1866 3161 1867
rect 3141 1868 3142 1869
rect 3163 1868 3164 1869
rect 2897 1870 2898 1871
rect 3142 1870 3143 1871
rect 3144 1870 3145 1871
rect 3184 1870 3185 1871
rect 2903 1872 2904 1873
rect 3145 1872 3146 1873
rect 3166 1872 3167 1873
rect 3216 1872 3217 1873
rect 3169 1874 3170 1875
rect 3180 1874 3181 1875
rect 3174 1876 3175 1877
rect 3214 1876 3215 1877
rect 3186 1878 3187 1879
rect 3220 1878 3221 1879
rect 3190 1880 3191 1881
rect 3201 1880 3202 1881
rect 3112 1882 3113 1883
rect 3202 1882 3203 1883
rect 3204 1882 3205 1883
rect 3238 1882 3239 1883
rect 3210 1884 3211 1885
rect 3244 1884 3245 1885
rect 3222 1886 3223 1887
rect 3262 1886 3263 1887
rect 3231 1888 3232 1889
rect 3298 1888 3299 1889
rect 3198 1890 3199 1891
rect 3232 1890 3233 1891
rect 3147 1892 3148 1893
rect 3199 1892 3200 1893
rect 3117 1894 3118 1895
rect 3148 1894 3149 1895
rect 2921 1896 2922 1897
rect 3118 1896 3119 1897
rect 3234 1896 3235 1897
rect 3268 1896 3269 1897
rect 3235 1898 3236 1899
rect 3474 1898 3475 1899
rect 3240 1900 3241 1901
rect 3286 1900 3287 1901
rect 3207 1902 3208 1903
rect 3241 1902 3242 1903
rect 3109 1904 3110 1905
rect 3208 1904 3209 1905
rect 3246 1904 3247 1905
rect 3280 1904 3281 1905
rect 3150 1906 3151 1907
rect 3247 1906 3248 1907
rect 3255 1906 3256 1907
rect 3351 1906 3352 1907
rect 3264 1908 3265 1909
rect 3544 1908 3545 1909
rect 3016 1910 3017 1911
rect 3265 1910 3266 1911
rect 3270 1910 3271 1911
rect 3304 1910 3305 1911
rect 3276 1912 3277 1913
rect 3310 1912 3311 1913
rect 3294 1914 3295 1915
rect 3328 1914 3329 1915
rect 3300 1916 3301 1917
rect 3525 1916 3526 1917
rect 3114 1918 3115 1919
rect 3301 1918 3302 1919
rect 3083 1920 3084 1921
rect 3115 1920 3116 1921
rect 3306 1920 3307 1921
rect 3352 1920 3353 1921
rect 3322 1922 3323 1923
rect 3339 1922 3340 1923
rect 3312 1924 3313 1925
rect 3340 1924 3341 1925
rect 3324 1926 3325 1927
rect 3382 1926 3383 1927
rect 3336 1928 3337 1929
rect 3415 1928 3416 1929
rect 3348 1930 3349 1931
rect 3400 1930 3401 1931
rect 3354 1932 3355 1933
rect 3430 1932 3431 1933
rect 3370 1934 3371 1935
rect 3481 1934 3482 1935
rect 3384 1936 3385 1937
rect 3565 1936 3566 1937
rect 3402 1938 3403 1939
rect 3484 1938 3485 1939
rect 3318 1940 3319 1941
rect 3403 1940 3404 1941
rect 3405 1940 3406 1941
rect 3487 1940 3488 1941
rect 3408 1942 3409 1943
rect 3490 1942 3491 1943
rect 3411 1944 3412 1945
rect 3493 1944 3494 1945
rect 3412 1946 3413 1947
rect 3547 1946 3548 1947
rect 3420 1948 3421 1949
rect 3496 1948 3497 1949
rect 3375 1950 3376 1951
rect 3421 1950 3422 1951
rect 2896 1952 2897 1953
rect 3376 1952 3377 1953
rect 3423 1952 3424 1953
rect 3499 1952 3500 1953
rect 3342 1954 3343 1955
rect 3424 1954 3425 1955
rect 3315 1956 3316 1957
rect 3343 1956 3344 1957
rect 3438 1956 3439 1957
rect 3508 1956 3509 1957
rect 3448 1958 3449 1959
rect 3646 1958 3647 1959
rect 3450 1960 3451 1961
rect 3520 1960 3521 1961
rect 3372 1962 3373 1963
rect 3451 1962 3452 1963
rect 3453 1962 3454 1963
rect 3523 1962 3524 1963
rect 3378 1964 3379 1965
rect 3454 1964 3455 1965
rect 3456 1964 3457 1965
rect 3526 1964 3527 1965
rect 3459 1966 3460 1967
rect 3529 1966 3530 1967
rect 3468 1968 3469 1969
rect 3538 1968 3539 1969
rect 3471 1970 3472 1971
rect 3541 1970 3542 1971
rect 3552 1970 3553 1971
rect 3636 1970 3637 1971
rect 3418 1972 3419 1973
rect 3551 1972 3552 1973
rect 3558 1972 3559 1973
rect 3583 1972 3584 1973
rect 3228 1974 3229 1975
rect 3558 1974 3559 1975
rect 2980 1976 2981 1977
rect 3229 1976 3230 1977
rect 2980 1978 2981 1979
rect 3105 1978 3106 1979
rect 3562 1978 3563 1979
rect 3574 1978 3575 1979
rect 3572 1980 3573 1981
rect 3633 1980 3634 1981
rect 3501 1982 3502 1983
rect 3571 1982 3572 1983
rect 3432 1984 3433 1985
rect 3502 1984 3503 1985
rect 3357 1986 3358 1987
rect 3433 1986 3434 1987
rect 3358 1988 3359 1989
rect 3603 1988 3604 1989
rect 2866 1997 2867 1998
rect 3010 1997 3011 1998
rect 2896 1999 2897 2000
rect 3175 1999 3176 2000
rect 2903 2001 2904 2002
rect 2958 2001 2959 2002
rect 2870 2003 2871 2004
rect 2957 2003 2958 2004
rect 2902 2005 2903 2006
rect 3070 2005 3071 2006
rect 2909 2007 2910 2008
rect 3034 2007 3035 2008
rect 2915 2009 2916 2010
rect 3052 2009 3053 2010
rect 2921 2011 2922 2012
rect 3064 2011 3065 2012
rect 2924 2013 2925 2014
rect 3196 2013 3197 2014
rect 2934 2015 2935 2016
rect 3055 2015 3056 2016
rect 2940 2017 2941 2018
rect 3039 2017 3040 2018
rect 2961 2019 2962 2020
rect 3247 2019 3248 2020
rect 2960 2021 2961 2022
rect 3157 2021 3158 2022
rect 2963 2023 2964 2024
rect 3073 2023 3074 2024
rect 2966 2025 2967 2026
rect 2989 2025 2990 2026
rect 2968 2027 2969 2028
rect 3283 2027 3284 2028
rect 2972 2029 2973 2030
rect 2998 2029 2999 2030
rect 2977 2031 2978 2032
rect 3199 2031 3200 2032
rect 2984 2033 2985 2034
rect 3145 2033 3146 2034
rect 2995 2035 2996 2036
rect 3002 2035 3003 2036
rect 3005 2035 3006 2036
rect 3130 2035 3131 2036
rect 3016 2037 3017 2038
rect 3067 2037 3068 2038
rect 3017 2039 3018 2040
rect 3079 2039 3080 2040
rect 3020 2041 3021 2042
rect 3241 2041 3242 2042
rect 3023 2043 3024 2044
rect 3112 2043 3113 2044
rect 3025 2045 3026 2046
rect 3238 2045 3239 2046
rect 3028 2047 3029 2048
rect 3151 2047 3152 2048
rect 3033 2049 3034 2050
rect 3289 2049 3290 2050
rect 3036 2051 3037 2052
rect 3049 2051 3050 2052
rect 3043 2053 3044 2054
rect 3054 2053 3055 2054
rect 3031 2055 3032 2056
rect 3042 2055 3043 2056
rect 3030 2057 3031 2058
rect 3295 2057 3296 2058
rect 3051 2059 3052 2060
rect 3061 2059 3062 2060
rect 3070 2059 3071 2060
rect 3085 2059 3086 2060
rect 3076 2061 3077 2062
rect 3091 2061 3092 2062
rect 3100 2061 3101 2062
rect 3121 2061 3122 2062
rect 3109 2063 3110 2064
rect 3190 2063 3191 2064
rect 3118 2065 3119 2066
rect 3130 2065 3131 2066
rect 3097 2067 3098 2068
rect 3118 2067 3119 2068
rect 3124 2067 3125 2068
rect 3148 2067 3149 2068
rect 3142 2069 3143 2070
rect 3199 2069 3200 2070
rect 2931 2071 2932 2072
rect 3142 2071 3143 2072
rect 3160 2071 3161 2072
rect 3181 2071 3182 2072
rect 3166 2073 3167 2074
rect 3433 2073 3434 2074
rect 3169 2075 3170 2076
rect 3349 2075 3350 2076
rect 3169 2077 3170 2078
rect 3454 2077 3455 2078
rect 3178 2079 3179 2080
rect 3193 2079 3194 2080
rect 3115 2081 3116 2082
rect 3178 2081 3179 2082
rect 3184 2081 3185 2082
rect 3241 2081 3242 2082
rect 3163 2083 3164 2084
rect 3184 2083 3185 2084
rect 3139 2085 3140 2086
rect 3163 2085 3164 2086
rect 3187 2085 3188 2086
rect 3403 2085 3404 2086
rect 3202 2087 3203 2088
rect 3211 2087 3212 2088
rect 2900 2089 2901 2090
rect 3202 2089 3203 2090
rect 3208 2089 3209 2090
rect 3217 2089 3218 2090
rect 3226 2089 3227 2090
rect 3337 2089 3338 2090
rect 3232 2091 3233 2092
rect 3313 2091 3314 2092
rect 3235 2093 3236 2094
rect 3316 2093 3317 2094
rect 3220 2095 3221 2096
rect 3235 2095 3236 2096
rect 3244 2095 3245 2096
rect 3277 2095 3278 2096
rect 3244 2097 3245 2098
rect 3301 2097 3302 2098
rect 3250 2099 3251 2100
rect 3274 2099 3275 2100
rect 3250 2101 3251 2102
rect 3253 2101 3254 2102
rect 3253 2103 3254 2104
rect 3298 2103 3299 2104
rect 3214 2105 3215 2106
rect 3298 2105 3299 2106
rect 3256 2107 3257 2108
rect 3430 2107 3431 2108
rect 3262 2109 3263 2110
rect 3331 2109 3332 2110
rect 3265 2111 3266 2112
rect 3346 2111 3347 2112
rect 3268 2113 3269 2114
rect 3364 2113 3365 2114
rect 3286 2115 3287 2116
rect 3319 2115 3320 2116
rect 3307 2117 3308 2118
rect 3382 2117 3383 2118
rect 3280 2119 3281 2120
rect 3382 2119 3383 2120
rect 3310 2121 3311 2122
rect 3639 2121 3640 2122
rect 3322 2123 3323 2124
rect 3388 2123 3389 2124
rect 3340 2125 3341 2126
rect 3403 2125 3404 2126
rect 3229 2127 3230 2128
rect 3340 2127 3341 2128
rect 3229 2129 3230 2130
rect 3523 2129 3524 2130
rect 3343 2131 3344 2132
rect 3409 2131 3410 2132
rect 3103 2133 3104 2134
rect 3343 2133 3344 2134
rect 3352 2133 3353 2134
rect 3535 2133 3536 2134
rect 3358 2135 3359 2136
rect 3433 2135 3434 2136
rect 3328 2137 3329 2138
rect 3358 2137 3359 2138
rect 3367 2137 3368 2138
rect 3400 2137 3401 2138
rect 3376 2139 3377 2140
rect 3427 2139 3428 2140
rect 3376 2141 3377 2142
rect 3526 2141 3527 2142
rect 3379 2143 3380 2144
rect 3529 2143 3530 2144
rect 3385 2145 3386 2146
rect 3520 2145 3521 2146
rect 3400 2147 3401 2148
rect 3412 2147 3413 2148
rect 3418 2147 3419 2148
rect 3545 2147 3546 2148
rect 3418 2149 3419 2150
rect 3548 2149 3549 2150
rect 3424 2151 3425 2152
rect 3442 2151 3443 2152
rect 3439 2153 3440 2154
rect 3496 2153 3497 2154
rect 3448 2155 3449 2156
rect 3523 2155 3524 2156
rect 3415 2157 3416 2158
rect 3448 2157 3449 2158
rect 3415 2159 3416 2160
rect 3577 2159 3578 2160
rect 3445 2161 3446 2162
rect 3578 2161 3579 2162
rect 3481 2163 3482 2164
rect 3670 2163 3671 2164
rect 3484 2165 3485 2166
rect 3496 2165 3497 2166
rect 3451 2167 3452 2168
rect 3484 2167 3485 2168
rect 3451 2169 3452 2170
rect 3618 2169 3619 2170
rect 3490 2171 3491 2172
rect 3532 2171 3533 2172
rect 3421 2173 3422 2174
rect 3490 2173 3491 2174
rect 3370 2175 3371 2176
rect 3421 2175 3422 2176
rect 3304 2177 3305 2178
rect 3370 2177 3371 2178
rect 3493 2177 3494 2178
rect 3535 2177 3536 2178
rect 3493 2179 3494 2180
rect 3639 2179 3640 2180
rect 3499 2181 3500 2182
rect 3565 2181 3566 2182
rect 3487 2183 3488 2184
rect 3499 2183 3500 2184
rect 3502 2183 3503 2184
rect 3526 2183 3527 2184
rect 3508 2185 3509 2186
rect 3529 2185 3530 2186
rect 3514 2187 3515 2188
rect 3653 2187 3654 2188
rect 3520 2189 3521 2190
rect 3664 2189 3665 2190
rect 3538 2191 3539 2192
rect 3558 2191 3559 2192
rect 3325 2193 3326 2194
rect 3538 2193 3539 2194
rect 3555 2193 3556 2194
rect 3612 2193 3613 2194
rect 3561 2195 3562 2196
rect 3567 2195 3568 2196
rect 3541 2197 3542 2198
rect 3561 2197 3562 2198
rect 3265 2199 3266 2200
rect 3541 2199 3542 2200
rect 3571 2199 3572 2200
rect 3603 2199 3604 2200
rect 3574 2201 3575 2202
rect 3606 2201 3607 2202
rect 3583 2203 3584 2204
rect 3609 2203 3610 2204
rect 3591 2205 3592 2206
rect 3654 2205 3655 2206
rect 3633 2207 3634 2208
rect 3648 2207 3649 2208
rect 3636 2209 3637 2210
rect 3651 2209 3652 2210
rect 2902 2218 2903 2219
rect 3130 2218 3131 2219
rect 2915 2220 2916 2221
rect 3039 2220 3040 2221
rect 2924 2222 2925 2223
rect 3073 2222 3074 2223
rect 2923 2224 2924 2225
rect 3046 2224 3047 2225
rect 2927 2226 2928 2227
rect 3227 2226 3228 2227
rect 2927 2228 2928 2229
rect 3118 2228 3119 2229
rect 2934 2230 2935 2231
rect 3248 2230 3249 2231
rect 2933 2232 2934 2233
rect 2957 2232 2958 2233
rect 2961 2232 2962 2233
rect 2984 2232 2985 2233
rect 2964 2234 2965 2235
rect 3202 2234 3203 2235
rect 2966 2236 2967 2237
rect 3040 2236 3041 2237
rect 2972 2238 2973 2239
rect 2979 2238 2980 2239
rect 2985 2238 2986 2239
rect 3283 2238 3284 2239
rect 2988 2240 2989 2241
rect 3112 2240 3113 2241
rect 2993 2242 2994 2243
rect 3092 2242 3093 2243
rect 2992 2244 2993 2245
rect 3036 2244 3037 2245
rect 2920 2246 2921 2247
rect 3037 2246 3038 2247
rect 3004 2248 3005 2249
rect 3311 2248 3312 2249
rect 3007 2250 3008 2251
rect 3100 2250 3101 2251
rect 3020 2252 3021 2253
rect 3095 2252 3096 2253
rect 3017 2254 3018 2255
rect 3019 2254 3020 2255
rect 3002 2256 3003 2257
rect 3016 2256 3017 2257
rect 3023 2256 3024 2257
rect 3316 2256 3317 2257
rect 3030 2258 3031 2259
rect 3277 2258 3278 2259
rect 3031 2260 3032 2261
rect 3054 2260 3055 2261
rect 3042 2262 3043 2263
rect 3049 2262 3050 2263
rect 3043 2264 3044 2265
rect 3051 2264 3052 2265
rect 2906 2266 2907 2267
rect 3052 2266 3053 2267
rect 2906 2268 2907 2269
rect 3199 2268 3200 2269
rect 2967 2270 2968 2271
rect 3200 2270 3201 2271
rect 3060 2272 3061 2273
rect 3346 2272 3347 2273
rect 3061 2274 3062 2275
rect 3070 2274 3071 2275
rect 3067 2276 3068 2277
rect 3250 2276 3251 2277
rect 3067 2278 3068 2279
rect 3076 2278 3077 2279
rect 3076 2280 3077 2281
rect 3121 2280 3122 2281
rect 2995 2282 2996 2283
rect 3122 2282 3123 2283
rect 3079 2284 3080 2285
rect 3313 2284 3314 2285
rect 3098 2286 3099 2287
rect 3548 2286 3549 2287
rect 3103 2288 3104 2289
rect 3193 2288 3194 2289
rect 2902 2290 2903 2291
rect 3104 2290 3105 2291
rect 3116 2290 3117 2291
rect 3124 2290 3125 2291
rect 3128 2290 3129 2291
rect 3151 2290 3152 2291
rect 3140 2292 3141 2293
rect 3175 2292 3176 2293
rect 3142 2294 3143 2295
rect 3146 2294 3147 2295
rect 3143 2296 3144 2297
rect 3178 2296 3179 2297
rect 3157 2298 3158 2299
rect 3161 2298 3162 2299
rect 3169 2298 3170 2299
rect 3530 2298 3531 2299
rect 3173 2300 3174 2301
rect 3367 2300 3368 2301
rect 3176 2302 3177 2303
rect 3305 2302 3306 2303
rect 3179 2304 3180 2305
rect 3181 2304 3182 2305
rect 3182 2306 3183 2307
rect 3184 2306 3185 2307
rect 3187 2306 3188 2307
rect 3272 2306 3273 2307
rect 3197 2308 3198 2309
rect 3241 2308 3242 2309
rect 3203 2310 3204 2311
rect 3211 2310 3212 2311
rect 3163 2312 3164 2313
rect 3212 2312 3213 2313
rect 3209 2314 3210 2315
rect 3217 2314 3218 2315
rect 3215 2316 3216 2317
rect 3298 2316 3299 2317
rect 3229 2318 3230 2319
rect 3526 2318 3527 2319
rect 3233 2320 3234 2321
rect 3244 2320 3245 2321
rect 3239 2322 3240 2323
rect 3289 2322 3290 2323
rect 3245 2324 3246 2325
rect 3295 2324 3296 2325
rect 3251 2326 3252 2327
rect 3349 2326 3350 2327
rect 3256 2328 3257 2329
rect 3287 2328 3288 2329
rect 3088 2330 3089 2331
rect 3257 2330 3258 2331
rect 3089 2332 3090 2333
rect 3235 2332 3236 2333
rect 3236 2334 3237 2335
rect 3253 2334 3254 2335
rect 3263 2334 3264 2335
rect 3319 2334 3320 2335
rect 3265 2336 3266 2337
rect 3539 2336 3540 2337
rect 3275 2338 3276 2339
rect 3331 2338 3332 2339
rect 3281 2340 3282 2341
rect 3337 2340 3338 2341
rect 3284 2342 3285 2343
rect 3340 2342 3341 2343
rect 3290 2344 3291 2345
rect 3579 2344 3580 2345
rect 3296 2346 3297 2347
rect 3358 2346 3359 2347
rect 3302 2348 3303 2349
rect 3364 2348 3365 2349
rect 3307 2350 3308 2351
rect 3320 2350 3321 2351
rect 3325 2350 3326 2351
rect 3479 2350 3480 2351
rect 3326 2352 3327 2353
rect 3382 2352 3383 2353
rect 3332 2354 3333 2355
rect 3567 2354 3568 2355
rect 3338 2356 3339 2357
rect 3388 2356 3389 2357
rect 3343 2358 3344 2359
rect 3555 2358 3556 2359
rect 3350 2360 3351 2361
rect 3576 2360 3577 2361
rect 3353 2362 3354 2363
rect 3403 2362 3404 2363
rect 3359 2364 3360 2365
rect 3409 2364 3410 2365
rect 3365 2366 3366 2367
rect 3415 2366 3416 2367
rect 3370 2368 3371 2369
rect 3555 2368 3556 2369
rect 3371 2370 3372 2371
rect 3421 2370 3422 2371
rect 3379 2372 3380 2373
rect 3541 2372 3542 2373
rect 3383 2374 3384 2375
rect 3433 2374 3434 2375
rect 3385 2376 3386 2377
rect 3527 2376 3528 2377
rect 3392 2378 3393 2379
rect 3545 2378 3546 2379
rect 3400 2380 3401 2381
rect 3585 2380 3586 2381
rect 3401 2382 3402 2383
rect 3451 2382 3452 2383
rect 3057 2384 3058 2385
rect 3452 2384 3453 2385
rect 3437 2386 3438 2387
rect 3484 2386 3485 2387
rect 3439 2388 3440 2389
rect 3586 2388 3587 2389
rect 3442 2390 3443 2391
rect 3458 2390 3459 2391
rect 3445 2392 3446 2393
rect 3542 2392 3543 2393
rect 3448 2394 3449 2395
rect 3545 2394 3546 2395
rect 3418 2396 3419 2397
rect 3449 2396 3450 2397
rect 3455 2396 3456 2397
rect 3583 2396 3584 2397
rect 3473 2398 3474 2399
rect 3493 2398 3494 2399
rect 3476 2400 3477 2401
rect 3581 2400 3582 2401
rect 3481 2402 3482 2403
rect 3677 2402 3678 2403
rect 3485 2404 3486 2405
rect 3520 2404 3521 2405
rect 3490 2406 3491 2407
rect 3643 2406 3644 2407
rect 3503 2408 3504 2409
rect 3561 2408 3562 2409
rect 3509 2410 3510 2411
rect 3567 2410 3568 2411
rect 3514 2412 3515 2413
rect 3661 2412 3662 2413
rect 3521 2414 3522 2415
rect 3532 2414 3533 2415
rect 3523 2416 3524 2417
rect 3664 2416 3665 2417
rect 3524 2418 3525 2419
rect 3535 2418 3536 2419
rect 3376 2420 3377 2421
rect 3536 2420 3537 2421
rect 3377 2422 3378 2423
rect 3427 2422 3428 2423
rect 3533 2422 3534 2423
rect 3629 2422 3630 2423
rect 3558 2424 3559 2425
rect 3617 2424 3618 2425
rect 3314 2426 3315 2427
rect 3558 2426 3559 2427
rect 3564 2426 3565 2427
rect 3614 2426 3615 2427
rect 3571 2428 3572 2429
rect 3674 2428 3675 2429
rect 3488 2430 3489 2431
rect 3673 2430 3674 2431
rect 3573 2432 3574 2433
rect 3663 2432 3664 2433
rect 3603 2434 3604 2435
rect 3620 2434 3621 2435
rect 3602 2436 3603 2437
rect 3654 2436 3655 2437
rect 3606 2438 3607 2439
rect 3623 2438 3624 2439
rect 3591 2440 3592 2441
rect 3605 2440 3606 2441
rect 3609 2440 3610 2441
rect 3625 2440 3626 2441
rect 3608 2442 3609 2443
rect 3651 2442 3652 2443
rect 3425 2444 3426 2445
rect 3650 2444 3651 2445
rect 3612 2446 3613 2447
rect 3657 2446 3658 2447
rect 3611 2448 3612 2449
rect 3626 2448 3627 2449
rect 3636 2448 3637 2449
rect 3670 2448 3671 2449
rect 3308 2450 3309 2451
rect 3636 2450 3637 2451
rect 3648 2450 3649 2451
rect 3653 2450 3654 2451
rect 3413 2452 3414 2453
rect 3647 2452 3648 2453
rect 2894 2461 2895 2462
rect 3106 2461 3107 2462
rect 2899 2463 2900 2464
rect 2933 2463 2934 2464
rect 2901 2465 2902 2466
rect 3278 2465 3279 2466
rect 2904 2467 2905 2468
rect 3109 2467 3110 2468
rect 2906 2469 2907 2470
rect 3230 2469 3231 2470
rect 2913 2471 2914 2472
rect 3058 2471 3059 2472
rect 2916 2473 2917 2474
rect 3073 2473 3074 2474
rect 2918 2475 2919 2476
rect 3076 2475 3077 2476
rect 2934 2477 2935 2478
rect 3046 2477 3047 2478
rect 2943 2479 2944 2480
rect 3242 2479 3243 2480
rect 2951 2481 2952 2482
rect 2988 2481 2989 2482
rect 2955 2483 2956 2484
rect 3028 2483 3029 2484
rect 2992 2485 2993 2486
rect 3116 2485 3117 2486
rect 2995 2487 2996 2488
rect 3323 2487 3324 2488
rect 3010 2489 3011 2490
rect 3293 2489 3294 2490
rect 3013 2491 3014 2492
rect 3179 2491 3180 2492
rect 3016 2493 3017 2494
rect 3076 2493 3077 2494
rect 3019 2495 3020 2496
rect 3034 2495 3035 2496
rect 3022 2497 3023 2498
rect 3254 2497 3255 2498
rect 3037 2499 3038 2500
rect 3070 2499 3071 2500
rect 3043 2501 3044 2502
rect 3079 2501 3080 2502
rect 3052 2503 3053 2504
rect 3118 2503 3119 2504
rect 3061 2505 3062 2506
rect 3064 2505 3065 2506
rect 2974 2507 2975 2508
rect 3061 2507 3062 2508
rect 3095 2507 3096 2508
rect 3130 2507 3131 2508
rect 3094 2509 3095 2510
rect 3392 2509 3393 2510
rect 3101 2511 3102 2512
rect 3227 2511 3228 2512
rect 3104 2513 3105 2514
rect 3164 2513 3165 2514
rect 3049 2515 3050 2516
rect 3103 2515 3104 2516
rect 3128 2515 3129 2516
rect 3194 2515 3195 2516
rect 3092 2517 3093 2518
rect 3127 2517 3128 2518
rect 3146 2517 3147 2518
rect 3206 2517 3207 2518
rect 3152 2519 3153 2520
rect 3236 2519 3237 2520
rect 3091 2521 3092 2522
rect 3236 2521 3237 2522
rect 3158 2523 3159 2524
rect 3212 2523 3213 2524
rect 3161 2525 3162 2526
rect 3224 2525 3225 2526
rect 3170 2527 3171 2528
rect 3200 2527 3201 2528
rect 3140 2529 3141 2530
rect 3200 2529 3201 2530
rect 3140 2531 3141 2532
rect 3362 2531 3363 2532
rect 3188 2533 3189 2534
rect 3305 2533 3306 2534
rect 3212 2535 3213 2536
rect 3272 2535 3273 2536
rect 3197 2537 3198 2538
rect 3272 2537 3273 2538
rect 3182 2539 3183 2540
rect 3197 2539 3198 2540
rect 3233 2539 3234 2540
rect 3576 2539 3577 2540
rect 2964 2541 2965 2542
rect 3233 2541 3234 2542
rect 3248 2541 3249 2542
rect 3260 2541 3261 2542
rect 3266 2541 3267 2542
rect 3287 2541 3288 2542
rect 3281 2543 3282 2544
rect 3344 2543 3345 2544
rect 2927 2545 2928 2546
rect 3281 2545 3282 2546
rect 3284 2545 3285 2546
rect 3347 2545 3348 2546
rect 3203 2547 3204 2548
rect 3284 2547 3285 2548
rect 3143 2549 3144 2550
rect 3203 2549 3204 2550
rect 3143 2551 3144 2552
rect 3251 2551 3252 2552
rect 3296 2551 3297 2552
rect 3555 2551 3556 2552
rect 3215 2553 3216 2554
rect 3296 2553 3297 2554
rect 3302 2553 3303 2554
rect 3368 2553 3369 2554
rect 3086 2555 3087 2556
rect 3302 2555 3303 2556
rect 3067 2557 3068 2558
rect 3085 2557 3086 2558
rect 3308 2557 3309 2558
rect 3374 2557 3375 2558
rect 3257 2559 3258 2560
rect 3308 2559 3309 2560
rect 3314 2559 3315 2560
rect 3386 2559 3387 2560
rect 3239 2561 3240 2562
rect 3314 2561 3315 2562
rect 3320 2561 3321 2562
rect 3380 2561 3381 2562
rect 3245 2563 3246 2564
rect 3320 2563 3321 2564
rect 3031 2565 3032 2566
rect 3245 2565 3246 2566
rect 3326 2565 3327 2566
rect 3392 2565 3393 2566
rect 2985 2567 2986 2568
rect 3326 2567 3327 2568
rect 2961 2569 2962 2570
rect 2986 2569 2987 2570
rect 3332 2569 3333 2570
rect 3398 2569 3399 2570
rect 3290 2571 3291 2572
rect 3332 2571 3333 2572
rect 3209 2573 3210 2574
rect 3290 2573 3291 2574
rect 3004 2575 3005 2576
rect 3209 2575 3210 2576
rect 3004 2577 3005 2578
rect 3040 2577 3041 2578
rect 3338 2577 3339 2578
rect 3410 2577 3411 2578
rect 3263 2579 3264 2580
rect 3338 2579 3339 2580
rect 3350 2579 3351 2580
rect 3692 2579 3693 2580
rect 3275 2581 3276 2582
rect 3350 2581 3351 2582
rect 2915 2583 2916 2584
rect 3275 2583 3276 2584
rect 3353 2583 3354 2584
rect 3482 2583 3483 2584
rect 3356 2585 3357 2586
rect 3551 2585 3552 2586
rect 3365 2587 3366 2588
rect 3431 2587 3432 2588
rect 3371 2589 3372 2590
rect 3443 2589 3444 2590
rect 3176 2591 3177 2592
rect 3371 2591 3372 2592
rect 3122 2593 3123 2594
rect 3176 2593 3177 2594
rect 2979 2595 2980 2596
rect 3121 2595 3122 2596
rect 3401 2595 3402 2596
rect 3467 2595 3468 2596
rect 3416 2597 3417 2598
rect 3419 2597 3420 2598
rect 3422 2597 3423 2598
rect 3661 2597 3662 2598
rect 3425 2599 3426 2600
rect 3667 2599 3668 2600
rect 3359 2601 3360 2602
rect 3425 2601 3426 2602
rect 3452 2601 3453 2602
rect 3593 2601 3594 2602
rect 3458 2603 3459 2604
rect 3506 2603 3507 2604
rect 3479 2605 3480 2606
rect 3515 2605 3516 2606
rect 3449 2607 3450 2608
rect 3479 2607 3480 2608
rect 3485 2607 3486 2608
rect 3551 2607 3552 2608
rect 3413 2609 3414 2610
rect 3485 2609 3486 2610
rect 3488 2609 3489 2610
rect 3554 2609 3555 2610
rect 3497 2611 3498 2612
rect 3611 2611 3612 2612
rect 3500 2613 3501 2614
rect 3608 2613 3609 2614
rect 3509 2615 3510 2616
rect 3557 2615 3558 2616
rect 3437 2617 3438 2618
rect 3509 2617 3510 2618
rect 3521 2617 3522 2618
rect 3578 2617 3579 2618
rect 3524 2619 3525 2620
rect 3581 2619 3582 2620
rect 3527 2621 3528 2622
rect 3563 2621 3564 2622
rect 3533 2623 3534 2624
rect 3656 2623 3657 2624
rect 3545 2625 3546 2626
rect 3567 2625 3568 2626
rect 3503 2627 3504 2628
rect 3545 2627 3546 2628
rect 3455 2629 3456 2630
rect 3503 2629 3504 2630
rect 3383 2631 3384 2632
rect 3455 2631 3456 2632
rect 3530 2631 3531 2632
rect 3566 2631 3567 2632
rect 3569 2631 3570 2632
rect 3586 2631 3587 2632
rect 3536 2633 3537 2634
rect 3587 2633 3588 2634
rect 3573 2635 3574 2636
rect 3637 2635 3638 2636
rect 3377 2637 3378 2638
rect 3572 2637 3573 2638
rect 3311 2639 3312 2640
rect 3377 2639 3378 2640
rect 3575 2639 3576 2640
rect 3743 2639 3744 2640
rect 3584 2641 3585 2642
rect 3590 2641 3591 2642
rect 3539 2643 3540 2644
rect 3590 2643 3591 2644
rect 3473 2645 3474 2646
rect 3539 2645 3540 2646
rect 3599 2645 3600 2646
rect 3650 2645 3651 2646
rect 3605 2647 3606 2648
rect 3655 2647 3656 2648
rect 3329 2649 3330 2650
rect 3605 2649 3606 2650
rect 3617 2649 3618 2650
rect 3679 2649 3680 2650
rect 3404 2651 3405 2652
rect 3617 2651 3618 2652
rect 3620 2651 3621 2652
rect 3664 2651 3665 2652
rect 3623 2653 3624 2654
rect 3647 2653 3648 2654
rect 3542 2655 3543 2656
rect 3624 2655 3625 2656
rect 3476 2657 3477 2658
rect 3542 2657 3543 2658
rect 3653 2657 3654 2658
rect 3695 2657 3696 2658
rect 3602 2659 3603 2660
rect 3652 2659 3653 2660
rect 3602 2661 3603 2662
rect 3640 2661 3641 2662
rect 3670 2661 3671 2662
rect 3689 2661 3690 2662
rect 3677 2663 3678 2664
rect 3733 2663 3734 2664
rect 3614 2665 3615 2666
rect 3676 2665 3677 2666
rect 2890 2674 2891 2675
rect 3200 2674 3201 2675
rect 2897 2676 2898 2677
rect 3109 2676 3110 2677
rect 2905 2678 2906 2679
rect 3133 2678 3134 2679
rect 2915 2680 2916 2681
rect 3006 2680 3007 2681
rect 2931 2682 2932 2683
rect 3070 2682 3071 2683
rect 2934 2684 2935 2685
rect 3281 2684 3282 2685
rect 2908 2686 2909 2687
rect 3280 2686 3281 2687
rect 2937 2688 2938 2689
rect 2967 2688 2968 2689
rect 2941 2690 2942 2691
rect 3206 2690 3207 2691
rect 2944 2692 2945 2693
rect 3268 2692 3269 2693
rect 2943 2694 2944 2695
rect 2948 2694 2949 2695
rect 2946 2696 2947 2697
rect 3209 2696 3210 2697
rect 2965 2698 2966 2699
rect 3433 2698 3434 2699
rect 2974 2700 2975 2701
rect 3197 2700 3198 2701
rect 2976 2702 2977 2703
rect 3194 2702 3195 2703
rect 2986 2704 2987 2705
rect 3018 2704 3019 2705
rect 2997 2706 2998 2707
rect 3212 2706 3213 2707
rect 3004 2708 3005 2709
rect 3358 2708 3359 2709
rect 3028 2710 3029 2711
rect 3055 2710 3056 2711
rect 3027 2712 3028 2713
rect 3158 2712 3159 2713
rect 3034 2714 3035 2715
rect 3049 2714 3050 2715
rect 3036 2716 3037 2717
rect 3064 2716 3065 2717
rect 3046 2718 3047 2719
rect 3302 2718 3303 2719
rect 3061 2720 3062 2721
rect 3088 2720 3089 2721
rect 3073 2722 3074 2723
rect 3245 2722 3246 2723
rect 3076 2724 3077 2725
rect 3112 2724 3113 2725
rect 3079 2726 3080 2727
rect 3097 2726 3098 2727
rect 3079 2728 3080 2729
rect 3109 2728 3110 2729
rect 3082 2730 3083 2731
rect 3314 2730 3315 2731
rect 3085 2732 3086 2733
rect 3091 2732 3092 2733
rect 3058 2734 3059 2735
rect 3085 2734 3086 2735
rect 3094 2734 3095 2735
rect 3136 2734 3137 2735
rect 3103 2736 3104 2737
rect 3148 2736 3149 2737
rect 3103 2738 3104 2739
rect 3460 2738 3461 2739
rect 3106 2740 3107 2741
rect 3121 2740 3122 2741
rect 3106 2742 3107 2743
rect 3266 2742 3267 2743
rect 3115 2744 3116 2745
rect 3127 2744 3128 2745
rect 3124 2746 3125 2747
rect 3308 2746 3309 2747
rect 3140 2748 3141 2749
rect 3617 2748 3618 2749
rect 3151 2750 3152 2751
rect 3188 2750 3189 2751
rect 3022 2752 3023 2753
rect 3187 2752 3188 2753
rect 3164 2754 3165 2755
rect 3181 2754 3182 2755
rect 3170 2756 3171 2757
rect 3205 2756 3206 2757
rect 3176 2758 3177 2759
rect 3193 2758 3194 2759
rect 3199 2758 3200 2759
rect 3566 2758 3567 2759
rect 3217 2760 3218 2761
rect 3254 2760 3255 2761
rect 3224 2762 3225 2763
rect 3244 2762 3245 2763
rect 2979 2764 2980 2765
rect 3223 2764 3224 2765
rect 3230 2764 3231 2765
rect 3298 2764 3299 2765
rect 3229 2766 3230 2767
rect 3515 2766 3516 2767
rect 3233 2768 3234 2769
rect 3301 2768 3302 2769
rect 3236 2770 3237 2771
rect 3250 2770 3251 2771
rect 3203 2772 3204 2773
rect 3235 2772 3236 2773
rect 3238 2772 3239 2773
rect 3590 2772 3591 2773
rect 3242 2774 3243 2775
rect 3286 2774 3287 2775
rect 3256 2776 3257 2777
rect 3326 2776 3327 2777
rect 3262 2778 3263 2779
rect 3404 2778 3405 2779
rect 3275 2780 3276 2781
rect 3325 2780 3326 2781
rect 3260 2782 3261 2783
rect 3274 2782 3275 2783
rect 3259 2784 3260 2785
rect 3329 2784 3330 2785
rect 2969 2786 2970 2787
rect 3328 2786 3329 2787
rect 3284 2788 3285 2789
rect 3316 2788 3317 2789
rect 3293 2790 3294 2791
rect 3334 2790 3335 2791
rect 3292 2792 3293 2793
rect 3587 2792 3588 2793
rect 3296 2794 3297 2795
rect 3310 2794 3311 2795
rect 3323 2794 3324 2795
rect 3394 2794 3395 2795
rect 3272 2796 3273 2797
rect 3322 2796 3323 2797
rect 3332 2796 3333 2797
rect 3620 2796 3621 2797
rect 3290 2798 3291 2799
rect 3331 2798 3332 2799
rect 2915 2800 2916 2801
rect 3289 2800 3290 2801
rect 3344 2800 3345 2801
rect 3427 2800 3428 2801
rect 3356 2802 3357 2803
rect 3687 2802 3688 2803
rect 3278 2804 3279 2805
rect 3355 2804 3356 2805
rect 3368 2804 3369 2805
rect 3451 2804 3452 2805
rect 3367 2806 3368 2807
rect 3661 2806 3662 2807
rect 3374 2808 3375 2809
rect 3463 2808 3464 2809
rect 3362 2810 3363 2811
rect 3373 2810 3374 2811
rect 3380 2810 3381 2811
rect 3403 2810 3404 2811
rect 2950 2812 2951 2813
rect 3379 2812 3380 2813
rect 3386 2812 3387 2813
rect 3457 2812 3458 2813
rect 3160 2814 3161 2815
rect 3385 2814 3386 2815
rect 3398 2814 3399 2815
rect 3487 2814 3488 2815
rect 3397 2816 3398 2817
rect 3605 2816 3606 2817
rect 3410 2818 3411 2819
rect 3662 2818 3663 2819
rect 3409 2820 3410 2821
rect 3754 2820 3755 2821
rect 3425 2822 3426 2823
rect 3517 2822 3518 2823
rect 3431 2824 3432 2825
rect 3523 2824 3524 2825
rect 3347 2826 3348 2827
rect 3430 2826 3431 2827
rect 3439 2826 3440 2827
rect 3672 2826 3673 2827
rect 3443 2828 3444 2829
rect 3493 2828 3494 2829
rect 2972 2830 2973 2831
rect 3442 2830 3443 2831
rect 3455 2830 3456 2831
rect 3547 2830 3548 2831
rect 3371 2832 3372 2833
rect 3454 2832 3455 2833
rect 3467 2832 3468 2833
rect 3559 2832 3560 2833
rect 3377 2834 3378 2835
rect 3466 2834 3467 2835
rect 3475 2834 3476 2835
rect 3624 2834 3625 2835
rect 3479 2836 3480 2837
rect 3691 2836 3692 2837
rect 3482 2838 3483 2839
rect 3658 2838 3659 2839
rect 3392 2840 3393 2841
rect 3481 2840 3482 2841
rect 3320 2842 3321 2843
rect 3391 2842 3392 2843
rect 3415 2842 3416 2843
rect 3658 2842 3659 2843
rect 3490 2844 3491 2845
rect 3563 2844 3564 2845
rect 3496 2846 3497 2847
rect 3503 2846 3504 2847
rect 3499 2848 3500 2849
rect 3557 2848 3558 2849
rect 3506 2850 3507 2851
rect 3640 2850 3641 2851
rect 3505 2852 3506 2853
rect 3631 2852 3632 2853
rect 3509 2854 3510 2855
rect 3595 2854 3596 2855
rect 3422 2856 3423 2857
rect 3508 2856 3509 2857
rect 3350 2858 3351 2859
rect 3421 2858 3422 2859
rect 2922 2860 2923 2861
rect 3349 2860 3350 2861
rect 3526 2860 3527 2861
rect 3684 2860 3685 2861
rect 3529 2862 3530 2863
rect 3572 2862 3573 2863
rect 3485 2864 3486 2865
rect 3571 2864 3572 2865
rect 3532 2866 3533 2867
rect 3569 2866 3570 2867
rect 3535 2868 3536 2869
rect 3545 2868 3546 2869
rect 3539 2870 3540 2871
rect 3607 2870 3608 2871
rect 3542 2872 3543 2873
rect 3610 2872 3611 2873
rect 3541 2874 3542 2875
rect 3682 2874 3683 2875
rect 3551 2876 3552 2877
rect 3625 2876 3626 2877
rect 3554 2878 3555 2879
rect 3628 2878 3629 2879
rect 3565 2880 3566 2881
rect 3581 2880 3582 2881
rect 3575 2882 3576 2883
rect 3768 2882 3769 2883
rect 3578 2884 3579 2885
rect 3640 2884 3641 2885
rect 3589 2886 3590 2887
rect 3599 2886 3600 2887
rect 3592 2888 3593 2889
rect 3602 2888 3603 2889
rect 3652 2888 3653 2889
rect 3681 2888 3682 2889
rect 3655 2890 3656 2891
rect 3718 2890 3719 2891
rect 3338 2892 3339 2893
rect 3655 2892 3656 2893
rect 3039 2894 3040 2895
rect 3337 2894 3338 2895
rect 3676 2894 3677 2895
rect 3712 2894 3713 2895
rect 3679 2896 3680 2897
rect 3715 2896 3716 2897
rect 3584 2898 3585 2899
rect 3678 2898 3679 2899
rect 3583 2900 3584 2901
rect 3667 2900 3668 2901
rect 3689 2900 3690 2901
rect 3758 2900 3759 2901
rect 3695 2902 3696 2903
rect 3738 2902 3739 2903
rect 3708 2904 3709 2905
rect 3726 2904 3727 2905
rect 3637 2906 3638 2907
rect 3709 2906 3710 2907
rect 3637 2908 3638 2909
rect 3698 2908 3699 2909
rect 3664 2910 3665 2911
rect 3697 2910 3698 2911
rect 3361 2912 3362 2913
rect 3665 2912 3666 2913
rect 3729 2912 3730 2913
rect 3736 2912 3737 2913
rect 3601 2914 3602 2915
rect 3735 2914 3736 2915
rect 3675 2916 3676 2917
rect 3728 2916 3729 2917
rect 3733 2916 3734 2917
rect 3786 2916 3787 2917
rect 3740 2918 3741 2919
rect 3747 2918 3748 2919
rect 3700 2920 3701 2921
rect 3747 2920 3748 2921
rect 3741 2922 3742 2923
rect 3772 2922 3773 2923
rect 2914 2931 2915 2932
rect 3085 2931 3086 2932
rect 2931 2933 2932 2934
rect 3286 2933 3287 2934
rect 2950 2935 2951 2936
rect 3363 2935 3364 2936
rect 2953 2937 2954 2938
rect 3358 2937 3359 2938
rect 2962 2939 2963 2940
rect 3073 2939 3074 2940
rect 2934 2941 2935 2942
rect 3072 2941 3073 2942
rect 2921 2943 2922 2944
rect 2933 2943 2934 2944
rect 2961 2943 2962 2944
rect 2994 2943 2995 2944
rect 2971 2945 2972 2946
rect 3427 2945 3428 2946
rect 2976 2947 2977 2948
rect 3193 2947 3194 2948
rect 2993 2949 2994 2950
rect 3468 2949 3469 2950
rect 3006 2951 3007 2952
rect 3029 2951 3030 2952
rect 3014 2953 3015 2954
rect 3244 2953 3245 2954
rect 3018 2955 3019 2956
rect 3023 2955 3024 2956
rect 3027 2955 3028 2956
rect 3187 2955 3188 2956
rect 3043 2957 3044 2958
rect 3421 2957 3422 2958
rect 3045 2959 3046 2960
rect 3162 2959 3163 2960
rect 3055 2961 3056 2962
rect 3060 2961 3061 2962
rect 3069 2961 3070 2962
rect 3103 2961 3104 2962
rect 3079 2963 3080 2964
rect 3303 2963 3304 2964
rect 2979 2965 2980 2966
rect 3078 2965 3079 2966
rect 2978 2967 2979 2968
rect 3379 2967 3380 2968
rect 3097 2969 3098 2970
rect 3099 2969 3100 2970
rect 3096 2971 3097 2972
rect 3112 2971 3113 2972
rect 3091 2973 3092 2974
rect 3111 2973 3112 2974
rect 3106 2975 3107 2976
rect 3259 2975 3260 2976
rect 3109 2977 3110 2978
rect 3123 2977 3124 2978
rect 3115 2979 3116 2980
rect 3144 2979 3145 2980
rect 3126 2981 3127 2982
rect 3148 2981 3149 2982
rect 3118 2983 3119 2984
rect 3147 2983 3148 2984
rect 3117 2985 3118 2986
rect 3475 2985 3476 2986
rect 3130 2987 3131 2988
rect 3138 2987 3139 2988
rect 3121 2989 3122 2990
rect 3129 2989 3130 2990
rect 3120 2991 3121 2992
rect 3378 2991 3379 2992
rect 3133 2993 3134 2994
rect 3141 2993 3142 2994
rect 3151 2993 3152 2994
rect 3174 2993 3175 2994
rect 3157 2995 3158 2996
rect 3238 2995 3239 2996
rect 3160 2997 3161 2998
rect 3373 2997 3374 2998
rect 3181 2999 3182 3000
rect 3186 2999 3187 3000
rect 3180 3001 3181 3002
rect 3442 3001 3443 3002
rect 3210 3003 3211 3004
rect 3223 3003 3224 3004
rect 3222 3005 3223 3006
rect 3229 3005 3230 3006
rect 3228 3007 3229 3008
rect 3250 3007 3251 3008
rect 2899 3009 2900 3010
rect 3249 3009 3250 3010
rect 3237 3011 3238 3012
rect 3765 3011 3766 3012
rect 3240 3013 3241 3014
rect 3262 3013 3263 3014
rect 3246 3015 3247 3016
rect 3256 3015 3257 3016
rect 3255 3017 3256 3018
rect 3274 3017 3275 3018
rect 3261 3019 3262 3020
rect 3658 3019 3659 3020
rect 3268 3021 3269 3022
rect 3273 3021 3274 3022
rect 3267 3023 3268 3024
rect 3310 3023 3311 3024
rect 3038 3025 3039 3026
rect 3309 3025 3310 3026
rect 3280 3027 3281 3028
rect 3285 3027 3286 3028
rect 3279 3029 3280 3030
rect 3316 3029 3317 3030
rect 3292 3031 3293 3032
rect 3357 3031 3358 3032
rect 3291 3033 3292 3034
rect 3298 3033 3299 3034
rect 2975 3035 2976 3036
rect 3297 3035 3298 3036
rect 3294 3037 3295 3038
rect 3301 3037 3302 3038
rect 3312 3037 3313 3038
rect 3430 3037 3431 3038
rect 3315 3039 3316 3040
rect 3331 3039 3332 3040
rect 3318 3041 3319 3042
rect 3334 3041 3335 3042
rect 3325 3043 3326 3044
rect 3369 3043 3370 3044
rect 2943 3045 2944 3046
rect 3324 3045 3325 3046
rect 3333 3045 3334 3046
rect 3337 3045 3338 3046
rect 3349 3045 3350 3046
rect 3351 3045 3352 3046
rect 3372 3045 3373 3046
rect 3685 3045 3686 3046
rect 3403 3047 3404 3048
rect 3660 3047 3661 3048
rect 3397 3049 3398 3050
rect 3402 3049 3403 3050
rect 2912 3051 2913 3052
rect 3396 3051 3397 3052
rect 2911 3053 2912 3054
rect 3084 3053 3085 3054
rect 3409 3053 3410 3054
rect 3420 3053 3421 3054
rect 3367 3055 3368 3056
rect 3408 3055 3409 3056
rect 2965 3057 2966 3058
rect 3366 3057 3367 3058
rect 2964 3059 2965 3060
rect 3205 3059 3206 3060
rect 3415 3059 3416 3060
rect 3426 3059 3427 3060
rect 3439 3059 3440 3060
rect 3444 3059 3445 3060
rect 3361 3061 3362 3062
rect 3438 3061 3439 3062
rect 3454 3061 3455 3062
rect 3483 3061 3484 3062
rect 2946 3063 2947 3064
rect 3453 3063 3454 3064
rect 3466 3063 3467 3064
rect 3471 3063 3472 3064
rect 3460 3065 3461 3066
rect 3465 3065 3466 3066
rect 3499 3065 3500 3066
rect 3756 3065 3757 3066
rect 3505 3067 3506 3068
rect 3510 3067 3511 3068
rect 3493 3069 3494 3070
rect 3504 3069 3505 3070
rect 3487 3071 3488 3072
rect 3492 3071 3493 3072
rect 3481 3073 3482 3074
rect 3486 3073 3487 3074
rect 3082 3075 3083 3076
rect 3480 3075 3481 3076
rect 3508 3075 3509 3076
rect 3513 3075 3514 3076
rect 3496 3077 3497 3078
rect 3507 3077 3508 3078
rect 3490 3079 3491 3080
rect 3495 3079 3496 3080
rect 3535 3079 3536 3080
rect 3728 3079 3729 3080
rect 3523 3081 3524 3082
rect 3534 3081 3535 3082
rect 3517 3083 3518 3084
rect 3522 3083 3523 3084
rect 3433 3085 3434 3086
rect 3516 3085 3517 3086
rect 3432 3087 3433 3088
rect 3451 3087 3452 3088
rect 3450 3089 3451 3090
rect 3669 3089 3670 3090
rect 3541 3091 3542 3092
rect 3687 3091 3688 3092
rect 3526 3093 3527 3094
rect 3540 3093 3541 3094
rect 3543 3093 3544 3094
rect 3691 3093 3692 3094
rect 3585 3095 3586 3096
rect 3703 3095 3704 3096
rect 3589 3097 3590 3098
rect 3621 3097 3622 3098
rect 3571 3099 3572 3100
rect 3588 3099 3589 3100
rect 3559 3101 3560 3102
rect 3570 3101 3571 3102
rect 3547 3103 3548 3104
rect 3558 3103 3559 3104
rect 3529 3105 3530 3106
rect 3546 3105 3547 3106
rect 3528 3107 3529 3108
rect 3727 3107 3728 3108
rect 3595 3109 3596 3110
rect 3615 3109 3616 3110
rect 3610 3111 3611 3112
rect 3630 3111 3631 3112
rect 3612 3113 3613 3114
rect 3796 3113 3797 3114
rect 3625 3115 3626 3116
rect 3791 3115 3792 3116
rect 3592 3117 3593 3118
rect 3624 3117 3625 3118
rect 3628 3117 3629 3118
rect 3793 3117 3794 3118
rect 3607 3119 3608 3120
rect 3627 3119 3628 3120
rect 3565 3121 3566 3122
rect 3606 3121 3607 3122
rect 3637 3121 3638 3122
rect 3746 3121 3747 3122
rect 3640 3123 3641 3124
rect 3645 3123 3646 3124
rect 3657 3123 3658 3124
rect 3749 3123 3750 3124
rect 3669 3125 3670 3126
rect 3779 3125 3780 3126
rect 3601 3127 3602 3128
rect 3778 3127 3779 3128
rect 3583 3129 3584 3130
rect 3600 3129 3601 3130
rect 3532 3131 3533 3132
rect 3582 3131 3583 3132
rect 3678 3131 3679 3132
rect 3718 3131 3719 3132
rect 3681 3133 3682 3134
rect 3703 3133 3704 3134
rect 3700 3135 3701 3136
rect 3718 3135 3719 3136
rect 3694 3137 3695 3138
rect 3700 3137 3701 3138
rect 3706 3137 3707 3138
rect 3794 3137 3795 3138
rect 3709 3139 3710 3140
rect 3721 3139 3722 3140
rect 3738 3139 3739 3140
rect 3762 3139 3763 3140
rect 3712 3141 3713 3142
rect 3737 3141 3738 3142
rect 3741 3141 3742 3142
rect 3765 3141 3766 3142
rect 3715 3143 3716 3144
rect 3740 3143 3741 3144
rect 3697 3145 3698 3146
rect 3715 3145 3716 3146
rect 3675 3147 3676 3148
rect 3697 3147 3698 3148
rect 3772 3147 3773 3148
rect 3789 3147 3790 3148
rect 3743 3149 3744 3150
rect 3771 3149 3772 3150
rect 3788 3149 3789 3150
rect 3808 3149 3809 3150
rect 3797 3151 3798 3152
rect 3801 3151 3802 3152
rect 3824 3151 3825 3152
rect 3831 3151 3832 3152
rect 2906 3160 2907 3161
rect 3069 3160 3070 3161
rect 2909 3162 2910 3163
rect 3129 3162 3130 3163
rect 2913 3164 2914 3165
rect 3141 3164 3142 3165
rect 2916 3166 2917 3167
rect 3075 3166 3076 3167
rect 2933 3168 2934 3169
rect 2949 3168 2950 3169
rect 2935 3170 2936 3171
rect 3258 3170 3259 3171
rect 2945 3172 2946 3173
rect 3029 3172 3030 3173
rect 2944 3174 2945 3175
rect 3321 3174 3322 3175
rect 2951 3176 2952 3177
rect 3363 3176 3364 3177
rect 2958 3178 2959 3179
rect 3369 3178 3370 3179
rect 2961 3180 2962 3181
rect 3312 3180 3313 3181
rect 2968 3182 2969 3183
rect 2980 3182 2981 3183
rect 2968 3184 2969 3185
rect 3309 3184 3310 3185
rect 2977 3186 2978 3187
rect 3501 3186 3502 3187
rect 2984 3188 2985 3189
rect 3156 3188 3157 3189
rect 2987 3190 2988 3191
rect 3144 3190 3145 3191
rect 2993 3192 2994 3193
rect 3002 3192 3003 3193
rect 3014 3192 3015 3193
rect 3105 3192 3106 3193
rect 3014 3194 3015 3195
rect 3023 3194 3024 3195
rect 3020 3196 3021 3197
rect 3306 3196 3307 3197
rect 3023 3198 3024 3199
rect 3414 3198 3415 3199
rect 3030 3200 3031 3201
rect 3468 3200 3469 3201
rect 3033 3202 3034 3203
rect 3048 3202 3049 3203
rect 3042 3204 3043 3205
rect 3168 3204 3169 3205
rect 3045 3206 3046 3207
rect 3471 3206 3472 3207
rect 3051 3208 3052 3209
rect 3060 3208 3061 3209
rect 3057 3210 3058 3211
rect 3727 3210 3728 3211
rect 3063 3212 3064 3213
rect 3072 3212 3073 3213
rect 3078 3212 3079 3213
rect 3339 3212 3340 3213
rect 3084 3214 3085 3215
rect 3102 3214 3103 3215
rect 3087 3216 3088 3217
rect 3105 3216 3106 3217
rect 3093 3218 3094 3219
rect 3096 3218 3097 3219
rect 2911 3220 2912 3221
rect 3096 3220 3097 3221
rect 3099 3220 3100 3221
rect 3114 3220 3115 3221
rect 3108 3222 3109 3223
rect 3117 3222 3118 3223
rect 3111 3224 3112 3225
rect 3129 3224 3130 3225
rect 3123 3226 3124 3227
rect 3165 3226 3166 3227
rect 3123 3228 3124 3229
rect 3150 3228 3151 3229
rect 3138 3230 3139 3231
rect 3141 3230 3142 3231
rect 3174 3230 3175 3231
rect 3429 3230 3430 3231
rect 3162 3232 3163 3233
rect 3174 3232 3175 3233
rect 3066 3234 3067 3235
rect 3162 3234 3163 3235
rect 3201 3234 3202 3235
rect 3276 3234 3277 3235
rect 3207 3236 3208 3237
rect 3324 3236 3325 3237
rect 3213 3238 3214 3239
rect 3237 3238 3238 3239
rect 3147 3240 3148 3241
rect 3237 3240 3238 3241
rect 3222 3242 3223 3243
rect 3633 3242 3634 3243
rect 3243 3244 3244 3245
rect 3294 3244 3295 3245
rect 3255 3246 3256 3247
rect 3300 3246 3301 3247
rect 3264 3248 3265 3249
rect 3285 3248 3286 3249
rect 3267 3250 3268 3251
rect 3342 3250 3343 3251
rect 3270 3252 3271 3253
rect 3273 3252 3274 3253
rect 3273 3254 3274 3255
rect 3288 3254 3289 3255
rect 3282 3256 3283 3257
rect 3354 3256 3355 3257
rect 3288 3258 3289 3259
rect 3351 3258 3352 3259
rect 3294 3260 3295 3261
rect 3327 3260 3328 3261
rect 3297 3262 3298 3263
rect 3336 3262 3337 3263
rect 3303 3264 3304 3265
rect 3330 3264 3331 3265
rect 3312 3266 3313 3267
rect 3366 3266 3367 3267
rect 3279 3268 3280 3269
rect 3366 3268 3367 3269
rect 3318 3270 3319 3271
rect 3381 3270 3382 3271
rect 3120 3272 3121 3273
rect 3318 3272 3319 3273
rect 3120 3274 3121 3275
rect 3126 3274 3127 3275
rect 3324 3274 3325 3275
rect 3396 3274 3397 3275
rect 3252 3276 3253 3277
rect 3396 3276 3397 3277
rect 3348 3278 3349 3279
rect 3444 3278 3445 3279
rect 3354 3280 3355 3281
rect 3450 3280 3451 3281
rect 3360 3282 3361 3283
rect 3390 3282 3391 3283
rect 3372 3284 3373 3285
rect 3756 3284 3757 3285
rect 3372 3286 3373 3287
rect 3456 3286 3457 3287
rect 3375 3288 3376 3289
rect 3712 3288 3713 3289
rect 3378 3290 3379 3291
rect 3660 3290 3661 3291
rect 3315 3292 3316 3293
rect 3378 3292 3379 3293
rect 2961 3294 2962 3295
rect 3315 3294 3316 3295
rect 3390 3294 3391 3295
rect 3480 3294 3481 3295
rect 3393 3296 3394 3297
rect 3423 3296 3424 3297
rect 3402 3298 3403 3299
rect 3688 3298 3689 3299
rect 3402 3300 3403 3301
rect 3486 3300 3487 3301
rect 3408 3302 3409 3303
rect 3657 3302 3658 3303
rect 3333 3304 3334 3305
rect 3408 3304 3409 3305
rect 3426 3304 3427 3305
rect 3681 3304 3682 3305
rect 3027 3306 3028 3307
rect 3426 3306 3427 3307
rect 3435 3306 3436 3307
rect 3528 3306 3529 3307
rect 3441 3308 3442 3309
rect 3462 3308 3463 3309
rect 3459 3310 3460 3311
rect 3534 3310 3535 3311
rect 3240 3312 3241 3313
rect 3534 3312 3535 3313
rect 3240 3314 3241 3315
rect 3291 3314 3292 3315
rect 2921 3316 2922 3317
rect 3291 3316 3292 3317
rect 2920 3318 2921 3319
rect 3483 3318 3484 3319
rect 3471 3320 3472 3321
rect 3540 3320 3541 3321
rect 3477 3322 3478 3323
rect 3797 3322 3798 3323
rect 3483 3324 3484 3325
rect 3706 3324 3707 3325
rect 3489 3326 3490 3327
rect 3570 3326 3571 3327
rect 3492 3328 3493 3329
rect 3723 3328 3724 3329
rect 3504 3330 3505 3331
rect 3709 3330 3710 3331
rect 3246 3332 3247 3333
rect 3504 3332 3505 3333
rect 3210 3334 3211 3335
rect 3246 3334 3247 3335
rect 3210 3336 3211 3337
rect 3234 3336 3235 3337
rect 3234 3338 3235 3339
rect 3785 3338 3786 3339
rect 3507 3340 3508 3341
rect 3642 3340 3643 3341
rect 3507 3342 3508 3343
rect 3546 3342 3547 3343
rect 3513 3344 3514 3345
rect 3685 3344 3686 3345
rect 3216 3346 3217 3347
rect 3513 3346 3514 3347
rect 3516 3346 3517 3347
rect 3648 3346 3649 3347
rect 3522 3348 3523 3349
rect 3784 3348 3785 3349
rect 3525 3350 3526 3351
rect 3612 3350 3613 3351
rect 3420 3352 3421 3353
rect 3612 3352 3613 3353
rect 3228 3354 3229 3355
rect 3420 3354 3421 3355
rect 3228 3356 3229 3357
rect 3249 3356 3250 3357
rect 3540 3356 3541 3357
rect 3600 3356 3601 3357
rect 3552 3358 3553 3359
rect 3585 3358 3586 3359
rect 3564 3360 3565 3361
rect 3897 3360 3898 3361
rect 3570 3362 3571 3363
rect 3627 3362 3628 3363
rect 3573 3364 3574 3365
rect 3630 3364 3631 3365
rect 3465 3366 3466 3367
rect 3630 3366 3631 3367
rect 3465 3368 3466 3369
rect 3780 3368 3781 3369
rect 3576 3370 3577 3371
rect 3827 3370 3828 3371
rect 3582 3372 3583 3373
rect 3687 3372 3688 3373
rect 3582 3374 3583 3375
rect 3791 3374 3792 3375
rect 3594 3376 3595 3377
rect 3606 3376 3607 3377
rect 3621 3376 3622 3377
rect 3693 3376 3694 3377
rect 3645 3378 3646 3379
rect 3660 3378 3661 3379
rect 3438 3380 3439 3381
rect 3645 3380 3646 3381
rect 3666 3380 3667 3381
rect 3669 3380 3670 3381
rect 3669 3382 3670 3383
rect 3746 3382 3747 3383
rect 3192 3384 3193 3385
rect 3747 3384 3748 3385
rect 3186 3386 3187 3387
rect 3192 3386 3193 3387
rect 3180 3388 3181 3389
rect 3186 3388 3187 3389
rect 2964 3390 2965 3391
rect 3180 3390 3181 3391
rect 2965 3392 2966 3393
rect 3204 3392 3205 3393
rect 3681 3392 3682 3393
rect 3765 3392 3766 3393
rect 3690 3394 3691 3395
rect 3766 3394 3767 3395
rect 3697 3396 3698 3397
rect 3732 3396 3733 3397
rect 3624 3398 3625 3399
rect 3696 3398 3697 3399
rect 3543 3400 3544 3401
rect 3624 3400 3625 3401
rect 3700 3400 3701 3401
rect 3735 3400 3736 3401
rect 3495 3402 3496 3403
rect 3699 3402 3700 3403
rect 3261 3404 3262 3405
rect 3495 3404 3496 3405
rect 3705 3404 3706 3405
rect 3721 3404 3722 3405
rect 3715 3406 3716 3407
rect 3844 3406 3845 3407
rect 3678 3408 3679 3409
rect 3714 3408 3715 3409
rect 3737 3408 3738 3409
rect 3790 3408 3791 3409
rect 3703 3410 3704 3411
rect 3738 3410 3739 3411
rect 3195 3412 3196 3413
rect 3702 3412 3703 3413
rect 3743 3412 3744 3413
rect 3796 3412 3797 3413
rect 3357 3414 3358 3415
rect 3744 3414 3745 3415
rect 3357 3416 3358 3417
rect 3453 3416 3454 3417
rect 3384 3418 3385 3419
rect 3453 3418 3454 3419
rect 3384 3420 3385 3421
rect 3432 3420 3433 3421
rect 3432 3422 3433 3423
rect 3510 3422 3511 3423
rect 3750 3422 3751 3423
rect 3841 3422 3842 3423
rect 3752 3424 3753 3425
rect 3794 3424 3795 3425
rect 3718 3426 3719 3427
rect 3753 3426 3754 3427
rect 3717 3428 3718 3429
rect 3851 3428 3852 3429
rect 3740 3430 3741 3431
rect 3793 3430 3794 3431
rect 3741 3432 3742 3433
rect 3866 3432 3867 3433
rect 3762 3434 3763 3435
rect 3863 3434 3864 3435
rect 3768 3436 3769 3437
rect 3817 3436 3818 3437
rect 3788 3438 3789 3439
rect 3854 3438 3855 3439
rect 3588 3440 3589 3441
rect 3787 3440 3788 3441
rect 3804 3440 3805 3441
rect 3887 3440 3888 3441
rect 3811 3442 3812 3443
rect 3876 3442 3877 3443
rect 3815 3444 3816 3445
rect 3857 3444 3858 3445
rect 3771 3446 3772 3447
rect 3814 3446 3815 3447
rect 3831 3446 3832 3447
rect 3838 3446 3839 3447
rect 3558 3448 3559 3449
rect 3830 3448 3831 3449
rect 3558 3450 3559 3451
rect 3615 3450 3616 3451
rect 3860 3450 3861 3451
rect 3880 3450 3881 3451
rect 2815 3459 2816 3460
rect 2822 3459 2823 3460
rect 2878 3459 2879 3460
rect 3219 3459 3220 3460
rect 2884 3461 2885 3462
rect 3216 3461 3217 3462
rect 2899 3463 2900 3464
rect 3084 3463 3085 3464
rect 2908 3465 2909 3466
rect 3102 3465 3103 3466
rect 2913 3467 2914 3468
rect 3069 3467 3070 3468
rect 2916 3469 2917 3470
rect 3063 3469 3064 3470
rect 2915 3471 2916 3472
rect 3075 3471 3076 3472
rect 2918 3473 2919 3474
rect 3282 3473 3283 3474
rect 2920 3475 2921 3476
rect 3291 3475 3292 3476
rect 2935 3477 2936 3478
rect 3264 3477 3265 3478
rect 2939 3479 2940 3480
rect 3204 3479 3205 3480
rect 2942 3481 2943 3482
rect 3129 3481 3130 3482
rect 2949 3483 2950 3484
rect 2954 3483 2955 3484
rect 2958 3483 2959 3484
rect 2972 3483 2973 3484
rect 2961 3485 2962 3486
rect 3267 3485 3268 3486
rect 2965 3487 2966 3488
rect 3330 3487 3331 3488
rect 2968 3489 2969 3490
rect 3336 3489 3337 3490
rect 2978 3491 2979 3492
rect 3315 3491 3316 3492
rect 2980 3493 2981 3494
rect 3324 3493 3325 3494
rect 2987 3495 2988 3496
rect 3162 3495 3163 3496
rect 2990 3497 2991 3498
rect 3357 3497 3358 3498
rect 2993 3499 2994 3500
rect 3315 3499 3316 3500
rect 3008 3501 3009 3502
rect 3014 3501 3015 3502
rect 3014 3503 3015 3504
rect 3027 3503 3028 3504
rect 3033 3503 3034 3504
rect 3075 3503 3076 3504
rect 3039 3505 3040 3506
rect 3093 3505 3094 3506
rect 3042 3507 3043 3508
rect 3168 3507 3169 3508
rect 3048 3509 3049 3510
rect 3096 3509 3097 3510
rect 3051 3511 3052 3512
rect 3060 3511 3061 3512
rect 3051 3513 3052 3514
rect 3105 3513 3106 3514
rect 3054 3515 3055 3516
rect 3252 3515 3253 3516
rect 3057 3517 3058 3518
rect 3138 3517 3139 3518
rect 3066 3519 3067 3520
rect 3114 3519 3115 3520
rect 3072 3521 3073 3522
rect 3120 3521 3121 3522
rect 3081 3523 3082 3524
rect 3141 3523 3142 3524
rect 3087 3525 3088 3526
rect 3207 3525 3208 3526
rect 3114 3527 3115 3528
rect 3156 3527 3157 3528
rect 3120 3529 3121 3530
rect 3180 3529 3181 3530
rect 3036 3531 3037 3532
rect 3180 3531 3181 3532
rect 3126 3533 3127 3534
rect 3165 3533 3166 3534
rect 3126 3535 3127 3536
rect 3186 3535 3187 3536
rect 3132 3537 3133 3538
rect 3192 3537 3193 3538
rect 2960 3539 2961 3540
rect 3192 3539 3193 3540
rect 3144 3541 3145 3542
rect 3234 3541 3235 3542
rect 2947 3543 2948 3544
rect 3234 3543 3235 3544
rect 3147 3545 3148 3546
rect 3237 3545 3238 3546
rect 3156 3547 3157 3548
rect 3210 3547 3211 3548
rect 3159 3549 3160 3550
rect 3213 3549 3214 3550
rect 3168 3551 3169 3552
rect 3246 3551 3247 3552
rect 2891 3553 2892 3554
rect 3246 3553 3247 3554
rect 3186 3555 3187 3556
rect 3240 3555 3241 3556
rect 3189 3557 3190 3558
rect 3243 3557 3244 3558
rect 3198 3559 3199 3560
rect 3426 3559 3427 3560
rect 3198 3561 3199 3562
rect 3420 3561 3421 3562
rect 3020 3563 3021 3564
rect 3420 3563 3421 3564
rect 3201 3565 3202 3566
rect 3450 3565 3451 3566
rect 3204 3567 3205 3568
rect 3258 3567 3259 3568
rect 3222 3569 3223 3570
rect 3270 3569 3271 3570
rect 3225 3571 3226 3572
rect 3273 3571 3274 3572
rect 3240 3573 3241 3574
rect 3294 3573 3295 3574
rect 3249 3575 3250 3576
rect 3288 3575 3289 3576
rect 3252 3577 3253 3578
rect 3300 3577 3301 3578
rect 3255 3579 3256 3580
rect 3432 3579 3433 3580
rect 3258 3581 3259 3582
rect 3342 3581 3343 3582
rect 3264 3583 3265 3584
rect 3312 3583 3313 3584
rect 3270 3585 3271 3586
rect 3408 3585 3409 3586
rect 3276 3587 3277 3588
rect 3766 3587 3767 3588
rect 3276 3589 3277 3590
rect 3318 3589 3319 3590
rect 3023 3591 3024 3592
rect 3318 3591 3319 3592
rect 3279 3593 3280 3594
rect 3339 3593 3340 3594
rect 3282 3595 3283 3596
rect 3366 3595 3367 3596
rect 3174 3597 3175 3598
rect 3366 3597 3367 3598
rect 3174 3599 3175 3600
rect 3228 3599 3229 3600
rect 3228 3601 3229 3602
rect 3306 3601 3307 3602
rect 3288 3603 3289 3604
rect 3378 3603 3379 3604
rect 3291 3605 3292 3606
rect 3381 3605 3382 3606
rect 3294 3607 3295 3608
rect 3360 3607 3361 3608
rect 3300 3609 3301 3610
rect 3414 3609 3415 3610
rect 3306 3611 3307 3612
rect 3348 3611 3349 3612
rect 3312 3613 3313 3614
rect 3354 3613 3355 3614
rect 3321 3615 3322 3616
rect 3423 3615 3424 3616
rect 3324 3617 3325 3618
rect 3363 3617 3364 3618
rect 3330 3619 3331 3620
rect 3372 3619 3373 3620
rect 3348 3621 3349 3622
rect 3390 3621 3391 3622
rect 3354 3623 3355 3624
rect 3396 3623 3397 3624
rect 3369 3625 3370 3626
rect 3375 3625 3376 3626
rect 3378 3625 3379 3626
rect 3453 3625 3454 3626
rect 3384 3627 3385 3628
rect 3453 3627 3454 3628
rect 3150 3629 3151 3630
rect 3384 3629 3385 3630
rect 2956 3631 2957 3632
rect 3150 3631 3151 3632
rect 3390 3631 3391 3632
rect 3723 3631 3724 3632
rect 3396 3633 3397 3634
rect 3459 3633 3460 3634
rect 3402 3635 3403 3636
rect 3720 3635 3721 3636
rect 3408 3637 3409 3638
rect 3777 3637 3778 3638
rect 3414 3639 3415 3640
rect 3504 3639 3505 3640
rect 3417 3641 3418 3642
rect 3501 3641 3502 3642
rect 3426 3643 3427 3644
rect 3489 3643 3490 3644
rect 3429 3645 3430 3646
rect 3748 3645 3749 3646
rect 3432 3647 3433 3648
rect 3477 3647 3478 3648
rect 3435 3649 3436 3650
rect 3894 3649 3895 3650
rect 3444 3651 3445 3652
rect 3507 3651 3508 3652
rect 3456 3653 3457 3654
rect 3552 3653 3553 3654
rect 3465 3655 3466 3656
rect 3787 3655 3788 3656
rect 3468 3657 3469 3658
rect 3540 3657 3541 3658
rect 3471 3659 3472 3660
rect 3780 3659 3781 3660
rect 3474 3661 3475 3662
rect 3525 3661 3526 3662
rect 3483 3663 3484 3664
rect 3723 3663 3724 3664
rect 3489 3665 3490 3666
rect 3558 3665 3559 3666
rect 3045 3667 3046 3668
rect 3558 3667 3559 3668
rect 3495 3669 3496 3670
rect 3531 3669 3532 3670
rect 3501 3671 3502 3672
rect 3576 3671 3577 3672
rect 3507 3673 3508 3674
rect 3570 3673 3571 3674
rect 3510 3675 3511 3676
rect 3573 3675 3574 3676
rect 3513 3677 3514 3678
rect 3567 3677 3568 3678
rect 3513 3679 3514 3680
rect 3594 3679 3595 3680
rect 3441 3681 3442 3682
rect 3594 3681 3595 3682
rect 3519 3683 3520 3684
rect 3582 3683 3583 3684
rect 3525 3685 3526 3686
rect 3763 3685 3764 3686
rect 3534 3687 3535 3688
rect 3591 3687 3592 3688
rect 3537 3689 3538 3690
rect 3857 3689 3858 3690
rect 3543 3691 3544 3692
rect 3897 3691 3898 3692
rect 3549 3693 3550 3694
rect 3821 3693 3822 3694
rect 3561 3695 3562 3696
rect 3624 3695 3625 3696
rect 3573 3697 3574 3698
rect 3612 3697 3613 3698
rect 3579 3699 3580 3700
rect 3756 3699 3757 3700
rect 3585 3701 3586 3702
rect 3759 3701 3760 3702
rect 3597 3703 3598 3704
rect 3753 3703 3754 3704
rect 3600 3705 3601 3706
rect 3835 3705 3836 3706
rect 3615 3707 3616 3708
rect 3660 3707 3661 3708
rect 3621 3709 3622 3710
rect 3699 3709 3700 3710
rect 3387 3711 3388 3712
rect 3699 3711 3700 3712
rect 3624 3713 3625 3714
rect 3702 3713 3703 3714
rect 3627 3715 3628 3716
rect 3669 3715 3670 3716
rect 3630 3717 3631 3718
rect 3744 3717 3745 3718
rect 3645 3719 3646 3720
rect 3755 3719 3756 3720
rect 3645 3721 3646 3722
rect 3705 3721 3706 3722
rect 3651 3723 3652 3724
rect 3752 3723 3753 3724
rect 3666 3725 3667 3726
rect 3857 3725 3858 3726
rect 3648 3727 3649 3728
rect 3666 3727 3667 3728
rect 3642 3729 3643 3730
rect 3648 3729 3649 3730
rect 3672 3729 3673 3730
rect 3687 3729 3688 3730
rect 3675 3731 3676 3732
rect 3690 3731 3691 3732
rect 3684 3733 3685 3734
rect 3693 3733 3694 3734
rect 3687 3735 3688 3736
rect 3696 3735 3697 3736
rect 3633 3737 3634 3738
rect 3696 3737 3697 3738
rect 3633 3739 3634 3740
rect 3681 3739 3682 3740
rect 3702 3739 3703 3740
rect 3714 3739 3715 3740
rect 3705 3741 3706 3742
rect 3717 3741 3718 3742
rect 3720 3741 3721 3742
rect 3738 3741 3739 3742
rect 3654 3743 3655 3744
rect 3738 3743 3739 3744
rect 3726 3745 3727 3746
rect 3732 3745 3733 3746
rect 3741 3745 3742 3746
rect 3842 3745 3843 3746
rect 3660 3747 3661 3748
rect 3741 3747 3742 3748
rect 3750 3747 3751 3748
rect 3873 3747 3874 3748
rect 3770 3749 3771 3750
rect 3851 3749 3852 3750
rect 3778 3751 3779 3752
rect 3831 3751 3832 3752
rect 3784 3753 3785 3754
rect 3790 3753 3791 3754
rect 3787 3755 3788 3756
rect 3793 3755 3794 3756
rect 3790 3757 3791 3758
rect 3796 3757 3797 3758
rect 3796 3759 3797 3760
rect 3863 3759 3864 3760
rect 3799 3761 3800 3762
rect 3868 3761 3869 3762
rect 3808 3763 3809 3764
rect 3814 3763 3815 3764
rect 3735 3765 3736 3766
rect 3814 3765 3815 3766
rect 3811 3767 3812 3768
rect 3817 3767 3818 3768
rect 3729 3769 3730 3770
rect 3817 3769 3818 3770
rect 3838 3769 3839 3770
rect 3848 3769 3849 3770
rect 3848 3771 3849 3772
rect 3854 3771 3855 3772
rect 3860 3771 3861 3772
rect 3887 3771 3888 3772
rect 3564 3773 3565 3774
rect 3861 3773 3862 3774
rect 2881 3782 2882 3783
rect 3219 3782 3220 3783
rect 2893 3784 2894 3785
rect 3246 3784 3247 3785
rect 2904 3786 2905 3787
rect 3361 3786 3362 3787
rect 2908 3788 2909 3789
rect 3430 3788 3431 3789
rect 2915 3790 2916 3791
rect 2926 3790 2927 3791
rect 2942 3790 2943 3791
rect 3238 3790 3239 3791
rect 2946 3792 2947 3793
rect 2957 3792 2958 3793
rect 2949 3794 2950 3795
rect 3346 3794 3347 3795
rect 2960 3796 2961 3797
rect 3198 3796 3199 3797
rect 2963 3798 2964 3799
rect 3008 3798 3009 3799
rect 2918 3800 2919 3801
rect 3008 3800 3009 3801
rect 2953 3802 2954 3803
rect 2964 3802 2965 3803
rect 2953 3804 2954 3805
rect 3189 3804 3190 3805
rect 2967 3806 2968 3807
rect 3412 3806 3413 3807
rect 2972 3808 2973 3809
rect 2990 3808 2991 3809
rect 2971 3810 2972 3811
rect 3279 3810 3280 3811
rect 2884 3812 2885 3813
rect 3280 3812 3281 3813
rect 2978 3814 2979 3815
rect 2996 3814 2997 3815
rect 2978 3816 2979 3817
rect 3163 3816 3164 3817
rect 2981 3818 2982 3819
rect 3132 3818 3133 3819
rect 3014 3820 3015 3821
rect 3382 3820 3383 3821
rect 3017 3822 3018 3823
rect 3436 3822 3437 3823
rect 2950 3824 2951 3825
rect 3017 3824 3018 3825
rect 3036 3824 3037 3825
rect 3321 3824 3322 3825
rect 3039 3826 3040 3827
rect 3130 3826 3131 3827
rect 3038 3828 3039 3829
rect 3315 3828 3316 3829
rect 3042 3830 3043 3831
rect 3472 3830 3473 3831
rect 3045 3832 3046 3833
rect 3324 3832 3325 3833
rect 3048 3834 3049 3835
rect 3058 3834 3059 3835
rect 3048 3836 3049 3837
rect 3310 3836 3311 3837
rect 3060 3838 3061 3839
rect 3064 3838 3065 3839
rect 3066 3838 3067 3839
rect 3070 3838 3071 3839
rect 3081 3838 3082 3839
rect 3106 3838 3107 3839
rect 3084 3840 3085 3841
rect 3364 3840 3365 3841
rect 3112 3842 3113 3843
rect 3138 3842 3139 3843
rect 3114 3844 3115 3845
rect 3118 3844 3119 3845
rect 3120 3844 3121 3845
rect 3190 3844 3191 3845
rect 3124 3846 3125 3847
rect 3648 3846 3649 3847
rect 3126 3848 3127 3849
rect 3487 3848 3488 3849
rect 3139 3850 3140 3851
rect 3366 3850 3367 3851
rect 3144 3852 3145 3853
rect 3232 3852 3233 3853
rect 3156 3854 3157 3855
rect 3274 3854 3275 3855
rect 2922 3856 2923 3857
rect 3157 3856 3158 3857
rect 3168 3856 3169 3857
rect 3244 3856 3245 3857
rect 3174 3858 3175 3859
rect 3298 3858 3299 3859
rect 3072 3860 3073 3861
rect 3175 3860 3176 3861
rect 3180 3860 3181 3861
rect 3184 3860 3185 3861
rect 3186 3860 3187 3861
rect 3328 3860 3329 3861
rect 3204 3862 3205 3863
rect 3334 3862 3335 3863
rect 3208 3864 3209 3865
rect 3567 3864 3568 3865
rect 3222 3866 3223 3867
rect 3316 3866 3317 3867
rect 3223 3868 3224 3869
rect 3624 3868 3625 3869
rect 3225 3870 3226 3871
rect 3337 3870 3338 3871
rect 3150 3872 3151 3873
rect 3226 3872 3227 3873
rect 3228 3872 3229 3873
rect 3262 3872 3263 3873
rect 3234 3874 3235 3875
rect 3304 3874 3305 3875
rect 3240 3876 3241 3877
rect 3367 3876 3368 3877
rect 3087 3878 3088 3879
rect 3241 3878 3242 3879
rect 3075 3880 3076 3881
rect 3088 3880 3089 3881
rect 3054 3882 3055 3883
rect 3076 3882 3077 3883
rect 3055 3884 3056 3885
rect 3439 3884 3440 3885
rect 3256 3886 3257 3887
rect 3480 3886 3481 3887
rect 3258 3888 3259 3889
rect 3340 3888 3341 3889
rect 3264 3890 3265 3891
rect 3394 3890 3395 3891
rect 3276 3892 3277 3893
rect 3406 3892 3407 3893
rect 3282 3894 3283 3895
rect 3373 3894 3374 3895
rect 3159 3896 3160 3897
rect 3283 3896 3284 3897
rect 3286 3896 3287 3897
rect 3300 3896 3301 3897
rect 3288 3898 3289 3899
rect 3755 3898 3756 3899
rect 3291 3900 3292 3901
rect 3376 3900 3377 3901
rect 3252 3902 3253 3903
rect 3292 3902 3293 3903
rect 3294 3902 3295 3903
rect 3442 3902 3443 3903
rect 3306 3904 3307 3905
rect 3478 3904 3479 3905
rect 3312 3906 3313 3907
rect 3484 3906 3485 3907
rect 3318 3908 3319 3909
rect 3322 3908 3323 3909
rect 3369 3908 3370 3909
rect 3505 3908 3506 3909
rect 3378 3910 3379 3911
rect 3448 3910 3449 3911
rect 3249 3912 3250 3913
rect 3379 3912 3380 3913
rect 3250 3914 3251 3915
rect 3531 3914 3532 3915
rect 3384 3916 3385 3917
rect 3403 3916 3404 3917
rect 3387 3918 3388 3919
rect 3400 3918 3401 3919
rect 3390 3920 3391 3921
rect 3553 3920 3554 3921
rect 3396 3922 3397 3923
rect 3547 3922 3548 3923
rect 3408 3924 3409 3925
rect 3762 3924 3763 3925
rect 2939 3926 2940 3927
rect 3409 3926 3410 3927
rect 2929 3928 2930 3929
rect 2938 3928 2939 3929
rect 3417 3928 3418 3929
rect 3424 3928 3425 3929
rect 3418 3930 3419 3931
rect 3585 3930 3586 3931
rect 3420 3932 3421 3933
rect 3466 3932 3467 3933
rect 3444 3934 3445 3935
rect 3571 3934 3572 3935
rect 3033 3936 3034 3937
rect 3445 3936 3446 3937
rect 3032 3938 3033 3939
rect 3147 3938 3148 3939
rect 3450 3938 3451 3939
rect 3523 3938 3524 3939
rect 3456 3940 3457 3941
rect 3589 3940 3590 3941
rect 3468 3942 3469 3943
rect 3613 3942 3614 3943
rect 3469 3944 3470 3945
rect 3621 3944 3622 3945
rect 3474 3946 3475 3947
rect 3943 3946 3944 3947
rect 3489 3948 3490 3949
rect 3637 3948 3638 3949
rect 3453 3950 3454 3951
rect 3490 3950 3491 3951
rect 3454 3952 3455 3953
rect 3708 3952 3709 3953
rect 3496 3954 3497 3955
rect 3654 3954 3655 3955
rect 3501 3956 3502 3957
rect 3619 3956 3620 3957
rect 3330 3958 3331 3959
rect 3502 3958 3503 3959
rect 2897 3960 2898 3961
rect 3331 3960 3332 3961
rect 2896 3962 2897 3963
rect 3216 3962 3217 3963
rect 3507 3962 3508 3963
rect 3649 3962 3650 3963
rect 3354 3964 3355 3965
rect 3508 3964 3509 3965
rect 3510 3964 3511 3965
rect 3896 3964 3897 3965
rect 3414 3966 3415 3967
rect 3511 3966 3512 3967
rect 3267 3968 3268 3969
rect 3415 3968 3416 3969
rect 3192 3970 3193 3971
rect 3268 3970 3269 3971
rect 3513 3970 3514 3971
rect 3655 3970 3656 3971
rect 3525 3972 3526 3973
rect 3882 3972 3883 3973
rect 3526 3974 3527 3975
rect 3731 3974 3732 3975
rect 3529 3976 3530 3977
rect 3594 3976 3595 3977
rect 3532 3978 3533 3979
rect 3660 3978 3661 3979
rect 3519 3980 3520 3981
rect 3661 3980 3662 3981
rect 3348 3982 3349 3983
rect 3520 3982 3521 3983
rect 3270 3984 3271 3985
rect 3349 3984 3350 3985
rect 3537 3984 3538 3985
rect 3915 3984 3916 3985
rect 3538 3986 3539 3987
rect 3734 3986 3735 3987
rect 3541 3988 3542 3989
rect 3558 3988 3559 3989
rect 3543 3990 3544 3991
rect 3918 3990 3919 3991
rect 3549 3992 3550 3993
rect 3770 3992 3771 3993
rect 3555 3994 3556 3995
rect 3591 3994 3592 3995
rect 3559 3996 3560 3997
rect 3842 3996 3843 3997
rect 3561 3998 3562 3999
rect 3631 3998 3632 3999
rect 3573 4000 3574 4001
rect 3577 4000 3578 4001
rect 3579 4000 3580 4001
rect 3711 4000 3712 4001
rect 3580 4002 3581 4003
rect 3752 4002 3753 4003
rect 3597 4004 3598 4005
rect 3764 4004 3765 4005
rect 3600 4006 3601 4007
rect 3625 4006 3626 4007
rect 3432 4008 3433 4009
rect 3601 4008 3602 4009
rect 3051 4010 3052 4011
rect 3433 4010 3434 4011
rect 3607 4010 3608 4011
rect 3675 4010 3676 4011
rect 3627 4012 3628 4013
rect 3868 4012 3869 4013
rect 3633 4014 3634 4015
rect 3743 4014 3744 4015
rect 3643 4016 3644 4017
rect 3861 4016 3862 4017
rect 3645 4018 3646 4019
rect 3773 4018 3774 4019
rect 3651 4020 3652 4021
rect 3821 4020 3822 4021
rect 3426 4022 3427 4023
rect 3652 4022 3653 4023
rect 3666 4022 3667 4023
rect 3741 4022 3742 4023
rect 3667 4024 3668 4025
rect 3946 4024 3947 4025
rect 3670 4026 3671 4027
rect 3885 4026 3886 4027
rect 3684 4028 3685 4029
rect 3691 4028 3692 4029
rect 3694 4030 3695 4031
rect 3857 4030 3858 4031
rect 3705 4032 3706 4033
rect 3752 4032 3753 4033
rect 3615 4034 3616 4035
rect 3706 4034 3707 4035
rect 3720 4034 3721 4035
rect 3776 4034 3777 4035
rect 3721 4036 3722 4037
rect 3766 4036 3767 4037
rect 3726 4038 3727 4039
rect 3817 4038 3818 4039
rect 3696 4040 3697 4041
rect 3727 4040 3728 4041
rect 3729 4040 3730 4041
rect 3767 4040 3768 4041
rect 3737 4042 3738 4043
rect 3787 4042 3788 4043
rect 3748 4044 3749 4045
rect 3759 4044 3760 4045
rect 3460 4046 3461 4047
rect 3758 4046 3759 4047
rect 3702 4048 3703 4049
rect 3749 4048 3750 4049
rect 3761 4048 3762 4049
rect 3889 4048 3890 4049
rect 3778 4050 3779 4051
rect 3814 4050 3815 4051
rect 3723 4052 3724 4053
rect 3779 4052 3780 4053
rect 3784 4052 3785 4053
rect 3862 4052 3863 4053
rect 3790 4054 3791 4055
rect 3838 4054 3839 4055
rect 3796 4056 3797 4057
rect 3844 4056 3845 4057
rect 3808 4058 3809 4059
rect 3856 4058 3857 4059
rect 3718 4060 3719 4061
rect 3808 4060 3809 4061
rect 3811 4060 3812 4061
rect 3859 4060 3860 4061
rect 3672 4062 3673 4063
rect 3811 4062 3812 4063
rect 3820 4062 3821 4063
rect 3831 4062 3832 4063
rect 3848 4062 3849 4063
rect 3902 4062 3903 4063
rect 3799 4064 3800 4065
rect 3847 4064 3848 4065
rect 3851 4064 3852 4065
rect 3905 4064 3906 4065
rect 3865 4066 3866 4067
rect 3878 4066 3879 4067
rect 3925 4066 3926 4067
rect 3929 4066 3930 4067
rect 2809 4075 2810 4076
rect 3175 4075 3176 4076
rect 2887 4077 2888 4078
rect 3280 4077 3281 4078
rect 2907 4079 2908 4080
rect 3058 4079 3059 4080
rect 2918 4081 2919 4082
rect 3433 4081 3434 4082
rect 2922 4083 2923 4084
rect 3430 4083 3431 4084
rect 2926 4085 2927 4086
rect 3457 4085 3458 4086
rect 2925 4087 2926 4088
rect 3394 4087 3395 4088
rect 2928 4089 2929 4090
rect 3391 4089 3392 4090
rect 2935 4091 2936 4092
rect 3316 4091 3317 4092
rect 2941 4093 2942 4094
rect 3298 4093 3299 4094
rect 2944 4095 2945 4096
rect 3385 4095 3386 4096
rect 2947 4097 2948 4098
rect 3286 4097 3287 4098
rect 2954 4099 2955 4100
rect 3346 4099 3347 4100
rect 2961 4101 2962 4102
rect 3190 4101 3191 4102
rect 2971 4103 2972 4104
rect 3430 4103 3431 4104
rect 2981 4105 2982 4106
rect 3487 4105 3488 4106
rect 2984 4107 2985 4108
rect 2990 4107 2991 4108
rect 2996 4107 2997 4108
rect 3739 4107 3740 4108
rect 2996 4109 2997 4110
rect 3172 4109 3173 4110
rect 3026 4111 3027 4112
rect 3032 4111 3033 4112
rect 3038 4111 3039 4112
rect 3472 4111 3473 4112
rect 3041 4113 3042 4114
rect 3436 4113 3437 4114
rect 3042 4115 3043 4116
rect 3382 4115 3383 4116
rect 3045 4117 3046 4118
rect 3064 4117 3065 4118
rect 2899 4119 2900 4120
rect 3045 4119 3046 4120
rect 3048 4119 3049 4120
rect 3292 4119 3293 4120
rect 2896 4121 2897 4122
rect 3292 4121 3293 4122
rect 3052 4123 3053 4124
rect 3403 4123 3404 4124
rect 2903 4125 2904 4126
rect 3051 4125 3052 4126
rect 3057 4125 3058 4126
rect 3310 4125 3311 4126
rect 3076 4127 3077 4128
rect 3081 4127 3082 4128
rect 3070 4129 3071 4130
rect 3075 4129 3076 4130
rect 3088 4129 3089 4130
rect 3093 4129 3094 4130
rect 3112 4129 3113 4130
rect 3132 4129 3133 4130
rect 3111 4131 3112 4132
rect 3147 4131 3148 4132
rect 3124 4133 3125 4134
rect 3517 4133 3518 4134
rect 3151 4135 3152 4136
rect 3487 4135 3488 4136
rect 3154 4137 3155 4138
rect 3286 4137 3287 4138
rect 3160 4139 3161 4140
rect 3163 4139 3164 4140
rect 3178 4139 3179 4140
rect 3184 4139 3185 4140
rect 2958 4141 2959 4142
rect 3184 4141 3185 4142
rect 3190 4141 3191 4142
rect 3523 4141 3524 4142
rect 3196 4143 3197 4144
rect 3211 4143 3212 4144
rect 3202 4145 3203 4146
rect 3409 4145 3410 4146
rect 3214 4147 3215 4148
rect 3232 4147 3233 4148
rect 3220 4149 3221 4150
rect 3226 4149 3227 4150
rect 3014 4151 3015 4152
rect 3226 4151 3227 4152
rect 3229 4151 3230 4152
rect 3439 4151 3440 4152
rect 3232 4153 3233 4154
rect 3238 4153 3239 4154
rect 3238 4155 3239 4156
rect 3244 4155 3245 4156
rect 3208 4157 3209 4158
rect 3244 4157 3245 4158
rect 3208 4159 3209 4160
rect 3424 4159 3425 4160
rect 3250 4161 3251 4162
rect 3727 4161 3728 4162
rect 3256 4163 3257 4164
rect 3316 4163 3317 4164
rect 3256 4165 3257 4166
rect 3262 4165 3263 4166
rect 3262 4167 3263 4168
rect 3274 4167 3275 4168
rect 3265 4169 3266 4170
rect 3283 4169 3284 4170
rect 3268 4171 3269 4172
rect 3274 4171 3275 4172
rect 2950 4173 2951 4174
rect 3268 4173 3269 4174
rect 3280 4173 3281 4174
rect 3322 4173 3323 4174
rect 3298 4175 3299 4176
rect 3304 4175 3305 4176
rect 2910 4177 2911 4178
rect 3304 4177 3305 4178
rect 3310 4177 3311 4178
rect 3334 4177 3335 4178
rect 3223 4179 3224 4180
rect 3334 4179 3335 4180
rect 3322 4181 3323 4182
rect 3328 4181 3329 4182
rect 2951 4183 2952 4184
rect 3328 4183 3329 4184
rect 3325 4185 3326 4186
rect 3331 4185 3332 4186
rect 3337 4185 3338 4186
rect 3352 4185 3353 4186
rect 2906 4187 2907 4188
rect 3337 4187 3338 4188
rect 3340 4187 3341 4188
rect 3343 4187 3344 4188
rect 3355 4187 3356 4188
rect 3367 4187 3368 4188
rect 3349 4189 3350 4190
rect 3367 4189 3368 4190
rect 2938 4191 2939 4192
rect 3349 4191 3350 4192
rect 3373 4191 3374 4192
rect 3397 4191 3398 4192
rect 3379 4193 3380 4194
rect 3394 4193 3395 4194
rect 3403 4193 3404 4194
rect 3496 4193 3497 4194
rect 3406 4195 3407 4196
rect 3427 4195 3428 4196
rect 3412 4197 3413 4198
rect 3421 4197 3422 4198
rect 3415 4199 3416 4200
rect 3424 4199 3425 4200
rect 3169 4201 3170 4202
rect 3415 4201 3416 4202
rect 3433 4201 3434 4202
rect 3466 4201 3467 4202
rect 3439 4203 3440 4204
rect 3442 4203 3443 4204
rect 3442 4205 3443 4206
rect 3445 4205 3446 4206
rect 3448 4205 3449 4206
rect 3734 4205 3735 4206
rect 3451 4207 3452 4208
rect 3460 4207 3461 4208
rect 3241 4209 3242 4210
rect 3460 4209 3461 4210
rect 3454 4211 3455 4212
rect 3463 4211 3464 4212
rect 3466 4211 3467 4212
rect 3469 4211 3470 4212
rect 3475 4211 3476 4212
rect 3526 4211 3527 4212
rect 3478 4213 3479 4214
rect 3493 4213 3494 4214
rect 3481 4215 3482 4216
rect 3490 4215 3491 4216
rect 3484 4217 3485 4218
rect 3499 4217 3500 4218
rect 3505 4217 3506 4218
rect 3526 4217 3527 4218
rect 3505 4219 3506 4220
rect 3529 4219 3530 4220
rect 3508 4221 3509 4222
rect 3529 4221 3530 4222
rect 3508 4223 3509 4224
rect 3797 4223 3798 4224
rect 3520 4225 3521 4226
rect 3535 4225 3536 4226
rect 3400 4227 3401 4228
rect 3520 4227 3521 4228
rect 3376 4229 3377 4230
rect 3400 4229 3401 4230
rect 3532 4229 3533 4230
rect 3709 4229 3710 4230
rect 3511 4231 3512 4232
rect 3532 4231 3533 4232
rect 3502 4233 3503 4234
rect 3511 4233 3512 4234
rect 2975 4235 2976 4236
rect 3502 4235 3503 4236
rect 3538 4235 3539 4236
rect 3782 4235 3783 4236
rect 3032 4237 3033 4238
rect 3538 4237 3539 4238
rect 3541 4237 3542 4238
rect 3562 4237 3563 4238
rect 3547 4239 3548 4240
rect 3568 4239 3569 4240
rect 3547 4241 3548 4242
rect 3801 4241 3802 4242
rect 3418 4243 3419 4244
rect 3800 4243 3801 4244
rect 3553 4245 3554 4246
rect 3574 4245 3575 4246
rect 3553 4247 3554 4248
rect 3577 4247 3578 4248
rect 3571 4249 3572 4250
rect 3586 4249 3587 4250
rect 3577 4251 3578 4252
rect 3580 4251 3581 4252
rect 3559 4253 3560 4254
rect 3580 4253 3581 4254
rect 3559 4255 3560 4256
rect 3816 4255 3817 4256
rect 3589 4257 3590 4258
rect 3598 4257 3599 4258
rect 3601 4257 3602 4258
rect 3616 4257 3617 4258
rect 3604 4259 3605 4260
rect 3652 4259 3653 4260
rect 3607 4261 3608 4262
rect 3610 4261 3611 4262
rect 3613 4261 3614 4262
rect 3628 4261 3629 4262
rect 3619 4263 3620 4264
rect 3622 4263 3623 4264
rect 3625 4263 3626 4264
rect 3634 4263 3635 4264
rect 3631 4265 3632 4266
rect 3755 4265 3756 4266
rect 3637 4267 3638 4268
rect 3652 4267 3653 4268
rect 3643 4269 3644 4270
rect 3658 4269 3659 4270
rect 3646 4271 3647 4272
rect 3649 4271 3650 4272
rect 3655 4271 3656 4272
rect 3664 4271 3665 4272
rect 3667 4271 3668 4272
rect 3685 4271 3686 4272
rect 3682 4273 3683 4274
rect 3941 4273 3942 4274
rect 3694 4275 3695 4276
rect 3712 4275 3713 4276
rect 3694 4277 3695 4278
rect 3871 4277 3872 4278
rect 3706 4279 3707 4280
rect 3724 4279 3725 4280
rect 3691 4281 3692 4282
rect 3706 4281 3707 4282
rect 3721 4281 3722 4282
rect 3808 4281 3809 4282
rect 3721 4283 3722 4284
rect 3915 4283 3916 4284
rect 3731 4285 3732 4286
rect 3826 4285 3827 4286
rect 3743 4287 3744 4288
rect 3922 4287 3923 4288
rect 3749 4289 3750 4290
rect 3758 4289 3759 4290
rect 3749 4291 3750 4292
rect 3951 4291 3952 4292
rect 3767 4293 3768 4294
rect 3788 4293 3789 4294
rect 3773 4295 3774 4296
rect 3794 4295 3795 4296
rect 3776 4297 3777 4298
rect 3874 4297 3875 4298
rect 3761 4299 3762 4300
rect 3776 4299 3777 4300
rect 3752 4301 3753 4302
rect 3761 4301 3762 4302
rect 3779 4301 3780 4302
rect 3908 4301 3909 4302
rect 3764 4303 3765 4304
rect 3779 4303 3780 4304
rect 3782 4303 3783 4304
rect 3927 4303 3928 4304
rect 3785 4305 3786 4306
rect 3792 4305 3793 4306
rect 3770 4307 3771 4308
rect 3791 4307 3792 4308
rect 3688 4309 3689 4310
rect 3770 4309 3771 4310
rect 3661 4311 3662 4312
rect 3688 4311 3689 4312
rect 3785 4311 3786 4312
rect 3931 4311 3932 4312
rect 3814 4313 3815 4314
rect 3889 4313 3890 4314
rect 3670 4315 3671 4316
rect 3888 4315 3889 4316
rect 3670 4317 3671 4318
rect 3899 4317 3900 4318
rect 3820 4319 3821 4320
rect 3835 4319 3836 4320
rect 3523 4321 3524 4322
rect 3819 4321 3820 4322
rect 3838 4321 3839 4322
rect 3871 4321 3872 4322
rect 3844 4323 3845 4324
rect 3868 4323 3869 4324
rect 3847 4325 3848 4326
rect 3850 4325 3851 4326
rect 3847 4327 3848 4328
rect 3918 4327 3919 4328
rect 3853 4329 3854 4330
rect 3865 4329 3866 4330
rect 3856 4331 3857 4332
rect 3865 4331 3866 4332
rect 3737 4333 3738 4334
rect 3856 4333 3857 4334
rect 3859 4333 3860 4334
rect 3868 4333 3869 4334
rect 3862 4335 3863 4336
rect 3878 4335 3879 4336
rect 3882 4335 3883 4336
rect 3924 4335 3925 4336
rect 3898 4337 3899 4338
rect 3936 4337 3937 4338
rect 3905 4339 3906 4340
rect 3907 4339 3908 4340
rect 3902 4341 3903 4342
rect 3904 4341 3905 4342
rect 3901 4343 3902 4344
rect 3917 4343 3918 4344
rect 2882 4352 2883 4353
rect 2991 4352 2992 4353
rect 2890 4354 2891 4355
rect 3262 4354 3263 4355
rect 2896 4356 2897 4357
rect 3322 4356 3323 4357
rect 2899 4358 2900 4359
rect 2921 4358 2922 4359
rect 2906 4360 2907 4361
rect 3364 4360 3365 4361
rect 2909 4362 2910 4363
rect 3340 4362 3341 4363
rect 2925 4364 2926 4365
rect 2972 4364 2973 4365
rect 2924 4366 2925 4367
rect 3406 4366 3407 4367
rect 2928 4368 2929 4369
rect 3385 4368 3386 4369
rect 2932 4370 2933 4371
rect 3292 4370 3293 4371
rect 2933 4372 2934 4373
rect 3310 4372 3311 4373
rect 2947 4374 2948 4375
rect 3349 4374 3350 4375
rect 2954 4376 2955 4377
rect 3238 4376 3239 4377
rect 2957 4378 2958 4379
rect 3427 4378 3428 4379
rect 2961 4380 2962 4381
rect 3331 4380 3332 4381
rect 2961 4382 2962 4383
rect 3493 4382 3494 4383
rect 2964 4384 2965 4385
rect 3181 4384 3182 4385
rect 2973 4386 2974 4387
rect 2984 4386 2985 4387
rect 2975 4388 2976 4389
rect 3211 4388 3212 4389
rect 2979 4390 2980 4391
rect 2996 4390 2997 4391
rect 2994 4392 2995 4393
rect 3265 4392 3266 4393
rect 2876 4394 2877 4395
rect 3265 4394 3266 4395
rect 2997 4396 2998 4397
rect 3008 4396 3009 4397
rect 2872 4398 2873 4399
rect 3009 4398 3010 4399
rect 3003 4400 3004 4401
rect 3226 4400 3227 4401
rect 3017 4402 3018 4403
rect 3502 4402 3503 4403
rect 3018 4404 3019 4405
rect 3026 4404 3027 4405
rect 3024 4406 3025 4407
rect 3256 4406 3257 4407
rect 3032 4408 3033 4409
rect 3421 4408 3422 4409
rect 3035 4410 3036 4411
rect 3583 4410 3584 4411
rect 2943 4412 2944 4413
rect 3036 4412 3037 4413
rect 3045 4412 3046 4413
rect 3048 4412 3049 4413
rect 3051 4412 3052 4413
rect 3054 4412 3055 4413
rect 3057 4412 3058 4413
rect 3502 4412 3503 4413
rect 3057 4414 3058 4415
rect 3325 4414 3326 4415
rect 3075 4416 3076 4417
rect 3078 4416 3079 4417
rect 3090 4416 3091 4417
rect 3093 4416 3094 4417
rect 3096 4416 3097 4417
rect 3111 4416 3112 4417
rect 3105 4418 3106 4419
rect 3108 4418 3109 4419
rect 3117 4418 3118 4419
rect 3120 4418 3121 4419
rect 3126 4418 3127 4419
rect 3132 4418 3133 4419
rect 3132 4420 3133 4421
rect 3160 4420 3161 4421
rect 3135 4422 3136 4423
rect 3814 4422 3815 4423
rect 3138 4424 3139 4425
rect 3934 4424 3935 4425
rect 3139 4426 3140 4427
rect 3196 4426 3197 4427
rect 2892 4428 2893 4429
rect 3196 4428 3197 4429
rect 3142 4430 3143 4431
rect 3199 4430 3200 4431
rect 3144 4432 3145 4433
rect 3217 4432 3218 4433
rect 3129 4434 3130 4435
rect 3145 4434 3146 4435
rect 3151 4434 3152 4435
rect 3816 4434 3817 4435
rect 3154 4436 3155 4437
rect 3481 4436 3482 4437
rect 3166 4438 3167 4439
rect 3190 4438 3191 4439
rect 3178 4440 3179 4441
rect 3190 4440 3191 4441
rect 3157 4442 3158 4443
rect 3178 4442 3179 4443
rect 3157 4444 3158 4445
rect 3310 4444 3311 4445
rect 3184 4446 3185 4447
rect 3205 4446 3206 4447
rect 3214 4446 3215 4447
rect 3253 4446 3254 4447
rect 3220 4448 3221 4449
rect 3235 4448 3236 4449
rect 3223 4450 3224 4451
rect 3244 4450 3245 4451
rect 3229 4452 3230 4453
rect 3409 4452 3410 4453
rect 3202 4454 3203 4455
rect 3229 4454 3230 4455
rect 3232 4454 3233 4455
rect 3241 4454 3242 4455
rect 3247 4454 3248 4455
rect 3316 4454 3317 4455
rect 3262 4456 3263 4457
rect 3334 4456 3335 4457
rect 3274 4458 3275 4459
rect 3292 4458 3293 4459
rect 3274 4460 3275 4461
rect 3280 4460 3281 4461
rect 3268 4462 3269 4463
rect 3280 4462 3281 4463
rect 3147 4464 3148 4465
rect 3268 4464 3269 4465
rect 3295 4464 3296 4465
rect 3430 4464 3431 4465
rect 3304 4466 3305 4467
rect 3316 4466 3317 4467
rect 3298 4468 3299 4469
rect 3304 4468 3305 4469
rect 3322 4468 3323 4469
rect 3403 4468 3404 4469
rect 3334 4470 3335 4471
rect 3343 4470 3344 4471
rect 3337 4472 3338 4473
rect 3346 4472 3347 4473
rect 3355 4472 3356 4473
rect 3370 4472 3371 4473
rect 3358 4474 3359 4475
rect 3361 4474 3362 4475
rect 3081 4476 3082 4477
rect 3361 4476 3362 4477
rect 3081 4478 3082 4479
rect 3352 4478 3353 4479
rect 3352 4480 3353 4481
rect 3367 4480 3368 4481
rect 3364 4482 3365 4483
rect 3433 4482 3434 4483
rect 3367 4484 3368 4485
rect 3466 4484 3467 4485
rect 2947 4486 2948 4487
rect 3466 4486 3467 4487
rect 3382 4488 3383 4489
rect 3391 4488 3392 4489
rect 3385 4490 3386 4491
rect 3394 4490 3395 4491
rect 3388 4492 3389 4493
rect 3397 4492 3398 4493
rect 3391 4494 3392 4495
rect 3400 4494 3401 4495
rect 3042 4496 3043 4497
rect 3400 4496 3401 4497
rect 3412 4496 3413 4497
rect 3520 4496 3521 4497
rect 3415 4498 3416 4499
rect 3418 4498 3419 4499
rect 3424 4498 3425 4499
rect 3469 4498 3470 4499
rect 3424 4500 3425 4501
rect 3508 4500 3509 4501
rect 3430 4502 3431 4503
rect 3439 4502 3440 4503
rect 3433 4504 3434 4505
rect 3442 4504 3443 4505
rect 3442 4506 3443 4507
rect 3457 4506 3458 4507
rect 3445 4508 3446 4509
rect 3460 4508 3461 4509
rect 3451 4510 3452 4511
rect 3454 4510 3455 4511
rect 3460 4510 3461 4511
rect 3761 4510 3762 4511
rect 3463 4512 3464 4513
rect 3739 4512 3740 4513
rect 3472 4514 3473 4515
rect 3475 4514 3476 4515
rect 3478 4514 3479 4515
rect 3505 4514 3506 4515
rect 3481 4516 3482 4517
rect 3751 4516 3752 4517
rect 3484 4518 3485 4519
rect 3499 4518 3500 4519
rect 3487 4520 3488 4521
rect 3743 4520 3744 4521
rect 3487 4522 3488 4523
rect 3529 4522 3530 4523
rect 3490 4524 3491 4525
rect 3532 4524 3533 4525
rect 3493 4526 3494 4527
rect 3511 4526 3512 4527
rect 3499 4528 3500 4529
rect 3517 4528 3518 4529
rect 3505 4530 3506 4531
rect 3523 4530 3524 4531
rect 3508 4532 3509 4533
rect 3526 4532 3527 4533
rect 3511 4534 3512 4535
rect 3547 4534 3548 4535
rect 3517 4536 3518 4537
rect 3535 4536 3536 4537
rect 3520 4538 3521 4539
rect 3538 4538 3539 4539
rect 3523 4540 3524 4541
rect 3804 4540 3805 4541
rect 3529 4542 3530 4543
rect 3770 4542 3771 4543
rect 3532 4544 3533 4545
rect 3709 4544 3710 4545
rect 3535 4546 3536 4547
rect 3562 4546 3563 4547
rect 3541 4548 3542 4549
rect 3568 4548 3569 4549
rect 3547 4550 3548 4551
rect 3574 4550 3575 4551
rect 3553 4552 3554 4553
rect 3821 4552 3822 4553
rect 3553 4554 3554 4555
rect 3885 4554 3886 4555
rect 3556 4556 3557 4557
rect 3577 4556 3578 4557
rect 3559 4558 3560 4559
rect 3797 4558 3798 4559
rect 3559 4560 3560 4561
rect 3871 4560 3872 4561
rect 3565 4562 3566 4563
rect 3580 4562 3581 4563
rect 3571 4564 3572 4565
rect 3586 4564 3587 4565
rect 3589 4564 3590 4565
rect 3598 4564 3599 4565
rect 3595 4566 3596 4567
rect 3622 4566 3623 4567
rect 3601 4568 3602 4569
rect 3604 4568 3605 4569
rect 3613 4568 3614 4569
rect 3628 4568 3629 4569
rect 3616 4570 3617 4571
rect 3917 4570 3918 4571
rect 3625 4572 3626 4573
rect 3664 4572 3665 4573
rect 3631 4574 3632 4575
rect 3935 4574 3936 4575
rect 3634 4576 3635 4577
rect 3832 4576 3833 4577
rect 3643 4578 3644 4579
rect 3646 4578 3647 4579
rect 3649 4578 3650 4579
rect 3652 4578 3653 4579
rect 3655 4578 3656 4579
rect 3658 4578 3659 4579
rect 3667 4578 3668 4579
rect 3688 4578 3689 4579
rect 3673 4580 3674 4581
rect 3961 4580 3962 4581
rect 3682 4582 3683 4583
rect 3953 4582 3954 4583
rect 3682 4584 3683 4585
rect 3938 4584 3939 4585
rect 3685 4586 3686 4587
rect 3941 4586 3942 4587
rect 3685 4588 3686 4589
rect 3694 4588 3695 4589
rect 3691 4590 3692 4591
rect 3886 4590 3887 4591
rect 3697 4592 3698 4593
rect 3712 4592 3713 4593
rect 3703 4594 3704 4595
rect 3718 4594 3719 4595
rect 3706 4596 3707 4597
rect 3773 4596 3774 4597
rect 3610 4598 3611 4599
rect 3706 4598 3707 4599
rect 3709 4598 3710 4599
rect 3924 4598 3925 4599
rect 3721 4600 3722 4601
rect 3826 4600 3827 4601
rect 3715 4602 3716 4603
rect 3825 4602 3826 4603
rect 3733 4604 3734 4605
rect 3749 4604 3750 4605
rect 3754 4604 3755 4605
rect 3758 4604 3759 4605
rect 3757 4606 3758 4607
rect 3878 4606 3879 4607
rect 3760 4608 3761 4609
rect 3776 4608 3777 4609
rect 3577 4610 3578 4611
rect 3775 4610 3776 4611
rect 3766 4612 3767 4613
rect 3782 4612 3783 4613
rect 3769 4614 3770 4615
rect 3920 4614 3921 4615
rect 3779 4616 3780 4617
rect 3874 4616 3875 4617
rect 3791 4618 3792 4619
rect 3889 4618 3890 4619
rect 3790 4620 3791 4621
rect 3927 4620 3928 4621
rect 3785 4622 3786 4623
rect 3928 4622 3929 4623
rect 3784 4624 3785 4625
rect 3794 4624 3795 4625
rect 3793 4626 3794 4627
rect 3823 4626 3824 4627
rect 3805 4628 3806 4629
rect 3974 4628 3975 4629
rect 3808 4630 3809 4631
rect 3942 4630 3943 4631
rect 3811 4632 3812 4633
rect 3828 4632 3829 4633
rect 3835 4632 3836 4633
rect 3844 4632 3845 4633
rect 3856 4632 3857 4633
rect 3859 4632 3860 4633
rect 3853 4634 3854 4635
rect 3856 4634 3857 4635
rect 3670 4636 3671 4637
rect 3853 4636 3854 4637
rect 3865 4636 3866 4637
rect 3880 4636 3881 4637
rect 3868 4638 3869 4639
rect 3883 4638 3884 4639
rect 3874 4640 3875 4641
rect 3948 4640 3949 4641
rect 3661 4642 3662 4643
rect 3949 4642 3950 4643
rect 3877 4644 3878 4645
rect 3945 4644 3946 4645
rect 3898 4646 3899 4647
rect 3913 4646 3914 4647
rect 3901 4648 3902 4649
rect 3916 4648 3917 4649
rect 3850 4650 3851 4651
rect 3900 4650 3901 4651
rect 3847 4652 3848 4653
rect 3850 4652 3851 4653
rect 3904 4652 3905 4653
rect 3919 4652 3920 4653
rect 3724 4654 3725 4655
rect 3903 4654 3904 4655
rect 3907 4654 3908 4655
rect 3922 4654 3923 4655
rect 3763 4656 3764 4657
rect 3907 4656 3908 4657
rect 3951 4656 3952 4657
rect 3977 4656 3978 4657
rect 2876 4665 2877 4666
rect 3009 4665 3010 4666
rect 2869 4667 2870 4668
rect 2876 4667 2877 4668
rect 2872 4669 2873 4670
rect 3009 4669 3010 4670
rect 2885 4671 2886 4672
rect 2994 4671 2995 4672
rect 2892 4673 2893 4674
rect 3346 4673 3347 4674
rect 2896 4675 2897 4676
rect 3196 4675 3197 4676
rect 2899 4677 2900 4678
rect 3316 4677 3317 4678
rect 2903 4679 2904 4680
rect 2918 4679 2919 4680
rect 2906 4681 2907 4682
rect 3278 4681 3279 4682
rect 2912 4683 2913 4684
rect 3260 4683 3261 4684
rect 2926 4685 2927 4686
rect 3048 4685 3049 4686
rect 2936 4687 2937 4688
rect 3235 4687 3236 4688
rect 2936 4689 2937 4690
rect 3081 4689 3082 4690
rect 2940 4691 2941 4692
rect 2950 4691 2951 4692
rect 2943 4693 2944 4694
rect 3331 4693 3332 4694
rect 2947 4695 2948 4696
rect 3166 4695 3167 4696
rect 2959 4697 2960 4698
rect 3385 4697 3386 4698
rect 2961 4699 2962 4700
rect 3541 4699 3542 4700
rect 2964 4701 2965 4702
rect 3643 4701 3644 4702
rect 2973 4703 2974 4704
rect 3045 4703 3046 4704
rect 2991 4705 2992 4706
rect 3012 4705 3013 4706
rect 2979 4707 2980 4708
rect 2991 4707 2992 4708
rect 3003 4707 3004 4708
rect 3221 4707 3222 4708
rect 3018 4709 3019 4710
rect 3021 4709 3022 4710
rect 3024 4709 3025 4710
rect 3299 4709 3300 4710
rect 3044 4711 3045 4712
rect 3164 4711 3165 4712
rect 3047 4713 3048 4714
rect 3054 4713 3055 4714
rect 3057 4713 3058 4714
rect 3149 4713 3150 4714
rect 3065 4715 3066 4716
rect 3361 4715 3362 4716
rect 3071 4717 3072 4718
rect 3508 4717 3509 4718
rect 3078 4719 3079 4720
rect 3080 4719 3081 4720
rect 3077 4721 3078 4722
rect 3145 4721 3146 4722
rect 2903 4723 2904 4724
rect 3146 4723 3147 4724
rect 3083 4725 3084 4726
rect 3108 4725 3109 4726
rect 3090 4727 3091 4728
rect 3107 4727 3108 4728
rect 3122 4727 3123 4728
rect 3181 4727 3182 4728
rect 2933 4729 2934 4730
rect 3182 4729 3183 4730
rect 3135 4731 3136 4732
rect 3217 4731 3218 4732
rect 3120 4733 3121 4734
rect 3134 4733 3135 4734
rect 3119 4735 3120 4736
rect 3178 4735 3179 4736
rect 3139 4737 3140 4738
rect 3520 4737 3521 4738
rect 3126 4739 3127 4740
rect 3140 4739 3141 4740
rect 3096 4741 3097 4742
rect 3125 4741 3126 4742
rect 3154 4741 3155 4742
rect 3490 4741 3491 4742
rect 3158 4743 3159 4744
rect 3205 4743 3206 4744
rect 3170 4745 3171 4746
rect 3433 4745 3434 4746
rect 3176 4747 3177 4748
rect 3241 4747 3242 4748
rect 3188 4749 3189 4750
rect 3229 4749 3230 4750
rect 3190 4751 3191 4752
rect 3197 4751 3198 4752
rect 3194 4753 3195 4754
rect 3265 4753 3266 4754
rect 3036 4755 3037 4756
rect 3266 4755 3267 4756
rect 3037 4757 3038 4758
rect 3344 4757 3345 4758
rect 3203 4759 3204 4760
rect 3280 4759 3281 4760
rect 3209 4761 3210 4762
rect 3253 4761 3254 4762
rect 3215 4763 3216 4764
rect 3292 4763 3293 4764
rect 3027 4765 3028 4766
rect 3293 4765 3294 4766
rect 3027 4767 3028 4768
rect 3286 4767 3287 4768
rect 3223 4769 3224 4770
rect 3458 4769 3459 4770
rect 3230 4771 3231 4772
rect 3502 4771 3503 4772
rect 3233 4773 3234 4774
rect 3304 4773 3305 4774
rect 2957 4775 2958 4776
rect 3305 4775 3306 4776
rect 3245 4777 3246 4778
rect 3340 4777 3341 4778
rect 3247 4779 3248 4780
rect 3380 4779 3381 4780
rect 3251 4781 3252 4782
rect 3334 4781 3335 4782
rect 3257 4783 3258 4784
rect 3358 4783 3359 4784
rect 3268 4785 3269 4786
rect 3772 4785 3773 4786
rect 3269 4787 3270 4788
rect 3352 4787 3353 4788
rect 3274 4789 3275 4790
rect 3750 4789 3751 4790
rect 3275 4791 3276 4792
rect 3382 4791 3383 4792
rect 3281 4793 3282 4794
rect 3370 4793 3371 4794
rect 3132 4795 3133 4796
rect 3371 4795 3372 4796
rect 2886 4797 2887 4798
rect 3131 4797 3132 4798
rect 3295 4797 3296 4798
rect 3308 4797 3309 4798
rect 3302 4799 3303 4800
rect 3391 4799 3392 4800
rect 3310 4801 3311 4802
rect 3398 4801 3399 4802
rect 3311 4803 3312 4804
rect 3442 4803 3443 4804
rect 3314 4805 3315 4806
rect 3445 4805 3446 4806
rect 3317 4807 3318 4808
rect 3406 4807 3407 4808
rect 3320 4809 3321 4810
rect 3409 4809 3410 4810
rect 3322 4811 3323 4812
rect 3599 4811 3600 4812
rect 3199 4813 3200 4814
rect 3323 4813 3324 4814
rect 3335 4813 3336 4814
rect 3466 4813 3467 4814
rect 3338 4815 3339 4816
rect 3469 4815 3470 4816
rect 3341 4817 3342 4818
rect 3430 4817 3431 4818
rect 3347 4819 3348 4820
rect 3412 4819 3413 4820
rect 3353 4821 3354 4822
rect 3484 4821 3485 4822
rect 3356 4823 3357 4824
rect 3418 4823 3419 4824
rect 3362 4825 3363 4826
rect 3493 4825 3494 4826
rect 3374 4827 3375 4828
rect 3505 4827 3506 4828
rect 3377 4829 3378 4830
rect 3772 4829 3773 4830
rect 3386 4831 3387 4832
rect 3517 4831 3518 4832
rect 3388 4833 3389 4834
rect 3739 4833 3740 4834
rect 3142 4835 3143 4836
rect 3389 4835 3390 4836
rect 3404 4835 3405 4836
rect 3671 4835 3672 4836
rect 3416 4837 3417 4838
rect 3424 4837 3425 4838
rect 3422 4839 3423 4840
rect 3553 4839 3554 4840
rect 3428 4841 3429 4842
rect 3472 4841 3473 4842
rect 3431 4843 3432 4844
rect 3481 4843 3482 4844
rect 3434 4845 3435 4846
rect 3535 4845 3536 4846
rect 3446 4847 3447 4848
rect 3454 4847 3455 4848
rect 3452 4849 3453 4850
rect 3896 4849 3897 4850
rect 3460 4851 3461 4852
rect 3699 4851 3700 4852
rect 3464 4853 3465 4854
rect 3583 4853 3584 4854
rect 3476 4855 3477 4856
rect 3939 4855 3940 4856
rect 3482 4857 3483 4858
rect 3571 4857 3572 4858
rect 3494 4859 3495 4860
rect 3589 4859 3590 4860
rect 3506 4861 3507 4862
rect 3595 4861 3596 4862
rect 3523 4863 3524 4864
rect 3775 4863 3776 4864
rect 3524 4865 3525 4866
rect 3631 4865 3632 4866
rect 3532 4867 3533 4868
rect 3659 4867 3660 4868
rect 3536 4869 3537 4870
rect 3649 4869 3650 4870
rect 3542 4871 3543 4872
rect 3655 4871 3656 4872
rect 3529 4873 3530 4874
rect 3656 4873 3657 4874
rect 3530 4875 3531 4876
rect 3625 4875 3626 4876
rect 3547 4877 3548 4878
rect 3596 4877 3597 4878
rect 3548 4879 3549 4880
rect 3661 4879 3662 4880
rect 3554 4881 3555 4882
rect 3673 4881 3674 4882
rect 3556 4883 3557 4884
rect 3593 4883 3594 4884
rect 3367 4885 3368 4886
rect 3557 4885 3558 4886
rect 3368 4887 3369 4888
rect 3499 4887 3500 4888
rect 3500 4889 3501 4890
rect 3559 4889 3560 4890
rect 3262 4891 3263 4892
rect 3560 4891 3561 4892
rect 3263 4893 3264 4894
rect 3328 4893 3329 4894
rect 3329 4895 3330 4896
rect 3400 4895 3401 4896
rect 3401 4897 3402 4898
rect 3487 4897 3488 4898
rect 3488 4899 3489 4900
rect 3601 4899 3602 4900
rect 3563 4901 3564 4902
rect 3667 4901 3668 4902
rect 3364 4903 3365 4904
rect 3668 4903 3669 4904
rect 3565 4905 3566 4906
rect 3782 4905 3783 4906
rect 3569 4907 3570 4908
rect 3853 4907 3854 4908
rect 3577 4909 3578 4910
rect 3893 4909 3894 4910
rect 3587 4911 3588 4912
rect 3685 4911 3686 4912
rect 3605 4913 3606 4914
rect 3709 4913 3710 4914
rect 3478 4915 3479 4916
rect 3708 4915 3709 4916
rect 3611 4917 3612 4918
rect 3775 4917 3776 4918
rect 3623 4919 3624 4920
rect 3960 4919 3961 4920
rect 3629 4921 3630 4922
rect 3733 4921 3734 4922
rect 3632 4923 3633 4924
rect 3769 4923 3770 4924
rect 3511 4925 3512 4926
rect 3768 4925 3769 4926
rect 3512 4927 3513 4928
rect 3613 4927 3614 4928
rect 3638 4927 3639 4928
rect 3697 4927 3698 4928
rect 3644 4929 3645 4930
rect 3900 4929 3901 4930
rect 3581 4931 3582 4932
rect 3899 4931 3900 4932
rect 3662 4933 3663 4934
rect 3703 4933 3704 4934
rect 3665 4935 3666 4936
rect 3706 4935 3707 4936
rect 3678 4937 3679 4938
rect 3846 4937 3847 4938
rect 3682 4939 3683 4940
rect 3932 4939 3933 4940
rect 3691 4941 3692 4942
rect 3839 4941 3840 4942
rect 3693 4943 3694 4944
rect 3983 4943 3984 4944
rect 3696 4945 3697 4946
rect 3754 4945 3755 4946
rect 3702 4947 3703 4948
rect 3928 4947 3929 4948
rect 3715 4949 3716 4950
rect 3832 4949 3833 4950
rect 3714 4951 3715 4952
rect 3760 4951 3761 4952
rect 3717 4953 3718 4954
rect 3903 4953 3904 4954
rect 3726 4955 3727 4956
rect 3766 4955 3767 4956
rect 3419 4957 3420 4958
rect 3765 4957 3766 4958
rect 3738 4959 3739 4960
rect 3787 4959 3788 4960
rect 3741 4961 3742 4962
rect 3790 4961 3791 4962
rect 3744 4963 3745 4964
rect 3863 4963 3864 4964
rect 3757 4965 3758 4966
rect 3828 4965 3829 4966
rect 3759 4967 3760 4968
rect 3922 4967 3923 4968
rect 3763 4969 3764 4970
rect 3835 4969 3836 4970
rect 3762 4971 3763 4972
rect 3793 4971 3794 4972
rect 3779 4973 3780 4974
rect 3886 4973 3887 4974
rect 3797 4975 3798 4976
rect 3893 4975 3894 4976
rect 3800 4977 3801 4978
rect 3902 4977 3903 4978
rect 3803 4979 3804 4980
rect 3844 4979 3845 4980
rect 3805 4981 3806 4982
rect 3909 4981 3910 4982
rect 3808 4983 3809 4984
rect 3970 4983 3971 4984
rect 3809 4985 3810 4986
rect 3856 4985 3857 4986
rect 3812 4987 3813 4988
rect 3859 4987 3860 4988
rect 3821 4989 3822 4990
rect 3874 4989 3875 4990
rect 3824 4991 3825 4992
rect 3877 4991 3878 4992
rect 3833 4993 3834 4994
rect 3880 4993 3881 4994
rect 3836 4995 3837 4996
rect 3883 4995 3884 4996
rect 3729 4997 3730 4998
rect 3882 4997 3883 4998
rect 3850 4999 3851 5000
rect 3896 4999 3897 5000
rect 3866 5001 3867 5002
rect 3913 5001 3914 5002
rect 3784 5003 3785 5004
rect 3912 5003 3913 5004
rect 3747 5005 3748 5006
rect 3785 5005 3786 5006
rect 3869 5005 3870 5006
rect 3916 5005 3917 5006
rect 3889 5007 3890 5008
rect 3919 5007 3920 5008
rect 3935 5007 3936 5008
rect 3967 5007 3968 5008
rect 2863 5016 2864 5017
rect 2876 5016 2877 5017
rect 2870 5018 2871 5019
rect 3009 5018 3010 5019
rect 2873 5020 2874 5021
rect 3047 5020 3048 5021
rect 2879 5022 2880 5023
rect 3194 5022 3195 5023
rect 2882 5024 2883 5025
rect 3012 5024 3013 5025
rect 2896 5026 2897 5027
rect 3131 5026 3132 5027
rect 2905 5028 2906 5029
rect 3275 5028 3276 5029
rect 2912 5030 2913 5031
rect 3146 5030 3147 5031
rect 2922 5032 2923 5033
rect 3149 5032 3150 5033
rect 2922 5034 2923 5035
rect 3278 5034 3279 5035
rect 2919 5036 2920 5037
rect 3279 5036 3280 5037
rect 2929 5038 2930 5039
rect 3335 5038 3336 5039
rect 2933 5040 2934 5041
rect 3069 5040 3070 5041
rect 2940 5042 2941 5043
rect 3311 5042 3312 5043
rect 2941 5044 2942 5045
rect 2950 5044 2951 5045
rect 2947 5046 2948 5047
rect 3263 5046 3264 5047
rect 2960 5048 2961 5049
rect 3386 5048 3387 5049
rect 2973 5050 2974 5051
rect 3221 5050 3222 5051
rect 2972 5052 2973 5053
rect 3192 5052 3193 5053
rect 2988 5054 2989 5055
rect 2991 5054 2992 5055
rect 2994 5054 2995 5055
rect 2997 5054 2998 5055
rect 3000 5054 3001 5055
rect 3308 5054 3309 5055
rect 3003 5056 3004 5057
rect 3317 5056 3318 5057
rect 3006 5058 3007 5059
rect 3027 5058 3028 5059
rect 3012 5060 3013 5061
rect 3021 5060 3022 5061
rect 3021 5062 3022 5063
rect 3125 5062 3126 5063
rect 3037 5064 3038 5065
rect 3164 5064 3165 5065
rect 3041 5066 3042 5067
rect 3140 5066 3141 5067
rect 2893 5068 2894 5069
rect 3141 5068 3142 5069
rect 3018 5070 3019 5071
rect 3042 5070 3043 5071
rect 3044 5070 3045 5071
rect 3071 5070 3072 5071
rect 3048 5072 3049 5073
rect 3107 5072 3108 5073
rect 3057 5074 3058 5075
rect 3269 5074 3270 5075
rect 2979 5076 2980 5077
rect 3270 5076 3271 5077
rect 3060 5078 3061 5079
rect 3065 5078 3066 5079
rect 3066 5080 3067 5081
rect 3080 5080 3081 5081
rect 3077 5082 3078 5083
rect 3114 5082 3115 5083
rect 3078 5084 3079 5085
rect 3083 5084 3084 5085
rect 3102 5084 3103 5085
rect 3134 5084 3135 5085
rect 3119 5086 3120 5087
rect 3129 5086 3130 5087
rect 3122 5088 3123 5089
rect 3132 5088 3133 5089
rect 3156 5088 3157 5089
rect 3170 5088 3171 5089
rect 3158 5090 3159 5091
rect 3162 5090 3163 5091
rect 3168 5090 3169 5091
rect 3197 5090 3198 5091
rect 3180 5092 3181 5093
rect 3182 5092 3183 5093
rect 3183 5094 3184 5095
rect 3266 5094 3267 5095
rect 3198 5096 3199 5097
rect 3458 5096 3459 5097
rect 3203 5098 3204 5099
rect 3240 5098 3241 5099
rect 3108 5100 3109 5101
rect 3204 5100 3205 5101
rect 3219 5100 3220 5101
rect 3320 5100 3321 5101
rect 3222 5102 3223 5103
rect 3371 5102 3372 5103
rect 3227 5104 3228 5105
rect 3372 5104 3373 5105
rect 3231 5106 3232 5107
rect 3560 5106 3561 5107
rect 3233 5108 3234 5109
rect 3273 5108 3274 5109
rect 3030 5110 3031 5111
rect 3234 5110 3235 5111
rect 3030 5112 3031 5113
rect 3096 5112 3097 5113
rect 3243 5112 3244 5113
rect 3314 5112 3315 5113
rect 3245 5114 3246 5115
rect 3675 5114 3676 5115
rect 3246 5116 3247 5117
rect 3380 5116 3381 5117
rect 3249 5118 3250 5119
rect 3389 5118 3390 5119
rect 3251 5120 3252 5121
rect 3291 5120 3292 5121
rect 3215 5122 3216 5123
rect 3252 5122 3253 5123
rect 3209 5124 3210 5125
rect 3216 5124 3217 5125
rect 3176 5126 3177 5127
rect 3210 5126 3211 5127
rect 3257 5126 3258 5127
rect 3309 5126 3310 5127
rect 3260 5128 3261 5129
rect 3312 5128 3313 5129
rect 3281 5130 3282 5131
rect 3321 5130 3322 5131
rect 2919 5132 2920 5133
rect 3282 5132 3283 5133
rect 3297 5132 3298 5133
rect 3404 5132 3405 5133
rect 3299 5134 3300 5135
rect 3315 5134 3316 5135
rect 3300 5136 3301 5137
rect 3557 5136 3558 5137
rect 3302 5138 3303 5139
rect 3318 5138 3319 5139
rect 3293 5140 3294 5141
rect 3303 5140 3304 5141
rect 3323 5140 3324 5141
rect 3722 5140 3723 5141
rect 3324 5142 3325 5143
rect 3338 5142 3339 5143
rect 3327 5144 3328 5145
rect 3599 5144 3600 5145
rect 3333 5146 3334 5147
rect 3446 5146 3447 5147
rect 3339 5148 3340 5149
rect 3347 5148 3348 5149
rect 3188 5150 3189 5151
rect 3348 5150 3349 5151
rect 3344 5152 3345 5153
rect 3360 5152 3361 5153
rect 3305 5154 3306 5155
rect 3345 5154 3346 5155
rect 3351 5154 3352 5155
rect 3356 5154 3357 5155
rect 3329 5156 3330 5157
rect 3357 5156 3358 5157
rect 3353 5158 3354 5159
rect 3393 5158 3394 5159
rect 3362 5160 3363 5161
rect 3408 5160 3409 5161
rect 3363 5162 3364 5163
rect 3659 5162 3660 5163
rect 3368 5164 3369 5165
rect 3678 5164 3679 5165
rect 3369 5166 3370 5167
rect 3431 5166 3432 5167
rect 3374 5168 3375 5169
rect 3414 5168 3415 5169
rect 3381 5170 3382 5171
rect 3611 5170 3612 5171
rect 3387 5172 3388 5173
rect 3782 5172 3783 5173
rect 3398 5174 3399 5175
rect 3432 5174 3433 5175
rect 3401 5176 3402 5177
rect 3429 5176 3430 5177
rect 3416 5178 3417 5179
rect 3636 5178 3637 5179
rect 3377 5180 3378 5181
rect 3417 5180 3418 5181
rect 3419 5180 3420 5181
rect 3426 5180 3427 5181
rect 3420 5182 3421 5183
rect 3817 5182 3818 5183
rect 3434 5184 3435 5185
rect 3459 5184 3460 5185
rect 3438 5186 3439 5187
rect 3775 5186 3776 5187
rect 3447 5188 3448 5189
rect 3708 5188 3709 5189
rect 3450 5190 3451 5191
rect 3656 5190 3657 5191
rect 3468 5192 3469 5193
rect 3842 5192 3843 5193
rect 3471 5194 3472 5195
rect 3665 5194 3666 5195
rect 3480 5196 3481 5197
rect 3662 5196 3663 5197
rect 3488 5198 3489 5199
rect 3519 5198 3520 5199
rect 3489 5200 3490 5201
rect 3711 5200 3712 5201
rect 3435 5202 3436 5203
rect 3711 5202 3712 5203
rect 3530 5204 3531 5205
rect 3779 5204 3780 5205
rect 3512 5206 3513 5207
rect 3531 5206 3532 5207
rect 3542 5206 3543 5207
rect 3561 5206 3562 5207
rect 3543 5208 3544 5209
rect 3838 5208 3839 5209
rect 3554 5210 3555 5211
rect 3585 5210 3586 5211
rect 3536 5212 3537 5213
rect 3555 5212 3556 5213
rect 3537 5214 3538 5215
rect 3638 5214 3639 5215
rect 3563 5216 3564 5217
rect 3579 5216 3580 5217
rect 3581 5216 3582 5217
rect 3768 5216 3769 5217
rect 3587 5218 3588 5219
rect 3687 5218 3688 5219
rect 3593 5220 3594 5221
rect 3671 5220 3672 5221
rect 3569 5222 3570 5223
rect 3594 5222 3595 5223
rect 3612 5222 3613 5223
rect 3747 5222 3748 5223
rect 3623 5224 3624 5225
rect 3902 5224 3903 5225
rect 3605 5226 3606 5227
rect 3624 5226 3625 5227
rect 3629 5226 3630 5227
rect 3648 5226 3649 5227
rect 3632 5228 3633 5229
rect 3875 5228 3876 5229
rect 3642 5230 3643 5231
rect 3702 5230 3703 5231
rect 3657 5232 3658 5233
rect 3714 5232 3715 5233
rect 3422 5234 3423 5235
rect 3715 5234 3716 5235
rect 3660 5236 3661 5237
rect 3831 5236 3832 5237
rect 3669 5238 3670 5239
rect 3726 5238 3727 5239
rect 3672 5240 3673 5241
rect 3729 5240 3730 5241
rect 3500 5242 3501 5243
rect 3729 5242 3730 5243
rect 3464 5244 3465 5245
rect 3501 5244 3502 5245
rect 3465 5246 3466 5247
rect 3596 5246 3597 5247
rect 3675 5246 3676 5247
rect 3696 5246 3697 5247
rect 3678 5248 3679 5249
rect 3732 5248 3733 5249
rect 3681 5250 3682 5251
rect 3744 5250 3745 5251
rect 3684 5252 3685 5253
rect 3741 5252 3742 5253
rect 3693 5254 3694 5255
rect 3912 5254 3913 5255
rect 3699 5256 3700 5257
rect 3772 5256 3773 5257
rect 3702 5258 3703 5259
rect 3759 5258 3760 5259
rect 3705 5260 3706 5261
rect 3762 5260 3763 5261
rect 3717 5262 3718 5263
rect 3863 5262 3864 5263
rect 3441 5264 3442 5265
rect 3718 5264 3719 5265
rect 3725 5264 3726 5265
rect 3806 5264 3807 5265
rect 3735 5266 3736 5267
rect 3785 5266 3786 5267
rect 3738 5268 3739 5269
rect 3853 5268 3854 5269
rect 3747 5270 3748 5271
rect 3797 5270 3798 5271
rect 3644 5272 3645 5273
rect 3796 5272 3797 5273
rect 3750 5274 3751 5275
rect 3800 5274 3801 5275
rect 3588 5276 3589 5277
rect 3799 5276 3800 5277
rect 3753 5278 3754 5279
rect 3869 5278 3870 5279
rect 3759 5280 3760 5281
rect 3803 5280 3804 5281
rect 3567 5282 3568 5283
rect 3803 5282 3804 5283
rect 3765 5284 3766 5285
rect 3821 5284 3822 5285
rect 3630 5286 3631 5287
rect 3820 5286 3821 5287
rect 3771 5288 3772 5289
rect 3809 5288 3810 5289
rect 3476 5290 3477 5291
rect 3810 5290 3811 5291
rect 3477 5292 3478 5293
rect 3482 5292 3483 5293
rect 3452 5294 3453 5295
rect 3483 5294 3484 5295
rect 3453 5296 3454 5297
rect 3494 5296 3495 5297
rect 3495 5298 3496 5299
rect 3506 5298 3507 5299
rect 3507 5300 3508 5301
rect 3856 5300 3857 5301
rect 3774 5302 3775 5303
rect 3846 5302 3847 5303
rect 3756 5304 3757 5305
rect 3845 5304 3846 5305
rect 3783 5306 3784 5307
rect 3833 5306 3834 5307
rect 3786 5308 3787 5309
rect 3836 5308 3837 5309
rect 3812 5310 3813 5311
rect 3849 5310 3850 5311
rect 3341 5312 3342 5313
rect 3813 5312 3814 5313
rect 3824 5312 3825 5313
rect 3896 5312 3897 5313
rect 3827 5314 3828 5315
rect 3866 5314 3867 5315
rect 3834 5316 3835 5317
rect 3889 5316 3890 5317
rect 2884 5325 2885 5326
rect 3270 5325 3271 5326
rect 2888 5327 2889 5328
rect 3141 5327 3142 5328
rect 2891 5329 2892 5330
rect 2895 5329 2896 5330
rect 2908 5329 2909 5330
rect 3210 5329 3211 5330
rect 2912 5331 2913 5332
rect 2922 5331 2923 5332
rect 2911 5333 2912 5334
rect 3129 5333 3130 5334
rect 2929 5335 2930 5336
rect 2934 5335 2935 5336
rect 2941 5335 2942 5336
rect 3211 5335 3212 5336
rect 2945 5337 2946 5338
rect 3180 5337 3181 5338
rect 2965 5339 2966 5340
rect 3229 5339 3230 5340
rect 2969 5341 2970 5342
rect 3042 5341 3043 5342
rect 2972 5343 2973 5344
rect 3348 5343 3349 5344
rect 2975 5345 2976 5346
rect 3102 5345 3103 5346
rect 2979 5347 2980 5348
rect 3765 5347 3766 5348
rect 2984 5349 2985 5350
rect 2988 5349 2989 5350
rect 2990 5349 2991 5350
rect 2994 5349 2995 5350
rect 2996 5349 2997 5350
rect 3048 5349 3049 5350
rect 2999 5351 3000 5352
rect 3042 5351 3043 5352
rect 3003 5353 3004 5354
rect 3381 5353 3382 5354
rect 3008 5355 3009 5356
rect 3012 5355 3013 5356
rect 3018 5355 3019 5356
rect 3318 5355 3319 5356
rect 3021 5357 3022 5358
rect 3268 5357 3269 5358
rect 3020 5359 3021 5360
rect 3114 5359 3115 5360
rect 3023 5361 3024 5362
rect 3096 5361 3097 5362
rect 3030 5363 3031 5364
rect 3360 5363 3361 5364
rect 3030 5365 3031 5366
rect 3187 5365 3188 5366
rect 3036 5367 3037 5368
rect 3060 5367 3061 5368
rect 3048 5369 3049 5370
rect 3066 5369 3067 5370
rect 3054 5371 3055 5372
rect 3385 5371 3386 5372
rect 3054 5373 3055 5374
rect 3078 5373 3079 5374
rect 3069 5375 3070 5376
rect 3208 5375 3209 5376
rect 3072 5377 3073 5378
rect 3286 5377 3287 5378
rect 3075 5379 3076 5380
rect 3417 5379 3418 5380
rect 3099 5381 3100 5382
rect 3400 5381 3401 5382
rect 3106 5383 3107 5384
rect 3175 5383 3176 5384
rect 3111 5385 3112 5386
rect 3369 5385 3370 5386
rect 3115 5387 3116 5388
rect 3204 5387 3205 5388
rect 2922 5389 2923 5390
rect 3205 5389 3206 5390
rect 3121 5391 3122 5392
rect 3162 5391 3163 5392
rect 3132 5393 3133 5394
rect 3178 5393 3179 5394
rect 3144 5395 3145 5396
rect 3357 5395 3358 5396
rect 3145 5397 3146 5398
rect 3168 5397 3169 5398
rect 3147 5399 3148 5400
rect 3781 5399 3782 5400
rect 3151 5401 3152 5402
rect 3240 5401 3241 5402
rect 2960 5403 2961 5404
rect 3241 5403 3242 5404
rect 3154 5405 3155 5406
rect 3243 5405 3244 5406
rect 3160 5407 3161 5408
rect 3219 5407 3220 5408
rect 3163 5409 3164 5410
rect 3252 5409 3253 5410
rect 3169 5411 3170 5412
rect 3279 5411 3280 5412
rect 3172 5413 3173 5414
rect 3282 5413 3283 5414
rect 3057 5415 3058 5416
rect 3283 5415 3284 5416
rect 3181 5417 3182 5418
rect 3309 5417 3310 5418
rect 3156 5419 3157 5420
rect 3310 5419 3311 5420
rect 3157 5421 3158 5422
rect 3216 5421 3217 5422
rect 3183 5423 3184 5424
rect 3214 5423 3215 5424
rect 3184 5425 3185 5426
rect 3312 5425 3313 5426
rect 3192 5427 3193 5428
rect 3244 5427 3245 5428
rect 3193 5429 3194 5430
rect 3234 5429 3235 5430
rect 3217 5431 3218 5432
rect 3321 5431 3322 5432
rect 3220 5433 3221 5434
rect 3324 5433 3325 5434
rect 3226 5435 3227 5436
rect 3514 5435 3515 5436
rect 3235 5437 3236 5438
rect 3345 5437 3346 5438
rect 3246 5439 3247 5440
rect 3319 5439 3320 5440
rect 3247 5441 3248 5442
rect 3393 5441 3394 5442
rect 3249 5443 3250 5444
rect 3397 5443 3398 5444
rect 3033 5445 3034 5446
rect 3250 5445 3251 5446
rect 3253 5445 3254 5446
rect 3291 5445 3292 5446
rect 3259 5447 3260 5448
rect 3303 5447 3304 5448
rect 3265 5449 3266 5450
rect 3315 5449 3316 5450
rect 3271 5451 3272 5452
rect 3414 5451 3415 5452
rect 3277 5453 3278 5454
rect 3408 5453 3409 5454
rect 3289 5455 3290 5456
rect 3333 5455 3334 5456
rect 3295 5457 3296 5458
rect 3429 5457 3430 5458
rect 3300 5459 3301 5460
rect 3610 5459 3611 5460
rect 3313 5461 3314 5462
rect 3690 5461 3691 5462
rect 3325 5463 3326 5464
rect 3351 5463 3352 5464
rect 3331 5465 3332 5466
rect 3447 5465 3448 5466
rect 3337 5467 3338 5468
rect 3426 5467 3427 5468
rect 3339 5469 3340 5470
rect 3349 5469 3350 5470
rect 3355 5469 3356 5470
rect 3489 5469 3490 5470
rect 3361 5471 3362 5472
rect 3459 5471 3460 5472
rect 3363 5473 3364 5474
rect 3622 5473 3623 5474
rect 3367 5475 3368 5476
rect 3483 5475 3484 5476
rect 3391 5477 3392 5478
rect 3501 5477 3502 5478
rect 3297 5479 3298 5480
rect 3502 5479 3503 5480
rect 3409 5481 3410 5482
rect 3519 5481 3520 5482
rect 3424 5483 3425 5484
rect 3432 5483 3433 5484
rect 3433 5485 3434 5486
rect 3507 5485 3508 5486
rect 3435 5487 3436 5488
rect 3655 5487 3656 5488
rect 3450 5489 3451 5490
rect 3743 5489 3744 5490
rect 3451 5491 3452 5492
rect 3531 5491 3532 5492
rect 3453 5493 3454 5494
rect 3553 5493 3554 5494
rect 3463 5495 3464 5496
rect 3549 5495 3550 5496
rect 3441 5497 3442 5498
rect 3550 5497 3551 5498
rect 3465 5499 3466 5500
rect 3634 5499 3635 5500
rect 3471 5501 3472 5502
rect 3732 5501 3733 5502
rect 3475 5503 3476 5504
rect 3555 5503 3556 5504
rect 3420 5505 3421 5506
rect 3556 5505 3557 5506
rect 3421 5507 3422 5508
rect 3718 5507 3719 5508
rect 3480 5509 3481 5510
rect 3799 5509 3800 5510
rect 3481 5511 3482 5512
rect 3874 5511 3875 5512
rect 3487 5513 3488 5514
rect 3585 5513 3586 5514
rect 3490 5515 3491 5516
rect 3561 5515 3562 5516
rect 3495 5517 3496 5518
rect 3792 5517 3793 5518
rect 3387 5519 3388 5520
rect 3496 5519 3497 5520
rect 3372 5521 3373 5522
rect 3388 5521 3389 5522
rect 3373 5523 3374 5524
rect 3715 5523 3716 5524
rect 3508 5525 3509 5526
rect 3525 5525 3526 5526
rect 3532 5525 3533 5526
rect 3750 5525 3751 5526
rect 3343 5527 3344 5528
rect 3750 5527 3751 5528
rect 3535 5529 3536 5530
rect 3594 5529 3595 5530
rect 3541 5531 3542 5532
rect 3852 5531 3853 5532
rect 3562 5533 3563 5534
rect 3789 5533 3790 5534
rect 3567 5535 3568 5536
rect 3871 5535 3872 5536
rect 3198 5537 3199 5538
rect 3568 5537 3569 5538
rect 3199 5539 3200 5540
rect 3273 5539 3274 5540
rect 3574 5539 3575 5540
rect 3834 5539 3835 5540
rect 3583 5541 3584 5542
rect 3636 5541 3637 5542
rect 3588 5543 3589 5544
rect 3598 5543 3599 5544
rect 3624 5543 3625 5544
rect 3853 5543 3854 5544
rect 3327 5545 3328 5546
rect 3625 5545 3626 5546
rect 3628 5545 3629 5546
rect 3884 5545 3885 5546
rect 3642 5547 3643 5548
rect 3878 5547 3879 5548
rect 3612 5549 3613 5550
rect 3643 5549 3644 5550
rect 3231 5551 3232 5552
rect 3613 5551 3614 5552
rect 3648 5551 3649 5552
rect 3841 5551 3842 5552
rect 3301 5553 3302 5554
rect 3649 5553 3650 5554
rect 3657 5553 3658 5554
rect 3692 5553 3693 5554
rect 3438 5555 3439 5556
rect 3658 5555 3659 5556
rect 3660 5555 3661 5556
rect 3835 5555 3836 5556
rect 3661 5557 3662 5558
rect 3820 5557 3821 5558
rect 3537 5559 3538 5560
rect 3821 5559 3822 5560
rect 3538 5561 3539 5562
rect 3768 5561 3769 5562
rect 3672 5563 3673 5564
rect 3689 5563 3690 5564
rect 3675 5565 3676 5566
rect 3737 5565 3738 5566
rect 3678 5567 3679 5568
rect 3707 5567 3708 5568
rect 3681 5569 3682 5570
rect 3698 5569 3699 5570
rect 3684 5571 3685 5572
rect 3713 5571 3714 5572
rect 3687 5573 3688 5574
rect 3716 5573 3717 5574
rect 3669 5575 3670 5576
rect 3686 5575 3687 5576
rect 3695 5575 3696 5576
rect 3832 5575 3833 5576
rect 3705 5577 3706 5578
rect 3725 5577 3726 5578
rect 3735 5577 3736 5578
rect 3857 5577 3858 5578
rect 3747 5579 3748 5580
rect 3845 5579 3846 5580
rect 3415 5581 3416 5582
rect 3746 5581 3747 5582
rect 3753 5581 3754 5582
rect 3769 5581 3770 5582
rect 3756 5583 3757 5584
rect 3763 5583 3764 5584
rect 3427 5585 3428 5586
rect 3757 5585 3758 5586
rect 3771 5585 3772 5586
rect 3793 5585 3794 5586
rect 3774 5587 3775 5588
rect 3796 5587 3797 5588
rect 3477 5589 3478 5590
rect 3775 5589 3776 5590
rect 3778 5589 3779 5590
rect 3811 5589 3812 5590
rect 3783 5591 3784 5592
rect 3805 5591 3806 5592
rect 3702 5593 3703 5594
rect 3784 5593 3785 5594
rect 3701 5595 3702 5596
rect 3861 5595 3862 5596
rect 3786 5597 3787 5598
rect 3808 5597 3809 5598
rect 3759 5599 3760 5600
rect 3787 5599 3788 5600
rect 3307 5601 3308 5602
rect 3760 5601 3761 5602
rect 3824 5601 3825 5602
rect 3847 5601 3848 5602
rect 3630 5603 3631 5604
rect 3825 5603 3826 5604
rect 3468 5605 3469 5606
rect 3631 5605 3632 5606
rect 3469 5607 3470 5608
rect 3677 5607 3678 5608
rect 3827 5607 3828 5608
rect 3844 5607 3845 5608
rect 3867 5607 3868 5608
rect 3887 5607 3888 5608
rect 3543 5609 3544 5610
rect 3867 5609 3868 5610
rect 3544 5611 3545 5612
rect 3579 5611 3580 5612
rect 3580 5613 3581 5614
rect 3817 5613 3818 5614
rect 3740 5615 3741 5616
rect 3818 5615 3819 5616
rect 2904 5624 2905 5625
rect 3358 5624 3359 5625
rect 2905 5626 2906 5627
rect 3778 5626 3779 5627
rect 2908 5628 2909 5629
rect 3178 5628 3179 5629
rect 2915 5630 2916 5631
rect 3214 5630 3215 5631
rect 2922 5632 2923 5633
rect 3184 5632 3185 5633
rect 2937 5634 2938 5635
rect 2951 5634 2952 5635
rect 2929 5636 2930 5637
rect 2938 5636 2939 5637
rect 2941 5636 2942 5637
rect 3295 5636 3296 5637
rect 2944 5638 2945 5639
rect 3172 5638 3173 5639
rect 2947 5640 2948 5641
rect 3418 5640 3419 5641
rect 2953 5642 2954 5643
rect 3217 5642 3218 5643
rect 2956 5644 2957 5645
rect 3127 5644 3128 5645
rect 2965 5646 2966 5647
rect 3298 5646 3299 5647
rect 2972 5648 2973 5649
rect 2996 5648 2997 5649
rect 2975 5650 2976 5651
rect 3442 5650 3443 5651
rect 2975 5652 2976 5653
rect 3205 5652 3206 5653
rect 2984 5654 2985 5655
rect 3148 5654 3149 5655
rect 2984 5656 2985 5657
rect 2990 5656 2991 5657
rect 2990 5658 2991 5659
rect 3133 5658 3134 5659
rect 3002 5660 3003 5661
rect 3008 5660 3009 5661
rect 3008 5662 3009 5663
rect 3262 5662 3263 5663
rect 3015 5664 3016 5665
rect 3346 5664 3347 5665
rect 3020 5666 3021 5667
rect 3094 5666 3095 5667
rect 3021 5668 3022 5669
rect 3042 5668 3043 5669
rect 3023 5670 3024 5671
rect 3193 5670 3194 5671
rect 3026 5672 3027 5673
rect 3217 5672 3218 5673
rect 3030 5674 3031 5675
rect 3283 5674 3284 5675
rect 3033 5676 3034 5677
rect 3472 5676 3473 5677
rect 3048 5678 3049 5679
rect 3070 5678 3071 5679
rect 3048 5680 3049 5681
rect 3490 5680 3491 5681
rect 3054 5682 3055 5683
rect 3082 5682 3083 5683
rect 3106 5682 3107 5683
rect 3220 5682 3221 5683
rect 3157 5684 3158 5685
rect 3193 5684 3194 5685
rect 3145 5686 3146 5687
rect 3157 5686 3158 5687
rect 3121 5688 3122 5689
rect 3145 5688 3146 5689
rect 3076 5690 3077 5691
rect 3121 5690 3122 5691
rect 3169 5690 3170 5691
rect 3295 5690 3296 5691
rect 3175 5692 3176 5693
rect 3340 5692 3341 5693
rect 3181 5694 3182 5695
rect 3370 5694 3371 5695
rect 3115 5696 3116 5697
rect 3181 5696 3182 5697
rect 3199 5696 3200 5697
rect 3256 5696 3257 5697
rect 3103 5698 3104 5699
rect 3199 5698 3200 5699
rect 3079 5700 3080 5701
rect 3103 5700 3104 5701
rect 3202 5700 3203 5701
rect 3421 5700 3422 5701
rect 3154 5702 3155 5703
rect 3421 5702 3422 5703
rect 3205 5704 3206 5705
rect 3568 5704 3569 5705
rect 3208 5706 3209 5707
rect 3403 5706 3404 5707
rect 3226 5708 3227 5709
rect 3670 5708 3671 5709
rect 3229 5710 3230 5711
rect 3430 5710 3431 5711
rect 3151 5712 3152 5713
rect 3229 5712 3230 5713
rect 3235 5712 3236 5713
rect 3406 5712 3407 5713
rect 3235 5714 3236 5715
rect 3385 5714 3386 5715
rect 3250 5716 3251 5717
rect 3499 5716 3500 5717
rect 3268 5718 3269 5719
rect 3316 5718 3317 5719
rect 2888 5720 2889 5721
rect 3268 5720 3269 5721
rect 3271 5720 3272 5721
rect 3520 5720 3521 5721
rect 3283 5722 3284 5723
rect 3307 5722 3308 5723
rect 3259 5724 3260 5725
rect 3307 5724 3308 5725
rect 3286 5726 3287 5727
rect 3523 5726 3524 5727
rect 3289 5728 3290 5729
rect 3334 5728 3335 5729
rect 3289 5730 3290 5731
rect 3502 5730 3503 5731
rect 3325 5732 3326 5733
rect 3364 5732 3365 5733
rect 3241 5734 3242 5735
rect 3325 5734 3326 5735
rect 2891 5736 2892 5737
rect 3241 5736 3242 5737
rect 3343 5736 3344 5737
rect 3586 5736 3587 5737
rect 2915 5738 2916 5739
rect 3343 5738 3344 5739
rect 3349 5738 3350 5739
rect 3352 5738 3353 5739
rect 3310 5740 3311 5741
rect 3349 5740 3350 5741
rect 3361 5740 3362 5741
rect 3890 5740 3891 5741
rect 3367 5742 3368 5743
rect 3604 5742 3605 5743
rect 3367 5744 3368 5745
rect 3388 5744 3389 5745
rect 3376 5746 3377 5747
rect 3469 5746 3470 5747
rect 3385 5748 3386 5749
rect 3613 5748 3614 5749
rect 3388 5750 3389 5751
rect 3625 5750 3626 5751
rect 3394 5752 3395 5753
rect 3574 5752 3575 5753
rect 3412 5754 3413 5755
rect 3957 5754 3958 5755
rect 3415 5756 3416 5757
rect 3448 5756 3449 5757
rect 3424 5758 3425 5759
rect 3674 5758 3675 5759
rect 3424 5760 3425 5761
rect 3790 5760 3791 5761
rect 3427 5762 3428 5763
rect 3574 5762 3575 5763
rect 3433 5764 3434 5765
rect 3616 5764 3617 5765
rect 3244 5766 3245 5767
rect 3433 5766 3434 5767
rect 3163 5768 3164 5769
rect 3244 5768 3245 5769
rect 3163 5770 3164 5771
rect 3187 5770 3188 5771
rect 3187 5772 3188 5773
rect 3397 5772 3398 5773
rect 3436 5772 3437 5773
rect 3496 5772 3497 5773
rect 3247 5774 3248 5775
rect 3496 5774 3497 5775
rect 3451 5776 3452 5777
rect 3640 5776 3641 5777
rect 3451 5778 3452 5779
rect 3658 5778 3659 5779
rect 3454 5780 3455 5781
rect 3825 5780 3826 5781
rect 3460 5782 3461 5783
rect 3649 5782 3650 5783
rect 3463 5784 3464 5785
rect 3664 5784 3665 5785
rect 3400 5786 3401 5787
rect 3463 5786 3464 5787
rect 2925 5788 2926 5789
rect 3400 5788 3401 5789
rect 3466 5788 3467 5789
rect 3514 5788 3515 5789
rect 3277 5790 3278 5791
rect 3514 5790 3515 5791
rect 3253 5792 3254 5793
rect 3277 5792 3278 5793
rect 3475 5792 3476 5793
rect 3658 5792 3659 5793
rect 3160 5794 3161 5795
rect 3475 5794 3476 5795
rect 3478 5794 3479 5795
rect 3911 5794 3912 5795
rect 3484 5796 3485 5797
rect 3908 5796 3909 5797
rect 3502 5798 3503 5799
rect 3556 5798 3557 5799
rect 3313 5800 3314 5801
rect 3556 5800 3557 5801
rect 3265 5802 3266 5803
rect 3313 5802 3314 5803
rect 3526 5802 3527 5803
rect 3893 5802 3894 5803
rect 3529 5804 3530 5805
rect 3580 5804 3581 5805
rect 3508 5806 3509 5807
rect 3580 5806 3581 5807
rect 3337 5808 3338 5809
rect 3508 5808 3509 5809
rect 3535 5808 3536 5809
rect 4013 5808 4014 5809
rect 3538 5810 3539 5811
rect 3864 5810 3865 5811
rect 3301 5812 3302 5813
rect 3538 5812 3539 5813
rect 3301 5814 3302 5815
rect 3850 5814 3851 5815
rect 3541 5816 3542 5817
rect 3670 5816 3671 5817
rect 3547 5818 3548 5819
rect 3610 5818 3611 5819
rect 3373 5820 3374 5821
rect 3610 5820 3611 5821
rect 3036 5822 3037 5823
rect 3373 5822 3374 5823
rect 3550 5822 3551 5823
rect 3589 5822 3590 5823
rect 3562 5824 3563 5825
rect 3568 5824 3569 5825
rect 3598 5824 3599 5825
rect 3730 5824 3731 5825
rect 3355 5826 3356 5827
rect 3598 5826 3599 5827
rect 3628 5826 3629 5827
rect 4030 5826 4031 5827
rect 3628 5828 3629 5829
rect 3695 5828 3696 5829
rect 3634 5830 3635 5831
rect 3745 5830 3746 5831
rect 3409 5832 3410 5833
rect 3634 5832 3635 5833
rect 3643 5832 3644 5833
rect 3748 5832 3749 5833
rect 3655 5834 3656 5835
rect 3743 5834 3744 5835
rect 3631 5836 3632 5837
rect 3742 5836 3743 5837
rect 3661 5838 3662 5839
rect 3766 5838 3767 5839
rect 3673 5840 3674 5841
rect 3960 5840 3961 5841
rect 3679 5842 3680 5843
rect 3874 5842 3875 5843
rect 3689 5844 3690 5845
rect 3799 5844 3800 5845
rect 3692 5846 3693 5847
rect 3823 5846 3824 5847
rect 3691 5848 3692 5849
rect 3871 5848 3872 5849
rect 3139 5850 3140 5851
rect 3871 5850 3872 5851
rect 3698 5852 3699 5853
rect 3820 5852 3821 5853
rect 3487 5854 3488 5855
rect 3697 5854 3698 5855
rect 3713 5854 3714 5855
rect 3862 5854 3863 5855
rect 3712 5856 3713 5857
rect 4010 5856 4011 5857
rect 3716 5858 3717 5859
rect 3811 5858 3812 5859
rect 3532 5860 3533 5861
rect 3715 5860 3716 5861
rect 3331 5862 3332 5863
rect 3532 5862 3533 5863
rect 3211 5864 3212 5865
rect 3331 5864 3332 5865
rect 3718 5864 3719 5865
rect 4017 5864 4018 5865
rect 3725 5866 3726 5867
rect 4003 5866 4004 5867
rect 3724 5868 3725 5869
rect 3814 5868 3815 5869
rect 3737 5870 3738 5871
rect 3865 5870 3866 5871
rect 3736 5872 3737 5873
rect 3935 5872 3936 5873
rect 3740 5874 3741 5875
rect 3868 5874 3869 5875
rect 3754 5876 3755 5877
rect 3828 5876 3829 5877
rect 3701 5878 3702 5879
rect 3829 5878 3830 5879
rect 3757 5880 3758 5881
rect 3884 5880 3885 5881
rect 3760 5882 3761 5883
rect 3808 5882 3809 5883
rect 3583 5884 3584 5885
rect 3760 5884 3761 5885
rect 3763 5884 3764 5885
rect 3860 5884 3861 5885
rect 3223 5886 3224 5887
rect 3859 5886 3860 5887
rect 3223 5888 3224 5889
rect 3319 5888 3320 5889
rect 3769 5888 3770 5889
rect 3914 5888 3915 5889
rect 3772 5890 3773 5891
rect 3996 5890 3997 5891
rect 3781 5892 3782 5893
rect 3926 5892 3927 5893
rect 3622 5894 3623 5895
rect 3781 5894 3782 5895
rect 3391 5896 3392 5897
rect 3622 5896 3623 5897
rect 3784 5896 3785 5897
rect 3929 5896 3930 5897
rect 3784 5898 3785 5899
rect 3887 5898 3888 5899
rect 3787 5900 3788 5901
rect 3947 5900 3948 5901
rect 3793 5902 3794 5903
rect 3938 5902 3939 5903
rect 3707 5904 3708 5905
rect 3793 5904 3794 5905
rect 3796 5904 3797 5905
rect 3941 5904 3942 5905
rect 3805 5906 3806 5907
rect 3944 5906 3945 5907
rect 3686 5908 3687 5909
rect 3805 5908 3806 5909
rect 3481 5910 3482 5911
rect 3685 5910 3686 5911
rect 3817 5910 3818 5911
rect 4020 5910 4021 5911
rect 3826 5912 3827 5913
rect 3932 5912 3933 5913
rect 3832 5914 3833 5915
rect 3841 5914 3842 5915
rect 3844 5914 3845 5915
rect 3983 5914 3984 5915
rect 3847 5916 3848 5917
rect 3986 5916 3987 5917
rect 3853 5918 3854 5919
rect 3902 5918 3903 5919
rect 3905 5918 3906 5919
rect 3989 5918 3990 5919
rect 2857 5927 2858 5928
rect 3150 5927 3151 5928
rect 2872 5929 2873 5930
rect 2879 5929 2880 5930
rect 2887 5929 2888 5930
rect 3053 5929 3054 5930
rect 2890 5931 2891 5932
rect 3277 5931 3278 5932
rect 2899 5933 2900 5934
rect 3241 5933 3242 5934
rect 2915 5935 2916 5936
rect 3117 5935 3118 5936
rect 2919 5937 2920 5938
rect 3295 5937 3296 5938
rect 2922 5939 2923 5940
rect 2926 5939 2927 5940
rect 2930 5939 2931 5940
rect 2990 5939 2991 5940
rect 2951 5941 2952 5942
rect 3207 5941 3208 5942
rect 2954 5943 2955 5944
rect 3331 5943 3332 5944
rect 2964 5945 2965 5946
rect 2984 5945 2985 5946
rect 2968 5947 2969 5948
rect 3279 5947 3280 5948
rect 2967 5949 2968 5950
rect 2990 5949 2991 5950
rect 2978 5951 2979 5952
rect 3499 5951 3500 5952
rect 2993 5953 2994 5954
rect 3313 5953 3314 5954
rect 2996 5955 2997 5956
rect 3127 5955 3128 5956
rect 3008 5957 3009 5958
rect 3256 5957 3257 5958
rect 3002 5959 3003 5960
rect 3008 5959 3009 5960
rect 3015 5959 3016 5960
rect 3334 5959 3335 5960
rect 3018 5961 3019 5962
rect 3264 5961 3265 5962
rect 3026 5963 3027 5964
rect 3094 5963 3095 5964
rect 3029 5965 3030 5966
rect 3070 5965 3071 5966
rect 3021 5967 3022 5968
rect 3071 5967 3072 5968
rect 3033 5969 3034 5970
rect 3163 5969 3164 5970
rect 3036 5971 3037 5972
rect 3126 5971 3127 5972
rect 3041 5973 3042 5974
rect 3082 5973 3083 5974
rect 3055 5975 3056 5976
rect 3223 5975 3224 5976
rect 3068 5977 3069 5978
rect 3273 5977 3274 5978
rect 3076 5979 3077 5980
rect 3202 5979 3203 5980
rect 3079 5981 3080 5982
rect 3385 5981 3386 5982
rect 2952 5983 2953 5984
rect 3080 5983 3081 5984
rect 3083 5983 3084 5984
rect 3139 5983 3140 5984
rect 3086 5985 3087 5986
rect 3133 5985 3134 5986
rect 2916 5987 2917 5988
rect 3132 5987 3133 5988
rect 3093 5989 3094 5990
rect 3349 5989 3350 5990
rect 3096 5991 3097 5992
rect 3145 5991 3146 5992
rect 3099 5993 3100 5994
rect 3148 5993 3149 5994
rect 3103 5995 3104 5996
rect 3540 5995 3541 5996
rect 2961 5997 2962 5998
rect 3102 5997 3103 5998
rect 3108 5997 3109 5998
rect 3298 5997 3299 5998
rect 3114 5999 3115 6000
rect 3181 5999 3182 6000
rect 3138 6001 3139 6002
rect 3343 6001 3344 6002
rect 3144 6003 3145 6004
rect 3433 6003 3434 6004
rect 3157 6005 3158 6006
rect 3787 6005 3788 6006
rect 3159 6007 3160 6008
rect 3268 6007 3269 6008
rect 3162 6009 3163 6010
rect 3229 6009 3230 6010
rect 3168 6011 3169 6012
rect 3217 6011 3218 6012
rect 3174 6013 3175 6014
rect 3193 6013 3194 6014
rect 3180 6015 3181 6016
rect 3244 6015 3245 6016
rect 3187 6017 3188 6018
rect 3935 6017 3936 6018
rect 2945 6019 2946 6020
rect 3186 6019 3187 6020
rect 3192 6019 3193 6020
rect 3463 6019 3464 6020
rect 3205 6021 3206 6022
rect 3642 6021 3643 6022
rect 3204 6023 3205 6024
rect 3340 6023 3341 6024
rect 3045 6025 3046 6026
rect 3339 6025 3340 6026
rect 3210 6027 3211 6028
rect 3262 6027 3263 6028
rect 3216 6029 3217 6030
rect 3370 6029 3371 6030
rect 3219 6031 3220 6032
rect 3373 6031 3374 6032
rect 3222 6033 3223 6034
rect 3283 6033 3284 6034
rect 3121 6035 3122 6036
rect 3282 6035 3283 6036
rect 2999 6037 3000 6038
rect 3120 6037 3121 6038
rect 3228 6037 3229 6038
rect 3358 6037 3359 6038
rect 3235 6039 3236 6040
rect 3348 6039 3349 6040
rect 3234 6041 3235 6042
rect 3325 6041 3326 6042
rect 3240 6043 3241 6044
rect 3307 6043 3308 6044
rect 3017 6045 3018 6046
rect 3306 6045 3307 6046
rect 3246 6047 3247 6048
rect 3400 6047 3401 6048
rect 3249 6049 3250 6050
rect 3403 6049 3404 6050
rect 3252 6051 3253 6052
rect 3406 6051 3407 6052
rect 3258 6053 3259 6054
rect 3418 6053 3419 6054
rect 3261 6055 3262 6056
rect 3421 6055 3422 6056
rect 3270 6057 3271 6058
rect 3346 6057 3347 6058
rect 3090 6059 3091 6060
rect 3345 6059 3346 6060
rect 3276 6061 3277 6062
rect 3430 6061 3431 6062
rect 3289 6063 3290 6064
rect 3480 6063 3481 6064
rect 3294 6065 3295 6066
rect 3472 6065 3473 6066
rect 3297 6067 3298 6068
rect 3475 6067 3476 6068
rect 3309 6069 3310 6070
rect 3316 6069 3317 6070
rect 3312 6071 3313 6072
rect 3496 6071 3497 6072
rect 3315 6073 3316 6074
rect 3442 6073 3443 6074
rect 3318 6075 3319 6076
rect 3364 6075 3365 6076
rect 3330 6077 3331 6078
rect 3514 6077 3515 6078
rect 3336 6079 3337 6080
rect 3520 6079 3521 6080
rect 3342 6081 3343 6082
rect 3460 6081 3461 6082
rect 3354 6083 3355 6084
rect 3702 6083 3703 6084
rect 3360 6085 3361 6086
rect 3544 6085 3545 6086
rect 3372 6087 3373 6088
rect 3556 6087 3557 6088
rect 3384 6089 3385 6090
rect 3508 6089 3509 6090
rect 3388 6091 3389 6092
rect 3699 6091 3700 6092
rect 3390 6093 3391 6094
rect 3526 6093 3527 6094
rect 3376 6095 3377 6096
rect 3525 6095 3526 6096
rect 3402 6097 3403 6098
rect 3630 6097 3631 6098
rect 3408 6099 3409 6100
rect 3610 6099 3611 6100
rect 3412 6101 3413 6102
rect 3606 6101 3607 6102
rect 3414 6103 3415 6104
rect 3598 6103 3599 6104
rect 3420 6105 3421 6106
rect 3604 6105 3605 6106
rect 3432 6107 3433 6108
rect 3484 6107 3485 6108
rect 3438 6109 3439 6110
rect 3622 6109 3623 6110
rect 3444 6111 3445 6112
rect 3932 6111 3933 6112
rect 3448 6113 3449 6114
rect 3636 6113 3637 6114
rect 3456 6115 3457 6116
rect 3634 6115 3635 6116
rect 3451 6117 3452 6118
rect 3633 6117 3634 6118
rect 3450 6119 3451 6120
rect 3616 6119 3617 6120
rect 3462 6121 3463 6122
rect 3574 6121 3575 6122
rect 3474 6123 3475 6124
rect 3960 6123 3961 6124
rect 3478 6125 3479 6126
rect 3957 6125 3958 6126
rect 3486 6127 3487 6128
rect 3658 6127 3659 6128
rect 3454 6129 3455 6130
rect 3657 6129 3658 6130
rect 3492 6131 3493 6132
rect 3670 6131 3671 6132
rect 3495 6133 3496 6134
rect 3664 6133 3665 6134
rect 3513 6135 3514 6136
rect 3685 6135 3686 6136
rect 3519 6137 3520 6138
rect 3691 6137 3692 6138
rect 3523 6139 3524 6140
rect 3705 6139 3706 6140
rect 3529 6141 3530 6142
rect 3603 6141 3604 6142
rect 3538 6143 3539 6144
rect 3760 6143 3761 6144
rect 3199 6145 3200 6146
rect 3537 6145 3538 6146
rect 3543 6145 3544 6146
rect 3652 6145 3653 6146
rect 3549 6147 3550 6148
rect 3580 6147 3581 6148
rect 3466 6149 3467 6150
rect 3579 6149 3580 6150
rect 3553 6151 3554 6152
rect 3576 6151 3577 6152
rect 3555 6153 3556 6154
rect 3712 6153 3713 6154
rect 3532 6155 3533 6156
rect 3712 6155 3713 6156
rect 3301 6157 3302 6158
rect 3531 6157 3532 6158
rect 3558 6157 3559 6158
rect 3679 6157 3680 6158
rect 3561 6159 3562 6160
rect 3673 6159 3674 6160
rect 3367 6161 3368 6162
rect 3672 6161 3673 6162
rect 3366 6163 3367 6164
rect 3424 6163 3425 6164
rect 3568 6163 3569 6164
rect 3591 6163 3592 6164
rect 3394 6165 3395 6166
rect 3567 6165 3568 6166
rect 3573 6165 3574 6166
rect 3589 6165 3590 6166
rect 3615 6165 3616 6166
rect 3724 6165 3725 6166
rect 3621 6167 3622 6168
rect 3730 6167 3731 6168
rect 3628 6169 3629 6170
rect 3874 6169 3875 6170
rect 3396 6171 3397 6172
rect 3627 6171 3628 6172
rect 3640 6171 3641 6172
rect 3893 6171 3894 6172
rect 3547 6173 3548 6174
rect 3639 6173 3640 6174
rect 3651 6173 3652 6174
rect 3748 6173 3749 6174
rect 3663 6175 3664 6176
rect 3999 6175 4000 6176
rect 3687 6177 3688 6178
rect 3754 6177 3755 6178
rect 3693 6179 3694 6180
rect 3742 6179 3743 6180
rect 3697 6181 3698 6182
rect 4037 6181 4038 6182
rect 3696 6183 3697 6184
rect 3778 6183 3779 6184
rect 3715 6185 3716 6186
rect 4013 6185 4014 6186
rect 3718 6187 3719 6188
rect 4027 6187 4028 6188
rect 3727 6189 3728 6190
rect 3805 6189 3806 6190
rect 3730 6191 3731 6192
rect 3799 6191 3800 6192
rect 3733 6193 3734 6194
rect 3817 6193 3818 6194
rect 3736 6195 3737 6196
rect 3950 6195 3951 6196
rect 3736 6197 3737 6198
rect 3823 6197 3824 6198
rect 3739 6199 3740 6200
rect 3826 6199 3827 6200
rect 3745 6201 3746 6202
rect 3890 6201 3891 6202
rect 3748 6203 3749 6204
rect 3823 6203 3824 6204
rect 3760 6205 3761 6206
rect 3859 6205 3860 6206
rect 3763 6207 3764 6208
rect 3862 6207 3863 6208
rect 3766 6209 3767 6210
rect 3996 6209 3997 6210
rect 3766 6211 3767 6212
rect 3868 6211 3869 6212
rect 3769 6213 3770 6214
rect 3793 6213 3794 6214
rect 3586 6215 3587 6216
rect 3793 6215 3794 6216
rect 3502 6217 3503 6218
rect 3585 6217 3586 6218
rect 3048 6219 3049 6220
rect 3501 6219 3502 6220
rect 3772 6219 3773 6220
rect 3814 6219 3815 6220
rect 3436 6221 3437 6222
rect 3772 6221 3773 6222
rect 3779 6221 3780 6222
rect 3790 6221 3791 6222
rect 3784 6223 3785 6224
rect 4040 6223 4041 6224
rect 3786 6225 3787 6226
rect 3865 6225 3866 6226
rect 3796 6227 3797 6228
rect 3844 6227 3845 6228
rect 3805 6229 3806 6230
rect 3938 6229 3939 6230
rect 3808 6231 3809 6232
rect 3941 6231 3942 6232
rect 3811 6233 3812 6234
rect 3926 6233 3927 6234
rect 3817 6235 3818 6236
rect 3944 6235 3945 6236
rect 3826 6237 3827 6238
rect 3841 6237 3842 6238
rect 3781 6239 3782 6240
rect 3840 6239 3841 6240
rect 3829 6241 3830 6242
rect 3853 6241 3854 6242
rect 3789 6243 3790 6244
rect 3830 6243 3831 6244
rect 3847 6243 3848 6244
rect 3905 6243 3906 6244
rect 3850 6245 3851 6246
rect 3986 6245 3987 6246
rect 3859 6247 3860 6248
rect 3884 6247 3885 6248
rect 3820 6249 3821 6250
rect 3884 6249 3885 6250
rect 3820 6251 3821 6252
rect 3947 6251 3948 6252
rect 3866 6253 3867 6254
rect 3914 6253 3915 6254
rect 3902 6255 3903 6256
rect 3992 6255 3993 6256
rect 3929 6257 3930 6258
rect 4003 6257 4004 6258
rect 3953 6259 3954 6260
rect 3983 6259 3984 6260
rect 2872 6268 2873 6269
rect 3150 6268 3151 6269
rect 2875 6270 2876 6271
rect 3064 6270 3065 6271
rect 2879 6272 2880 6273
rect 2913 6272 2914 6273
rect 2878 6274 2879 6275
rect 3053 6274 3054 6275
rect 2897 6276 2898 6277
rect 3159 6276 3160 6277
rect 2902 6278 2903 6279
rect 3096 6278 3097 6279
rect 2903 6280 2904 6281
rect 3080 6280 3081 6281
rect 2906 6282 2907 6283
rect 3219 6282 3220 6283
rect 2909 6284 2910 6285
rect 3699 6284 3700 6285
rect 2910 6286 2911 6287
rect 3190 6286 3191 6287
rect 2914 6288 2915 6289
rect 3246 6288 3247 6289
rect 2927 6290 2928 6291
rect 3132 6290 3133 6291
rect 2930 6292 2931 6293
rect 3138 6292 3139 6293
rect 2933 6294 2934 6295
rect 2939 6294 2940 6295
rect 2945 6294 2946 6295
rect 3220 6294 3221 6295
rect 2948 6296 2949 6297
rect 3162 6296 3163 6297
rect 2948 6298 2949 6299
rect 3154 6298 3155 6299
rect 2964 6300 2965 6301
rect 3258 6300 3259 6301
rect 2967 6302 2968 6303
rect 3099 6302 3100 6303
rect 2967 6304 2968 6305
rect 3238 6304 3239 6305
rect 2971 6306 2972 6307
rect 3014 6306 3015 6307
rect 2971 6308 2972 6309
rect 3256 6308 3257 6309
rect 2978 6310 2979 6311
rect 3106 6310 3107 6311
rect 2955 6312 2956 6313
rect 2978 6312 2979 6313
rect 2955 6314 2956 6315
rect 2981 6314 2982 6315
rect 2999 6314 3000 6315
rect 3102 6314 3103 6315
rect 3016 6316 3017 6317
rect 3304 6316 3305 6317
rect 3026 6318 3027 6319
rect 3031 6318 3032 6319
rect 3029 6320 3030 6321
rect 3058 6320 3059 6321
rect 3046 6322 3047 6323
rect 3117 6322 3118 6323
rect 3061 6324 3062 6325
rect 3249 6324 3250 6325
rect 3086 6326 3087 6327
rect 3136 6326 3137 6327
rect 3067 6328 3068 6329
rect 3085 6328 3086 6329
rect 3090 6328 3091 6329
rect 3318 6328 3319 6329
rect 2952 6330 2953 6331
rect 3091 6330 3092 6331
rect 2907 6332 2908 6333
rect 2952 6332 2953 6333
rect 3093 6332 3094 6333
rect 3351 6332 3352 6333
rect 3100 6334 3101 6335
rect 3192 6334 3193 6335
rect 3103 6336 3104 6337
rect 3345 6336 3346 6337
rect 3108 6338 3109 6339
rect 3112 6338 3113 6339
rect 3114 6338 3115 6339
rect 3118 6338 3119 6339
rect 3126 6338 3127 6339
rect 3342 6338 3343 6339
rect 3070 6340 3071 6341
rect 3343 6340 3344 6341
rect 3129 6342 3130 6343
rect 3396 6342 3397 6343
rect 3120 6344 3121 6345
rect 3130 6344 3131 6345
rect 2923 6346 2924 6347
rect 3121 6346 3122 6347
rect 3142 6346 3143 6347
rect 3144 6346 3145 6347
rect 3148 6346 3149 6347
rect 3168 6346 3169 6347
rect 3166 6348 3167 6349
rect 3180 6348 3181 6349
rect 3172 6350 3173 6351
rect 3174 6350 3175 6351
rect 3178 6350 3179 6351
rect 3282 6350 3283 6351
rect 3184 6352 3185 6353
rect 3186 6352 3187 6353
rect 3196 6352 3197 6353
rect 3204 6352 3205 6353
rect 3199 6354 3200 6355
rect 3207 6354 3208 6355
rect 3202 6356 3203 6357
rect 3210 6356 3211 6357
rect 3041 6358 3042 6359
rect 3211 6358 3212 6359
rect 3208 6360 3209 6361
rect 3216 6360 3217 6361
rect 3214 6362 3215 6363
rect 3228 6362 3229 6363
rect 3222 6364 3223 6365
rect 3232 6364 3233 6365
rect 3226 6366 3227 6367
rect 3537 6366 3538 6367
rect 3234 6368 3235 6369
rect 3244 6368 3245 6369
rect 3250 6368 3251 6369
rect 3252 6368 3253 6369
rect 3264 6368 3265 6369
rect 3286 6368 3287 6369
rect 3268 6370 3269 6371
rect 3315 6370 3316 6371
rect 3270 6372 3271 6373
rect 3316 6372 3317 6373
rect 3273 6374 3274 6375
rect 3319 6374 3320 6375
rect 3274 6376 3275 6377
rect 3276 6376 3277 6377
rect 3277 6378 3278 6379
rect 3279 6378 3280 6379
rect 3292 6378 3293 6379
rect 3294 6378 3295 6379
rect 3295 6380 3296 6381
rect 3297 6380 3298 6381
rect 3298 6382 3299 6383
rect 3306 6382 3307 6383
rect 3307 6384 3308 6385
rect 3309 6384 3310 6385
rect 3310 6386 3311 6387
rect 3312 6386 3313 6387
rect 2981 6388 2982 6389
rect 3313 6388 3314 6389
rect 3328 6388 3329 6389
rect 3330 6388 3331 6389
rect 3334 6388 3335 6389
rect 3336 6388 3337 6389
rect 3337 6390 3338 6391
rect 3339 6390 3340 6391
rect 3340 6392 3341 6393
rect 3348 6392 3349 6393
rect 3346 6394 3347 6395
rect 3402 6394 3403 6395
rect 3349 6396 3350 6397
rect 3540 6396 3541 6397
rect 3352 6398 3353 6399
rect 3674 6398 3675 6399
rect 3354 6400 3355 6401
rect 3394 6400 3395 6401
rect 3358 6402 3359 6403
rect 3360 6402 3361 6403
rect 3364 6402 3365 6403
rect 3480 6402 3481 6403
rect 3366 6404 3367 6405
rect 3388 6404 3389 6405
rect 3367 6406 3368 6407
rect 3642 6406 3643 6407
rect 3370 6408 3371 6409
rect 3372 6408 3373 6409
rect 3376 6408 3377 6409
rect 3384 6408 3385 6409
rect 3382 6410 3383 6411
rect 3390 6410 3391 6411
rect 3400 6410 3401 6411
rect 3712 6410 3713 6411
rect 3406 6412 3407 6413
rect 3752 6412 3753 6413
rect 3408 6414 3409 6415
rect 3778 6414 3779 6415
rect 3412 6416 3413 6417
rect 3414 6416 3415 6417
rect 3418 6416 3419 6417
rect 3420 6416 3421 6417
rect 3424 6416 3425 6417
rect 3772 6416 3773 6417
rect 3430 6418 3431 6419
rect 3432 6418 3433 6419
rect 3436 6418 3437 6419
rect 3462 6418 3463 6419
rect 3442 6420 3443 6421
rect 3456 6420 3457 6421
rect 3444 6422 3445 6423
rect 3448 6422 3449 6423
rect 3454 6422 3455 6423
rect 3525 6422 3526 6423
rect 3466 6424 3467 6425
rect 3782 6424 3783 6425
rect 3472 6426 3473 6427
rect 3495 6426 3496 6427
rect 3474 6428 3475 6429
rect 3830 6428 3831 6429
rect 3478 6430 3479 6431
rect 3492 6430 3493 6431
rect 3493 6432 3494 6433
rect 3513 6432 3514 6433
rect 3501 6434 3502 6435
rect 3627 6434 3628 6435
rect 3505 6436 3506 6437
rect 3579 6436 3580 6437
rect 3511 6438 3512 6439
rect 3591 6438 3592 6439
rect 3517 6440 3518 6441
rect 3543 6440 3544 6441
rect 3519 6442 3520 6443
rect 3526 6442 3527 6443
rect 3523 6444 3524 6445
rect 3555 6444 3556 6445
rect 3529 6446 3530 6447
rect 3585 6446 3586 6447
rect 3531 6448 3532 6449
rect 3583 6448 3584 6449
rect 3535 6450 3536 6451
rect 3549 6450 3550 6451
rect 3553 6450 3554 6451
rect 3802 6450 3803 6451
rect 3556 6452 3557 6453
rect 3576 6452 3577 6453
rect 3558 6454 3559 6455
rect 3880 6454 3881 6455
rect 3561 6456 3562 6457
rect 3845 6456 3846 6457
rect 3565 6458 3566 6459
rect 3615 6458 3616 6459
rect 3567 6460 3568 6461
rect 3571 6460 3572 6461
rect 3589 6460 3590 6461
rect 3603 6460 3604 6461
rect 3592 6462 3593 6463
rect 3608 6462 3609 6463
rect 3595 6464 3596 6465
rect 3633 6464 3634 6465
rect 3598 6466 3599 6467
rect 3639 6466 3640 6467
rect 3606 6468 3607 6469
rect 3702 6468 3703 6469
rect 3611 6470 3612 6471
rect 3657 6470 3658 6471
rect 3617 6472 3618 6473
rect 3840 6472 3841 6473
rect 3630 6474 3631 6475
rect 3793 6474 3794 6475
rect 3621 6476 3622 6477
rect 3793 6476 3794 6477
rect 3636 6478 3637 6479
rect 3755 6478 3756 6479
rect 3635 6480 3636 6481
rect 3651 6480 3652 6481
rect 3641 6482 3642 6483
rect 3663 6482 3664 6483
rect 3647 6484 3648 6485
rect 3687 6484 3688 6485
rect 3653 6486 3654 6487
rect 3814 6486 3815 6487
rect 3659 6488 3660 6489
rect 3696 6488 3697 6489
rect 3662 6490 3663 6491
rect 3665 6490 3666 6491
rect 3669 6490 3670 6491
rect 3705 6490 3706 6491
rect 3000 6492 3001 6493
rect 3668 6492 3669 6493
rect 3672 6492 3673 6493
rect 3775 6492 3776 6493
rect 3677 6494 3678 6495
rect 3693 6494 3694 6495
rect 3698 6494 3699 6495
rect 3727 6494 3728 6495
rect 3701 6496 3702 6497
rect 3823 6496 3824 6497
rect 3704 6498 3705 6499
rect 3736 6498 3737 6499
rect 3707 6500 3708 6501
rect 3739 6500 3740 6501
rect 3716 6502 3717 6503
rect 3760 6502 3761 6503
rect 3541 6504 3542 6505
rect 3759 6504 3760 6505
rect 3719 6506 3720 6507
rect 3748 6506 3749 6507
rect 3728 6508 3729 6509
rect 3769 6508 3770 6509
rect 3573 6510 3574 6511
rect 3769 6510 3770 6511
rect 3733 6512 3734 6513
rect 3887 6512 3888 6513
rect 3734 6514 3735 6515
rect 3766 6514 3767 6515
rect 3746 6516 3747 6517
rect 3789 6516 3790 6517
rect 3749 6518 3750 6519
rect 3786 6518 3787 6519
rect 3763 6520 3764 6521
rect 3826 6520 3827 6521
rect 3559 6522 3560 6523
rect 3762 6522 3763 6523
rect 3730 6524 3731 6525
rect 3826 6524 3827 6525
rect 3772 6526 3773 6527
rect 3811 6526 3812 6527
rect 3790 6528 3791 6529
rect 3805 6528 3806 6529
rect 3450 6530 3451 6531
rect 3805 6530 3806 6531
rect 3796 6532 3797 6533
rect 3837 6532 3838 6533
rect 3796 6534 3797 6535
rect 3817 6534 3818 6535
rect 3799 6536 3800 6537
rect 3820 6536 3821 6537
rect 3671 6538 3672 6539
rect 3819 6538 3820 6539
rect 3808 6540 3809 6541
rect 3842 6540 3843 6541
rect 3438 6542 3439 6543
rect 3809 6542 3810 6543
rect 3829 6542 3830 6543
rect 3850 6542 3851 6543
rect 3832 6544 3833 6545
rect 3853 6544 3854 6545
rect 3847 6546 3848 6547
rect 3866 6546 3867 6547
rect 3859 6548 3860 6549
rect 3870 6548 3871 6549
rect 3008 6550 3009 6551
rect 3869 6550 3870 6551
rect 3863 6552 3864 6553
rect 3873 6552 3874 6553
rect 2887 6561 2888 6562
rect 2896 6561 2897 6562
rect 2890 6563 2891 6564
rect 3064 6563 3065 6564
rect 2900 6565 2901 6566
rect 3268 6565 3269 6566
rect 2903 6567 2904 6568
rect 3144 6567 3145 6568
rect 2907 6569 2908 6570
rect 2921 6569 2922 6570
rect 2907 6571 2908 6572
rect 3154 6571 3155 6572
rect 2924 6573 2925 6574
rect 3202 6573 3203 6574
rect 2924 6575 2925 6576
rect 3046 6575 3047 6576
rect 2928 6577 2929 6578
rect 3045 6577 3046 6578
rect 2933 6579 2934 6580
rect 2940 6579 2941 6580
rect 2945 6579 2946 6580
rect 3214 6579 3215 6580
rect 2952 6581 2953 6582
rect 3081 6581 3082 6582
rect 2962 6583 2963 6584
rect 2991 6583 2992 6584
rect 2964 6585 2965 6586
rect 3258 6585 3259 6586
rect 2974 6587 2975 6588
rect 3250 6587 3251 6588
rect 2974 6589 2975 6590
rect 3246 6589 3247 6590
rect 2981 6591 2982 6592
rect 3241 6591 3242 6592
rect 2985 6593 2986 6594
rect 3190 6593 3191 6594
rect 2995 6595 2996 6596
rect 3292 6595 3293 6596
rect 3004 6597 3005 6598
rect 3031 6597 3032 6598
rect 3006 6599 3007 6600
rect 3106 6599 3107 6600
rect 2917 6601 2918 6602
rect 3105 6601 3106 6602
rect 3000 6603 3001 6604
rect 3007 6603 3008 6604
rect 3013 6603 3014 6604
rect 3605 6603 3606 6604
rect 3016 6605 3017 6606
rect 3252 6605 3253 6606
rect 3030 6607 3031 6608
rect 3334 6607 3335 6608
rect 3034 6609 3035 6610
rect 3337 6609 3338 6610
rect 3033 6611 3034 6612
rect 3058 6611 3059 6612
rect 3037 6613 3038 6614
rect 3321 6613 3322 6614
rect 3036 6615 3037 6616
rect 3061 6615 3062 6616
rect 3063 6615 3064 6616
rect 3330 6615 3331 6616
rect 3070 6617 3071 6618
rect 3333 6617 3334 6618
rect 3085 6619 3086 6620
rect 3349 6619 3350 6620
rect 3084 6621 3085 6622
rect 3091 6621 3092 6622
rect 3100 6621 3101 6622
rect 3189 6621 3190 6622
rect 3099 6623 3100 6624
rect 3112 6623 3113 6624
rect 3108 6625 3109 6626
rect 3118 6625 3119 6626
rect 3111 6627 3112 6628
rect 3121 6627 3122 6628
rect 3126 6627 3127 6628
rect 3130 6627 3131 6628
rect 3132 6627 3133 6628
rect 3142 6627 3143 6628
rect 3136 6629 3137 6630
rect 3234 6629 3235 6630
rect 3138 6631 3139 6632
rect 3148 6631 3149 6632
rect 3150 6631 3151 6632
rect 3166 6631 3167 6632
rect 3156 6633 3157 6634
rect 3343 6633 3344 6634
rect 3162 6635 3163 6636
rect 3172 6635 3173 6636
rect 3165 6637 3166 6638
rect 3295 6637 3296 6638
rect 3020 6639 3021 6640
rect 3294 6639 3295 6640
rect 3174 6641 3175 6642
rect 3184 6641 3185 6642
rect 3178 6643 3179 6644
rect 3438 6643 3439 6644
rect 3180 6645 3181 6646
rect 3196 6645 3197 6646
rect 3183 6647 3184 6648
rect 3199 6647 3200 6648
rect 3192 6649 3193 6650
rect 3208 6649 3209 6650
rect 3195 6651 3196 6652
rect 3211 6651 3212 6652
rect 3204 6653 3205 6654
rect 3220 6653 3221 6654
rect 3210 6655 3211 6656
rect 3232 6655 3233 6656
rect 3216 6657 3217 6658
rect 3244 6657 3245 6658
rect 3222 6659 3223 6660
rect 3238 6659 3239 6660
rect 3226 6661 3227 6662
rect 3355 6661 3356 6662
rect 2952 6663 2953 6664
rect 3225 6663 3226 6664
rect 3228 6663 3229 6664
rect 3262 6663 3263 6664
rect 3240 6665 3241 6666
rect 3256 6665 3257 6666
rect 3264 6665 3265 6666
rect 3274 6665 3275 6666
rect 3267 6667 3268 6668
rect 3277 6667 3278 6668
rect 3270 6669 3271 6670
rect 3286 6669 3287 6670
rect 3276 6671 3277 6672
rect 3316 6671 3317 6672
rect 3282 6673 3283 6674
rect 3298 6673 3299 6674
rect 3288 6675 3289 6676
rect 3304 6675 3305 6676
rect 3291 6677 3292 6678
rect 3307 6677 3308 6678
rect 3300 6679 3301 6680
rect 3310 6679 3311 6680
rect 3303 6681 3304 6682
rect 3313 6681 3314 6682
rect 3088 6683 3089 6684
rect 3312 6683 3313 6684
rect 2971 6685 2972 6686
rect 3087 6685 3088 6686
rect 2971 6687 2972 6688
rect 3261 6687 3262 6688
rect 3315 6687 3316 6688
rect 3319 6687 3320 6688
rect 3318 6689 3319 6690
rect 3328 6689 3329 6690
rect 3324 6691 3325 6692
rect 3340 6691 3341 6692
rect 3339 6693 3340 6694
rect 3352 6693 3353 6694
rect 3348 6695 3349 6696
rect 3358 6695 3359 6696
rect 3364 6695 3365 6696
rect 3390 6695 3391 6696
rect 3367 6697 3368 6698
rect 3597 6697 3598 6698
rect 3366 6699 3367 6700
rect 3370 6699 3371 6700
rect 3372 6699 3373 6700
rect 3863 6699 3864 6700
rect 3376 6701 3377 6702
rect 3378 6701 3379 6702
rect 3382 6701 3383 6702
rect 3384 6701 3385 6702
rect 3388 6701 3389 6702
rect 3396 6701 3397 6702
rect 3394 6703 3395 6704
rect 3420 6703 3421 6704
rect 3402 6705 3403 6706
rect 3412 6705 3413 6706
rect 3406 6707 3407 6708
rect 3426 6707 3427 6708
rect 3418 6709 3419 6710
rect 3585 6709 3586 6710
rect 3430 6711 3431 6712
rect 3456 6711 3457 6712
rect 3432 6713 3433 6714
rect 3744 6713 3745 6714
rect 3436 6715 3437 6716
rect 3450 6715 3451 6716
rect 3448 6717 3449 6718
rect 3462 6717 3463 6718
rect 3468 6717 3469 6718
rect 3807 6717 3808 6718
rect 3472 6719 3473 6720
rect 3489 6719 3490 6720
rect 3478 6721 3479 6722
rect 3480 6721 3481 6722
rect 3487 6721 3488 6722
rect 3501 6721 3502 6722
rect 3493 6723 3494 6724
rect 3507 6723 3508 6724
rect 3511 6723 3512 6724
rect 3810 6723 3811 6724
rect 3523 6725 3524 6726
rect 3816 6725 3817 6726
rect 3517 6727 3518 6728
rect 3522 6727 3523 6728
rect 3526 6727 3527 6728
rect 3852 6727 3853 6728
rect 3535 6729 3536 6730
rect 3546 6729 3547 6730
rect 3529 6731 3530 6732
rect 3534 6731 3535 6732
rect 3505 6733 3506 6734
rect 3528 6733 3529 6734
rect 3571 6733 3572 6734
rect 3759 6733 3760 6734
rect 3565 6735 3566 6736
rect 3570 6735 3571 6736
rect 3559 6737 3560 6738
rect 3564 6737 3565 6738
rect 3576 6737 3577 6738
rect 3583 6737 3584 6738
rect 3582 6739 3583 6740
rect 3793 6739 3794 6740
rect 3589 6741 3590 6742
rect 3608 6741 3609 6742
rect 3342 6743 3343 6744
rect 3609 6743 3610 6744
rect 3588 6745 3589 6746
rect 3592 6745 3593 6746
rect 3400 6747 3401 6748
rect 3591 6747 3592 6748
rect 3603 6747 3604 6748
rect 3617 6747 3618 6748
rect 3611 6749 3612 6750
rect 3621 6749 3622 6750
rect 3360 6751 3361 6752
rect 3612 6751 3613 6752
rect 3627 6751 3628 6752
rect 3659 6751 3660 6752
rect 3630 6753 3631 6754
rect 3668 6753 3669 6754
rect 3466 6755 3467 6756
rect 3669 6755 3670 6756
rect 3633 6757 3634 6758
rect 3641 6757 3642 6758
rect 3635 6759 3636 6760
rect 3639 6759 3640 6760
rect 3645 6759 3646 6760
rect 3653 6759 3654 6760
rect 3474 6761 3475 6762
rect 3654 6761 3655 6762
rect 3651 6763 3652 6764
rect 3768 6763 3769 6764
rect 3662 6765 3663 6766
rect 3840 6765 3841 6766
rect 3663 6767 3664 6768
rect 3671 6767 3672 6768
rect 3424 6769 3425 6770
rect 3672 6769 3673 6770
rect 3666 6771 3667 6772
rect 3674 6771 3675 6772
rect 3454 6773 3455 6774
rect 3675 6773 3676 6774
rect 3677 6773 3678 6774
rect 3777 6773 3778 6774
rect 3678 6775 3679 6776
rect 3775 6775 3776 6776
rect 3690 6777 3691 6778
rect 3716 6777 3717 6778
rect 3693 6779 3694 6780
rect 3719 6779 3720 6780
rect 3696 6781 3697 6782
rect 3701 6781 3702 6782
rect 3698 6783 3699 6784
rect 3826 6783 3827 6784
rect 3442 6785 3443 6786
rect 3699 6785 3700 6786
rect 3346 6787 3347 6788
rect 3441 6787 3442 6788
rect 3103 6789 3104 6790
rect 3345 6789 3346 6790
rect 3702 6789 3703 6790
rect 3704 6789 3705 6790
rect 3705 6791 3706 6792
rect 3707 6791 3708 6792
rect 3714 6791 3715 6792
rect 3784 6791 3785 6792
rect 3720 6793 3721 6794
rect 3728 6793 3729 6794
rect 3726 6795 3727 6796
rect 3734 6795 3735 6796
rect 3732 6797 3733 6798
rect 3749 6797 3750 6798
rect 3746 6799 3747 6800
rect 3753 6799 3754 6800
rect 3750 6801 3751 6802
rect 3805 6801 3806 6802
rect 3756 6803 3757 6804
rect 3772 6803 3773 6804
rect 3771 6805 3772 6806
rect 3819 6805 3820 6806
rect 3794 6807 3795 6808
rect 3796 6807 3797 6808
rect 3647 6809 3648 6810
rect 3797 6809 3798 6810
rect 3799 6809 3800 6810
rect 3845 6809 3846 6810
rect 3827 6811 3828 6812
rect 3829 6811 3830 6812
rect 3830 6813 3831 6814
rect 3835 6813 3836 6814
rect 3832 6815 3833 6816
rect 3838 6815 3839 6816
rect 3849 6815 3850 6816
rect 3864 6815 3865 6816
rect 3790 6817 3791 6818
rect 3850 6817 3851 6818
rect 3408 6819 3409 6820
rect 3791 6819 3792 6820
rect 2896 6828 2897 6829
rect 3105 6828 3106 6829
rect 2907 6830 2908 6831
rect 3144 6830 3145 6831
rect 2912 6832 2913 6833
rect 3180 6832 3181 6833
rect 2914 6834 2915 6835
rect 3242 6834 3243 6835
rect 2922 6836 2923 6837
rect 3264 6836 3265 6837
rect 2924 6838 2925 6839
rect 3045 6838 3046 6839
rect 2940 6840 2941 6841
rect 2971 6840 2972 6841
rect 2952 6842 2953 6843
rect 3113 6842 3114 6843
rect 2959 6844 2960 6845
rect 2966 6844 2967 6845
rect 2963 6846 2964 6847
rect 3183 6846 3184 6847
rect 2978 6848 2979 6849
rect 3258 6848 3259 6849
rect 2979 6850 2980 6851
rect 3138 6850 3139 6851
rect 2981 6852 2982 6853
rect 3027 6852 3028 6853
rect 2982 6854 2983 6855
rect 3004 6854 3005 6855
rect 2917 6856 2918 6857
rect 3004 6856 3005 6857
rect 2985 6858 2986 6859
rect 3252 6858 3253 6859
rect 2988 6860 2989 6861
rect 3013 6860 3014 6861
rect 2995 6862 2996 6863
rect 3284 6862 3285 6863
rect 3007 6864 3008 6865
rect 3010 6864 3011 6865
rect 3022 6864 3023 6865
rect 3033 6864 3034 6865
rect 3034 6866 3035 6867
rect 3315 6866 3316 6867
rect 3036 6868 3037 6869
rect 3251 6868 3252 6869
rect 3037 6870 3038 6871
rect 3254 6870 3255 6871
rect 3044 6872 3045 6873
rect 3278 6872 3279 6873
rect 3059 6874 3060 6875
rect 3081 6874 3082 6875
rect 3066 6876 3067 6877
rect 3291 6876 3292 6877
rect 3065 6878 3066 6879
rect 3087 6878 3088 6879
rect 3071 6880 3072 6881
rect 3290 6880 3291 6881
rect 3077 6882 3078 6883
rect 3099 6882 3100 6883
rect 3086 6884 3087 6885
rect 3111 6884 3112 6885
rect 3092 6886 3093 6887
rect 3324 6886 3325 6887
rect 3101 6888 3102 6889
rect 3132 6888 3133 6889
rect 3119 6890 3120 6891
rect 3150 6890 3151 6891
rect 3143 6892 3144 6893
rect 3174 6892 3175 6893
rect 3149 6894 3150 6895
rect 3156 6894 3157 6895
rect 3167 6894 3168 6895
rect 3210 6894 3211 6895
rect 3173 6896 3174 6897
rect 3216 6896 3217 6897
rect 3179 6898 3180 6899
rect 3192 6898 3193 6899
rect 2928 6900 2929 6901
rect 3191 6900 3192 6901
rect 2929 6902 2930 6903
rect 3248 6902 3249 6903
rect 3182 6904 3183 6905
rect 3195 6904 3196 6905
rect 3084 6906 3085 6907
rect 3194 6906 3195 6907
rect 3083 6908 3084 6909
rect 3108 6908 3109 6909
rect 3107 6910 3108 6911
rect 3126 6910 3127 6911
rect 3125 6912 3126 6913
rect 3162 6912 3163 6913
rect 3161 6914 3162 6915
rect 3204 6914 3205 6915
rect 2903 6916 2904 6917
rect 3203 6916 3204 6917
rect 3189 6918 3190 6919
rect 3345 6918 3346 6919
rect 3206 6920 3207 6921
rect 3270 6920 3271 6921
rect 3212 6922 3213 6923
rect 3222 6922 3223 6923
rect 3215 6924 3216 6925
rect 3225 6924 3226 6925
rect 2974 6926 2975 6927
rect 3224 6926 3225 6927
rect 3218 6928 3219 6929
rect 3276 6928 3277 6929
rect 3230 6930 3231 6931
rect 3240 6930 3241 6931
rect 3234 6932 3235 6933
rect 3314 6932 3315 6933
rect 3233 6934 3234 6935
rect 3267 6934 3268 6935
rect 3236 6936 3237 6937
rect 3246 6936 3247 6937
rect 3266 6936 3267 6937
rect 3282 6936 3283 6937
rect 3272 6938 3273 6939
rect 3288 6938 3289 6939
rect 3165 6940 3166 6941
rect 3287 6940 3288 6941
rect 3300 6940 3301 6941
rect 3308 6940 3309 6941
rect 3228 6942 3229 6943
rect 3299 6942 3300 6943
rect 3227 6944 3228 6945
rect 3261 6944 3262 6945
rect 3318 6944 3319 6945
rect 3326 6944 3327 6945
rect 3323 6946 3324 6947
rect 3675 6946 3676 6947
rect 3330 6948 3331 6949
rect 3338 6948 3339 6949
rect 3321 6950 3322 6951
rect 3329 6950 3330 6951
rect 3312 6952 3313 6953
rect 3320 6952 3321 6953
rect 3303 6954 3304 6955
rect 3311 6954 3312 6955
rect 3294 6956 3295 6957
rect 3302 6956 3303 6957
rect 3342 6956 3343 6957
rect 3344 6956 3345 6957
rect 3333 6958 3334 6959
rect 3341 6958 3342 6959
rect 3296 6960 3297 6961
rect 3332 6960 3333 6961
rect 3348 6960 3349 6961
rect 3353 6960 3354 6961
rect 3063 6962 3064 6963
rect 3347 6962 3348 6963
rect 3402 6962 3403 6963
rect 3834 6962 3835 6963
rect 3372 6964 3373 6965
rect 3401 6964 3402 6965
rect 3366 6966 3367 6967
rect 3371 6966 3372 6967
rect 3360 6968 3361 6969
rect 3365 6968 3366 6969
rect 3408 6968 3409 6969
rect 3413 6968 3414 6969
rect 3426 6968 3427 6969
rect 3788 6968 3789 6969
rect 3390 6970 3391 6971
rect 3425 6970 3426 6971
rect 3378 6972 3379 6973
rect 3389 6972 3390 6973
rect 3336 6974 3337 6975
rect 3377 6974 3378 6975
rect 3335 6976 3336 6977
rect 3474 6976 3475 6977
rect 3441 6978 3442 6979
rect 3464 6978 3465 6979
rect 3456 6980 3457 6981
rect 3810 6980 3811 6981
rect 3450 6982 3451 6983
rect 3455 6982 3456 6983
rect 3473 6982 3474 6983
rect 3862 6982 3863 6983
rect 3480 6984 3481 6985
rect 3485 6984 3486 6985
rect 3468 6986 3469 6987
rect 3479 6986 3480 6987
rect 3462 6988 3463 6989
rect 3467 6988 3468 6989
rect 3438 6990 3439 6991
rect 3461 6990 3462 6991
rect 3432 6992 3433 6993
rect 3437 6992 3438 6993
rect 3396 6994 3397 6995
rect 3431 6994 3432 6995
rect 3384 6996 3385 6997
rect 3395 6996 3396 6997
rect 3383 6998 3384 6999
rect 3614 6998 3615 6999
rect 3489 7000 3490 7001
rect 3840 7000 3841 7001
rect 3494 7002 3495 7003
rect 3672 7002 3673 7003
rect 3501 7004 3502 7005
rect 3512 7004 3513 7005
rect 3522 7004 3523 7005
rect 3530 7004 3531 7005
rect 3524 7006 3525 7007
rect 3669 7006 3670 7007
rect 3528 7008 3529 7009
rect 3542 7008 3543 7009
rect 3534 7010 3535 7011
rect 3548 7010 3549 7011
rect 3536 7012 3537 7013
rect 3576 7012 3577 7013
rect 3546 7014 3547 7015
rect 3560 7014 3561 7015
rect 3552 7016 3553 7017
rect 3566 7016 3567 7017
rect 3564 7018 3565 7019
rect 3575 7018 3576 7019
rect 3572 7020 3573 7021
rect 3705 7020 3706 7021
rect 3591 7022 3592 7023
rect 3654 7022 3655 7023
rect 3420 7024 3421 7025
rect 3590 7024 3591 7025
rect 3419 7026 3420 7027
rect 3585 7026 3586 7027
rect 3600 7026 3601 7027
rect 3728 7026 3729 7027
rect 3594 7028 3595 7029
rect 3599 7028 3600 7029
rect 3603 7028 3604 7029
rect 3623 7028 3624 7029
rect 3597 7030 3598 7031
rect 3602 7030 3603 7031
rect 3627 7030 3628 7031
rect 3653 7030 3654 7031
rect 3630 7032 3631 7033
rect 3656 7032 3657 7033
rect 3633 7034 3634 7035
rect 3873 7034 3874 7035
rect 3639 7036 3640 7037
rect 3647 7036 3648 7037
rect 3666 7036 3667 7037
rect 3683 7036 3684 7037
rect 3645 7038 3646 7039
rect 3665 7038 3666 7039
rect 3686 7038 3687 7039
rect 3777 7038 3778 7039
rect 3507 7040 3508 7041
rect 3778 7040 3779 7041
rect 3506 7042 3507 7043
rect 3817 7042 3818 7043
rect 3693 7044 3694 7045
rect 3716 7044 3717 7045
rect 2951 7046 2952 7047
rect 3692 7046 3693 7047
rect 3696 7046 3697 7047
rect 3707 7046 3708 7047
rect 3678 7048 3679 7049
rect 3695 7048 3696 7049
rect 3699 7048 3700 7049
rect 3710 7048 3711 7049
rect 3702 7050 3703 7051
rect 3843 7050 3844 7051
rect 3720 7052 3721 7053
rect 3781 7052 3782 7053
rect 3719 7054 3720 7055
rect 3830 7054 3831 7055
rect 3407 7056 3408 7057
rect 3831 7056 3832 7057
rect 3722 7058 3723 7059
rect 3836 7058 3837 7059
rect 3726 7060 3727 7061
rect 3784 7060 3785 7061
rect 3609 7062 3610 7063
rect 3725 7062 3726 7063
rect 3747 7062 3748 7063
rect 3824 7062 3825 7063
rect 3756 7064 3757 7065
rect 3781 7064 3782 7065
rect 3617 7066 3618 7067
rect 3755 7066 3756 7067
rect 3765 7066 3766 7067
rect 3807 7066 3808 7067
rect 3753 7068 3754 7069
rect 3808 7068 3809 7069
rect 3732 7070 3733 7071
rect 3752 7070 3753 7071
rect 3714 7072 3715 7073
rect 3731 7072 3732 7073
rect 3690 7074 3691 7075
rect 3713 7074 3714 7075
rect 3663 7076 3664 7077
rect 3689 7076 3690 7077
rect 3775 7076 3776 7077
rect 3866 7076 3867 7077
rect 3794 7078 3795 7079
rect 3799 7078 3800 7079
rect 3768 7080 3769 7081
rect 3793 7080 3794 7081
rect 3797 7080 3798 7081
rect 3802 7080 3803 7081
rect 3771 7082 3772 7083
rect 3796 7082 3797 7083
rect 3621 7084 3622 7085
rect 3772 7084 3773 7085
rect 3811 7084 3812 7085
rect 3850 7084 3851 7085
rect 3814 7086 3815 7087
rect 3827 7086 3828 7087
rect 3582 7088 3583 7089
rect 3814 7088 3815 7089
rect 3570 7090 3571 7091
rect 3581 7090 3582 7091
rect 3555 7092 3556 7093
rect 3569 7092 3570 7093
rect 3540 7094 3541 7095
rect 3554 7094 3555 7095
rect 3854 7094 3855 7095
rect 3864 7094 3865 7095
rect 2893 7103 2894 7104
rect 3203 7103 3204 7104
rect 2908 7105 2909 7106
rect 3204 7105 3205 7106
rect 2911 7107 2912 7108
rect 2963 7107 2964 7108
rect 2915 7109 2916 7110
rect 3101 7109 3102 7110
rect 2919 7111 2920 7112
rect 3194 7111 3195 7112
rect 2918 7113 2919 7114
rect 3083 7113 3084 7114
rect 2921 7115 2922 7116
rect 3077 7115 3078 7116
rect 2926 7117 2927 7118
rect 3251 7117 3252 7118
rect 2925 7119 2926 7120
rect 3248 7119 3249 7120
rect 2928 7121 2929 7122
rect 3105 7121 3106 7122
rect 2950 7123 2951 7124
rect 3189 7123 3190 7124
rect 2954 7125 2955 7126
rect 3191 7125 3192 7126
rect 2956 7127 2957 7128
rect 2966 7127 2967 7128
rect 2959 7129 2960 7130
rect 3081 7129 3082 7130
rect 2969 7131 2970 7132
rect 3096 7131 3097 7132
rect 2969 7133 2970 7134
rect 3461 7133 3462 7134
rect 2972 7135 2973 7136
rect 3227 7135 3228 7136
rect 2973 7137 2974 7138
rect 3236 7137 3237 7138
rect 2966 7139 2967 7140
rect 3237 7139 3238 7140
rect 2976 7141 2977 7142
rect 3113 7141 3114 7142
rect 2985 7143 2986 7144
rect 3306 7143 3307 7144
rect 2995 7145 2996 7146
rect 3093 7145 3094 7146
rect 2994 7147 2995 7148
rect 3010 7147 3011 7148
rect 3000 7149 3001 7150
rect 3004 7149 3005 7150
rect 3006 7149 3007 7150
rect 3063 7149 3064 7150
rect 3009 7151 3010 7152
rect 3254 7151 3255 7152
rect 3022 7153 3023 7154
rect 3258 7153 3259 7154
rect 3030 7155 3031 7156
rect 3065 7155 3066 7156
rect 3037 7157 3038 7158
rect 3272 7157 3273 7158
rect 2979 7159 2980 7160
rect 3036 7159 3037 7160
rect 2979 7161 2980 7162
rect 2982 7161 2983 7162
rect 3041 7161 3042 7162
rect 3161 7161 3162 7162
rect 3042 7163 3043 7164
rect 3320 7163 3321 7164
rect 3048 7165 3049 7166
rect 3059 7165 3060 7166
rect 3060 7167 3061 7168
rect 3165 7167 3166 7168
rect 3074 7169 3075 7170
rect 3338 7169 3339 7170
rect 3075 7171 3076 7172
rect 3311 7171 3312 7172
rect 3086 7173 3087 7174
rect 3240 7173 3241 7174
rect 3087 7175 3088 7176
rect 3314 7175 3315 7176
rect 3107 7177 3108 7178
rect 3677 7177 3678 7178
rect 3111 7179 3112 7180
rect 3119 7179 3120 7180
rect 3117 7181 3118 7182
rect 3125 7181 3126 7182
rect 3123 7183 3124 7184
rect 3149 7183 3150 7184
rect 3129 7185 3130 7186
rect 3278 7185 3279 7186
rect 3143 7187 3144 7188
rect 3153 7187 3154 7188
rect 3147 7189 3148 7190
rect 3215 7189 3216 7190
rect 3167 7191 3168 7192
rect 3177 7191 3178 7192
rect 3171 7193 3172 7194
rect 3179 7193 3180 7194
rect 3173 7195 3174 7196
rect 3195 7195 3196 7196
rect 3174 7197 3175 7198
rect 3182 7197 3183 7198
rect 3197 7197 3198 7198
rect 3261 7197 3262 7198
rect 3200 7199 3201 7200
rect 3425 7199 3426 7200
rect 3201 7201 3202 7202
rect 3212 7201 3213 7202
rect 3206 7203 3207 7204
rect 3213 7203 3214 7204
rect 3057 7205 3058 7206
rect 3207 7205 3208 7206
rect 3222 7205 3223 7206
rect 3233 7205 3234 7206
rect 3224 7207 3225 7208
rect 3743 7207 3744 7208
rect 3218 7209 3219 7210
rect 3225 7209 3226 7210
rect 3219 7211 3220 7212
rect 3230 7211 3231 7212
rect 3231 7213 3232 7214
rect 3329 7213 3330 7214
rect 3071 7215 3072 7216
rect 3330 7215 3331 7216
rect 3242 7217 3243 7218
rect 3255 7217 3256 7218
rect 3089 7219 3090 7220
rect 3243 7219 3244 7220
rect 3246 7219 3247 7220
rect 3341 7219 3342 7220
rect 3144 7221 3145 7222
rect 3342 7221 3343 7222
rect 3287 7223 3288 7224
rect 3294 7223 3295 7224
rect 3288 7225 3289 7226
rect 3344 7225 3345 7226
rect 3299 7227 3300 7228
rect 3312 7227 3313 7228
rect 3302 7229 3303 7230
rect 3315 7229 3316 7230
rect 3303 7231 3304 7232
rect 3308 7231 3309 7232
rect 3296 7233 3297 7234
rect 3309 7233 3310 7234
rect 3290 7235 3291 7236
rect 3297 7235 3298 7236
rect 3284 7237 3285 7238
rect 3291 7237 3292 7238
rect 3132 7239 3133 7240
rect 3285 7239 3286 7240
rect 3318 7239 3319 7240
rect 3323 7239 3324 7240
rect 3321 7241 3322 7242
rect 3335 7241 3336 7242
rect 3333 7243 3334 7244
rect 3602 7243 3603 7244
rect 3339 7245 3340 7246
rect 3347 7245 3348 7246
rect 3345 7247 3346 7248
rect 3383 7247 3384 7248
rect 3348 7249 3349 7250
rect 3599 7249 3600 7250
rect 3351 7251 3352 7252
rect 3389 7251 3390 7252
rect 3353 7253 3354 7254
rect 3736 7253 3737 7254
rect 3357 7255 3358 7256
rect 3377 7255 3378 7256
rect 3363 7257 3364 7258
rect 3365 7257 3366 7258
rect 3369 7257 3370 7258
rect 3371 7257 3372 7258
rect 3381 7257 3382 7258
rect 3590 7257 3591 7258
rect 3393 7259 3394 7260
rect 3494 7259 3495 7260
rect 3399 7261 3400 7262
rect 3413 7261 3414 7262
rect 3401 7263 3402 7264
rect 3611 7263 3612 7264
rect 3405 7265 3406 7266
rect 3407 7265 3408 7266
rect 3411 7265 3412 7266
rect 3762 7265 3763 7266
rect 3423 7267 3424 7268
rect 3536 7267 3537 7268
rect 3429 7269 3430 7270
rect 3455 7269 3456 7270
rect 3431 7271 3432 7272
rect 3746 7271 3747 7272
rect 3435 7273 3436 7274
rect 3817 7273 3818 7274
rect 3437 7275 3438 7276
rect 3765 7275 3766 7276
rect 3441 7277 3442 7278
rect 3710 7277 3711 7278
rect 3450 7279 3451 7280
rect 3467 7279 3468 7280
rect 3456 7281 3457 7282
rect 3569 7281 3570 7282
rect 3462 7283 3463 7284
rect 3772 7283 3773 7284
rect 3464 7285 3465 7286
rect 3703 7285 3704 7286
rect 3395 7287 3396 7288
rect 3465 7287 3466 7288
rect 3468 7287 3469 7288
rect 3542 7287 3543 7288
rect 3473 7289 3474 7290
rect 3866 7289 3867 7290
rect 3474 7291 3475 7292
rect 3485 7291 3486 7292
rect 3477 7293 3478 7294
rect 3512 7293 3513 7294
rect 3479 7295 3480 7296
rect 3862 7295 3863 7296
rect 3483 7297 3484 7298
rect 3778 7297 3779 7298
rect 3489 7299 3490 7300
rect 3575 7299 3576 7300
rect 3501 7301 3502 7302
rect 3530 7301 3531 7302
rect 3513 7303 3514 7304
rect 3728 7303 3729 7304
rect 3506 7305 3507 7306
rect 3729 7305 3730 7306
rect 3507 7307 3508 7308
rect 3560 7307 3561 7308
rect 3519 7309 3520 7310
rect 3572 7309 3573 7310
rect 3522 7311 3523 7312
rect 3581 7311 3582 7312
rect 3528 7313 3529 7314
rect 3617 7313 3618 7314
rect 3534 7315 3535 7316
rect 3805 7315 3806 7316
rect 3537 7317 3538 7318
rect 3566 7317 3567 7318
rect 3546 7319 3547 7320
rect 3686 7319 3687 7320
rect 3552 7321 3553 7322
rect 3653 7321 3654 7322
rect 3554 7323 3555 7324
rect 3651 7323 3652 7324
rect 3555 7325 3556 7326
rect 3656 7325 3657 7326
rect 3564 7327 3565 7328
rect 3722 7327 3723 7328
rect 3582 7329 3583 7330
rect 3658 7329 3659 7330
rect 3587 7331 3588 7332
rect 3758 7331 3759 7332
rect 3600 7333 3601 7334
rect 3713 7333 3714 7334
rect 3603 7335 3604 7336
rect 3716 7335 3717 7336
rect 3606 7337 3607 7338
rect 3689 7337 3690 7338
rect 3609 7339 3610 7340
rect 3692 7339 3693 7340
rect 3618 7341 3619 7342
rect 3695 7341 3696 7342
rect 3623 7343 3624 7344
rect 3859 7343 3860 7344
rect 3624 7345 3625 7346
rect 3719 7345 3720 7346
rect 3419 7347 3420 7348
rect 3719 7347 3720 7348
rect 3627 7349 3628 7350
rect 3852 7349 3853 7350
rect 3636 7351 3637 7352
rect 3749 7351 3750 7352
rect 3639 7353 3640 7354
rect 3731 7353 3732 7354
rect 3642 7355 3643 7356
rect 3655 7355 3656 7356
rect 3645 7357 3646 7358
rect 3725 7357 3726 7358
rect 3661 7359 3662 7360
rect 3799 7359 3800 7360
rect 3665 7361 3666 7362
rect 3764 7361 3765 7362
rect 3647 7363 3648 7364
rect 3664 7363 3665 7364
rect 3387 7365 3388 7366
rect 3648 7365 3649 7366
rect 3667 7365 3668 7366
rect 3683 7365 3684 7366
rect 3680 7367 3681 7368
rect 3802 7367 3803 7368
rect 3679 7369 3680 7370
rect 3775 7369 3776 7370
rect 3682 7371 3683 7372
rect 3771 7371 3772 7372
rect 3685 7373 3686 7374
rect 3781 7373 3782 7374
rect 3697 7375 3698 7376
rect 3793 7375 3794 7376
rect 3700 7377 3701 7378
rect 3796 7377 3797 7378
rect 3707 7379 3708 7380
rect 3841 7379 3842 7380
rect 3548 7381 3549 7382
rect 3706 7381 3707 7382
rect 3524 7383 3525 7384
rect 3549 7383 3550 7384
rect 3716 7383 3717 7384
rect 3811 7383 3812 7384
rect 3752 7385 3753 7386
rect 3755 7385 3756 7386
rect 3757 7385 3758 7386
rect 3838 7385 3839 7386
rect 3814 7387 3815 7388
rect 3820 7387 3821 7388
rect 2911 7396 2912 7397
rect 2956 7396 2957 7397
rect 2918 7398 2919 7399
rect 3000 7398 3001 7399
rect 2928 7400 2929 7401
rect 3255 7400 3256 7401
rect 2935 7402 2936 7403
rect 3189 7402 3190 7403
rect 2962 7404 2963 7405
rect 3345 7404 3346 7405
rect 2962 7406 2963 7407
rect 3333 7406 3334 7407
rect 2966 7408 2967 7409
rect 3291 7408 3292 7409
rect 2969 7410 2970 7411
rect 3315 7410 3316 7411
rect 2969 7412 2970 7413
rect 3036 7412 3037 7413
rect 2925 7414 2926 7415
rect 3035 7414 3036 7415
rect 2973 7416 2974 7417
rect 3004 7416 3005 7417
rect 2979 7418 2980 7419
rect 2989 7418 2990 7419
rect 2985 7420 2986 7421
rect 3294 7420 3295 7421
rect 2979 7422 2980 7423
rect 2986 7422 2987 7423
rect 2994 7422 2995 7423
rect 3135 7422 3136 7423
rect 3006 7424 3007 7425
rect 3252 7424 3253 7425
rect 3007 7426 3008 7427
rect 3050 7426 3051 7427
rect 3009 7428 3010 7429
rect 3231 7428 3232 7429
rect 3017 7430 3018 7431
rect 3045 7430 3046 7431
rect 3038 7432 3039 7433
rect 3258 7432 3259 7433
rect 3042 7434 3043 7435
rect 3411 7434 3412 7435
rect 3030 7436 3031 7437
rect 3041 7436 3042 7437
rect 3054 7436 3055 7437
rect 3090 7436 3091 7437
rect 2953 7438 2954 7439
rect 3090 7438 3091 7439
rect 3057 7440 3058 7441
rect 3330 7440 3331 7441
rect 3057 7442 3058 7443
rect 3168 7442 3169 7443
rect 3063 7444 3064 7445
rect 3078 7444 3079 7445
rect 3075 7446 3076 7447
rect 3102 7446 3103 7447
rect 3093 7448 3094 7449
rect 3108 7448 3109 7449
rect 3105 7450 3106 7451
rect 3120 7450 3121 7451
rect 3111 7452 3112 7453
rect 3126 7452 3127 7453
rect 3096 7454 3097 7455
rect 3111 7454 3112 7455
rect 3081 7456 3082 7457
rect 3096 7456 3097 7457
rect 3114 7456 3115 7457
rect 3417 7456 3418 7457
rect 3123 7458 3124 7459
rect 3138 7458 3139 7459
rect 3129 7460 3130 7461
rect 3243 7460 3244 7461
rect 3132 7462 3133 7463
rect 3399 7462 3400 7463
rect 3117 7464 3118 7465
rect 3132 7464 3133 7465
rect 3147 7464 3148 7465
rect 3150 7464 3151 7465
rect 3153 7464 3154 7465
rect 3156 7464 3157 7465
rect 3165 7464 3166 7465
rect 3315 7464 3316 7465
rect 3171 7466 3172 7467
rect 3186 7466 3187 7467
rect 3171 7468 3172 7469
rect 3246 7468 3247 7469
rect 3174 7470 3175 7471
rect 3189 7470 3190 7471
rect 2958 7472 2959 7473
rect 3174 7472 3175 7473
rect 3177 7472 3178 7473
rect 3210 7472 3211 7473
rect 3048 7474 3049 7475
rect 3177 7474 3178 7475
rect 3047 7476 3048 7477
rect 3300 7476 3301 7477
rect 3192 7478 3193 7479
rect 3195 7478 3196 7479
rect 3207 7478 3208 7479
rect 3258 7478 3259 7479
rect 3213 7480 3214 7481
rect 3228 7480 3229 7481
rect 3219 7482 3220 7483
rect 3246 7482 3247 7483
rect 2914 7484 2915 7485
rect 3219 7484 3220 7485
rect 2914 7486 2915 7487
rect 3216 7486 3217 7487
rect 3222 7486 3223 7487
rect 3249 7486 3250 7487
rect 3201 7488 3202 7489
rect 3222 7488 3223 7489
rect 3234 7488 3235 7489
rect 3237 7488 3238 7489
rect 3237 7490 3238 7491
rect 3240 7490 3241 7491
rect 3225 7492 3226 7493
rect 3240 7492 3241 7493
rect 3204 7494 3205 7495
rect 3225 7494 3226 7495
rect 2932 7496 2933 7497
rect 3204 7496 3205 7497
rect 3243 7496 3244 7497
rect 3318 7496 3319 7497
rect 3261 7498 3262 7499
rect 3276 7498 3277 7499
rect 3267 7500 3268 7501
rect 3270 7500 3271 7501
rect 3144 7502 3145 7503
rect 3267 7502 3268 7503
rect 3282 7502 3283 7503
rect 3297 7502 3298 7503
rect 3285 7504 3286 7505
rect 3345 7504 3346 7505
rect 3291 7506 3292 7507
rect 3306 7506 3307 7507
rect 3294 7508 3295 7509
rect 3309 7508 3310 7509
rect 3297 7510 3298 7511
rect 3312 7510 3313 7511
rect 3306 7512 3307 7513
rect 3321 7512 3322 7513
rect 3312 7514 3313 7515
rect 3327 7514 3328 7515
rect 3318 7516 3319 7517
rect 3330 7516 3331 7517
rect 3342 7516 3343 7517
rect 3360 7516 3361 7517
rect 3288 7518 3289 7519
rect 3342 7518 3343 7519
rect 3288 7520 3289 7521
rect 3303 7520 3304 7521
rect 3348 7520 3349 7521
rect 3384 7520 3385 7521
rect 3348 7522 3349 7523
rect 3363 7522 3364 7523
rect 3339 7524 3340 7525
rect 3363 7524 3364 7525
rect 3351 7526 3352 7527
rect 3372 7526 3373 7527
rect 3354 7528 3355 7529
rect 3357 7528 3358 7529
rect 3369 7528 3370 7529
rect 3736 7528 3737 7529
rect 3387 7530 3388 7531
rect 3414 7530 3415 7531
rect 3381 7532 3382 7533
rect 3387 7532 3388 7533
rect 3390 7532 3391 7533
rect 3405 7532 3406 7533
rect 3393 7534 3394 7535
rect 3408 7534 3409 7535
rect 3396 7536 3397 7537
rect 3558 7536 3559 7537
rect 3399 7538 3400 7539
rect 3465 7538 3466 7539
rect 3402 7540 3403 7541
rect 3719 7540 3720 7541
rect 3420 7542 3421 7543
rect 3549 7542 3550 7543
rect 3426 7544 3427 7545
rect 3441 7544 3442 7545
rect 3435 7546 3436 7547
rect 3441 7546 3442 7547
rect 3429 7548 3430 7549
rect 3435 7548 3436 7549
rect 3423 7550 3424 7551
rect 3429 7550 3430 7551
rect 3447 7550 3448 7551
rect 3456 7550 3457 7551
rect 3453 7552 3454 7553
rect 3468 7552 3469 7553
rect 3459 7554 3460 7555
rect 3474 7554 3475 7555
rect 3462 7556 3463 7557
rect 3561 7556 3562 7557
rect 3462 7558 3463 7559
rect 3710 7558 3711 7559
rect 3468 7560 3469 7561
rect 3528 7560 3529 7561
rect 3477 7562 3478 7563
rect 3480 7562 3481 7563
rect 3483 7562 3484 7563
rect 3486 7562 3487 7563
rect 3489 7562 3490 7563
rect 3648 7562 3649 7563
rect 3510 7564 3511 7565
rect 3704 7564 3705 7565
rect 3513 7566 3514 7567
rect 3622 7566 3623 7567
rect 3525 7568 3526 7569
rect 3534 7568 3535 7569
rect 3528 7570 3529 7571
rect 3537 7570 3538 7571
rect 3537 7572 3538 7573
rect 3629 7572 3630 7573
rect 3540 7574 3541 7575
rect 3546 7574 3547 7575
rect 3543 7576 3544 7577
rect 3552 7576 3553 7577
rect 3546 7578 3547 7579
rect 3555 7578 3556 7579
rect 3561 7578 3562 7579
rect 3664 7578 3665 7579
rect 3573 7580 3574 7581
rect 3582 7580 3583 7581
rect 3579 7582 3580 7583
rect 3600 7582 3601 7583
rect 3582 7584 3583 7585
rect 3603 7584 3604 7585
rect 3564 7586 3565 7587
rect 3603 7586 3604 7587
rect 3507 7588 3508 7589
rect 3564 7588 3565 7589
rect 3507 7590 3508 7591
rect 3519 7590 3520 7591
rect 3585 7590 3586 7591
rect 3609 7590 3610 7591
rect 3594 7592 3595 7593
rect 3618 7592 3619 7593
rect 3576 7594 3577 7595
rect 3619 7594 3620 7595
rect 3600 7596 3601 7597
rect 3624 7596 3625 7597
rect 3606 7598 3607 7599
rect 3781 7598 3782 7599
rect 3606 7600 3607 7601
rect 3639 7600 3640 7601
rect 3450 7602 3451 7603
rect 3640 7602 3641 7603
rect 3609 7604 3610 7605
rect 3729 7604 3730 7605
rect 3612 7606 3613 7607
rect 3661 7606 3662 7607
rect 3627 7608 3628 7609
rect 3725 7608 3726 7609
rect 3633 7610 3634 7611
rect 3636 7610 3637 7611
rect 3642 7610 3643 7611
rect 3658 7610 3659 7611
rect 3645 7612 3646 7613
rect 3655 7612 3656 7613
rect 3643 7614 3644 7615
rect 3655 7614 3656 7615
rect 3652 7616 3653 7617
rect 3716 7616 3717 7617
rect 3658 7618 3659 7619
rect 3685 7618 3686 7619
rect 3670 7620 3671 7621
rect 3722 7620 3723 7621
rect 3522 7622 3523 7623
rect 3721 7622 3722 7623
rect 3670 7624 3671 7625
rect 3697 7624 3698 7625
rect 3673 7626 3674 7627
rect 3700 7626 3701 7627
rect 3679 7628 3680 7629
rect 3774 7628 3775 7629
rect 3321 7630 3322 7631
rect 3679 7630 3680 7631
rect 3682 7630 3683 7631
rect 3727 7630 3728 7631
rect 3743 7630 3744 7631
rect 3760 7630 3761 7631
rect 2809 7639 2810 7640
rect 3447 7639 3448 7640
rect 2888 7641 2889 7642
rect 2894 7641 2895 7642
rect 2924 7641 2925 7642
rect 3060 7641 3061 7642
rect 2928 7643 2929 7644
rect 3038 7643 3039 7644
rect 2931 7645 2932 7646
rect 3219 7645 3220 7646
rect 2964 7647 2965 7648
rect 3273 7647 3274 7648
rect 2967 7649 2968 7650
rect 3246 7649 3247 7650
rect 2969 7651 2970 7652
rect 3041 7651 3042 7652
rect 2972 7653 2973 7654
rect 3017 7653 3018 7654
rect 2986 7655 2987 7656
rect 3321 7655 3322 7656
rect 2989 7657 2990 7658
rect 3013 7657 3014 7658
rect 3035 7657 3036 7658
rect 3063 7657 3064 7658
rect 3039 7659 3040 7660
rect 3405 7659 3406 7660
rect 3050 7661 3051 7662
rect 3276 7661 3277 7662
rect 3057 7663 3058 7664
rect 3144 7663 3145 7664
rect 2960 7665 2961 7666
rect 3144 7665 3145 7666
rect 3072 7667 3073 7668
rect 3078 7667 3079 7668
rect 3078 7669 3079 7670
rect 3114 7669 3115 7670
rect 3084 7671 3085 7672
rect 3102 7671 3103 7672
rect 3102 7673 3103 7674
rect 3108 7673 3109 7674
rect 3105 7675 3106 7676
rect 3111 7675 3112 7676
rect 3108 7677 3109 7678
rect 3138 7677 3139 7678
rect 3114 7679 3115 7680
rect 3132 7679 3133 7680
rect 3117 7681 3118 7682
rect 3135 7681 3136 7682
rect 3120 7683 3121 7684
rect 3138 7683 3139 7684
rect 3123 7685 3124 7686
rect 3351 7685 3352 7686
rect 3129 7687 3130 7688
rect 3171 7687 3172 7688
rect 3156 7689 3157 7690
rect 3180 7689 3181 7690
rect 2957 7691 2958 7692
rect 3156 7691 3157 7692
rect 3165 7691 3166 7692
rect 3363 7691 3364 7692
rect 3174 7693 3175 7694
rect 3198 7693 3199 7694
rect 3177 7695 3178 7696
rect 3201 7695 3202 7696
rect 3189 7697 3190 7698
rect 3213 7697 3214 7698
rect 3204 7699 3205 7700
rect 3318 7699 3319 7700
rect 3216 7701 3217 7702
rect 3264 7701 3265 7702
rect 3192 7703 3193 7704
rect 3216 7703 3217 7704
rect 3219 7703 3220 7704
rect 3249 7703 3250 7704
rect 3222 7705 3223 7706
rect 3246 7705 3247 7706
rect 3210 7707 3211 7708
rect 3222 7707 3223 7708
rect 3186 7709 3187 7710
rect 3210 7709 3211 7710
rect 3225 7709 3226 7710
rect 3249 7709 3250 7710
rect 3234 7711 3235 7712
rect 3285 7711 3286 7712
rect 3234 7713 3235 7714
rect 3240 7713 3241 7714
rect 3029 7715 3030 7716
rect 3240 7715 3241 7716
rect 3252 7715 3253 7716
rect 3267 7715 3268 7716
rect 3252 7717 3253 7718
rect 3258 7717 3259 7718
rect 3270 7717 3271 7718
rect 3309 7717 3310 7718
rect 3282 7719 3283 7720
rect 3333 7719 3334 7720
rect 3288 7721 3289 7722
rect 3357 7721 3358 7722
rect 2921 7723 2922 7724
rect 3288 7723 3289 7724
rect 2920 7725 2921 7726
rect 3016 7725 3017 7726
rect 3294 7725 3295 7726
rect 3339 7725 3340 7726
rect 3300 7727 3301 7728
rect 3303 7727 3304 7728
rect 3312 7727 3313 7728
rect 3363 7727 3364 7728
rect 3327 7729 3328 7730
rect 3345 7729 3346 7730
rect 3306 7731 3307 7732
rect 3345 7731 3346 7732
rect 3330 7733 3331 7734
rect 3381 7733 3382 7734
rect 3348 7735 3349 7736
rect 3423 7735 3424 7736
rect 3369 7737 3370 7738
rect 3468 7737 3469 7738
rect 3372 7739 3373 7740
rect 3393 7739 3394 7740
rect 3375 7741 3376 7742
rect 3387 7741 3388 7742
rect 3032 7743 3033 7744
rect 3387 7743 3388 7744
rect 3390 7743 3391 7744
rect 3465 7743 3466 7744
rect 3315 7745 3316 7746
rect 3390 7745 3391 7746
rect 3399 7745 3400 7746
rect 3417 7745 3418 7746
rect 3354 7747 3355 7748
rect 3399 7747 3400 7748
rect 3342 7749 3343 7750
rect 3354 7749 3355 7750
rect 3297 7751 3298 7752
rect 3342 7751 3343 7752
rect 3297 7753 3298 7754
rect 3429 7753 3430 7754
rect 3402 7755 3403 7756
rect 3471 7755 3472 7756
rect 3411 7757 3412 7758
rect 3414 7757 3415 7758
rect 3384 7759 3385 7760
rect 3414 7759 3415 7760
rect 3420 7759 3421 7760
rect 3721 7759 3722 7760
rect 3396 7761 3397 7762
rect 3420 7761 3421 7762
rect 3426 7761 3427 7762
rect 3495 7761 3496 7762
rect 3426 7763 3427 7764
rect 3546 7763 3547 7764
rect 3429 7765 3430 7766
rect 3462 7765 3463 7766
rect 3435 7767 3436 7768
rect 3665 7767 3666 7768
rect 3435 7769 3436 7770
rect 3453 7769 3454 7770
rect 3441 7771 3442 7772
rect 3477 7771 3478 7772
rect 3162 7773 3163 7774
rect 3441 7773 3442 7774
rect 3447 7773 3448 7774
rect 3650 7773 3651 7774
rect 3459 7775 3460 7776
rect 3522 7775 3523 7776
rect 3459 7777 3460 7778
rect 3640 7777 3641 7778
rect 3453 7779 3454 7780
rect 3639 7779 3640 7780
rect 3486 7781 3487 7782
rect 3633 7781 3634 7782
rect 3504 7783 3505 7784
rect 3712 7783 3713 7784
rect 3510 7785 3511 7786
rect 3700 7785 3701 7786
rect 3150 7787 3151 7788
rect 3510 7787 3511 7788
rect 3126 7789 3127 7790
rect 3150 7789 3151 7790
rect 3126 7791 3127 7792
rect 3168 7791 3169 7792
rect 3516 7791 3517 7792
rect 3707 7791 3708 7792
rect 3525 7793 3526 7794
rect 3552 7793 3553 7794
rect 3480 7795 3481 7796
rect 3525 7795 3526 7796
rect 3528 7795 3529 7796
rect 3555 7795 3556 7796
rect 3537 7797 3538 7798
rect 3567 7797 3568 7798
rect 3507 7799 3508 7800
rect 3537 7799 3538 7800
rect 3540 7799 3541 7800
rect 3619 7799 3620 7800
rect 3501 7801 3502 7802
rect 3540 7801 3541 7802
rect 3543 7801 3544 7802
rect 3597 7801 3598 7802
rect 3561 7803 3562 7804
rect 3588 7803 3589 7804
rect 3564 7805 3565 7806
rect 3591 7805 3592 7806
rect 3564 7807 3565 7808
rect 3629 7807 3630 7808
rect 3570 7809 3571 7810
rect 3573 7809 3574 7810
rect 3573 7811 3574 7812
rect 3576 7811 3577 7812
rect 3579 7811 3580 7812
rect 3695 7811 3696 7812
rect 3582 7813 3583 7814
rect 3662 7813 3663 7814
rect 3585 7815 3586 7816
rect 3727 7815 3728 7816
rect 3594 7817 3595 7818
rect 3618 7817 3619 7818
rect 3237 7819 3238 7820
rect 3594 7819 3595 7820
rect 3237 7821 3238 7822
rect 3243 7821 3244 7822
rect 3600 7821 3601 7822
rect 3624 7821 3625 7822
rect 3600 7823 3601 7824
rect 3609 7823 3610 7824
rect 3603 7825 3604 7826
rect 3627 7825 3628 7826
rect 3606 7827 3607 7828
rect 3615 7827 3616 7828
rect 3612 7829 3613 7830
rect 3636 7829 3637 7830
rect 3630 7831 3631 7832
rect 3730 7831 3731 7832
rect 3655 7833 3656 7834
rect 3702 7833 3703 7834
rect 3656 7835 3657 7836
rect 3733 7835 3734 7836
rect 3670 7837 3671 7838
rect 3689 7837 3690 7838
rect 3652 7839 3653 7840
rect 3671 7839 3672 7840
rect 3673 7839 3674 7840
rect 3692 7839 3693 7840
rect 3674 7841 3675 7842
rect 3686 7841 3687 7842
rect 3676 7843 3677 7844
rect 3705 7843 3706 7844
rect 3658 7845 3659 7846
rect 3677 7845 3678 7846
rect 3659 7847 3660 7848
rect 3679 7847 3680 7848
rect 2884 7856 2885 7857
rect 2894 7856 2895 7857
rect 2888 7858 2889 7859
rect 2917 7858 2918 7859
rect 2914 7860 2915 7861
rect 3063 7860 3064 7861
rect 2918 7862 2919 7863
rect 3285 7862 3286 7863
rect 2921 7864 2922 7865
rect 3198 7864 3199 7865
rect 2931 7866 2932 7867
rect 3006 7866 3007 7867
rect 2946 7868 2947 7869
rect 3288 7868 3289 7869
rect 2960 7870 2961 7871
rect 3138 7870 3139 7871
rect 2961 7872 2962 7873
rect 3108 7872 3109 7873
rect 2965 7874 2966 7875
rect 3267 7874 3268 7875
rect 2967 7876 2968 7877
rect 3234 7876 3235 7877
rect 2968 7878 2969 7879
rect 3129 7878 3130 7879
rect 2975 7880 2976 7881
rect 3136 7880 3137 7881
rect 2995 7882 2996 7883
rect 3213 7882 3214 7883
rect 2943 7884 2944 7885
rect 2994 7884 2995 7885
rect 2997 7884 2998 7885
rect 3013 7884 3014 7885
rect 3003 7886 3004 7887
rect 3345 7886 3346 7887
rect 3018 7888 3019 7889
rect 3390 7888 3391 7889
rect 3022 7890 3023 7891
rect 3156 7890 3157 7891
rect 3025 7892 3026 7893
rect 3268 7892 3269 7893
rect 3029 7894 3030 7895
rect 3385 7894 3386 7895
rect 3032 7896 3033 7897
rect 3331 7896 3332 7897
rect 3016 7898 3017 7899
rect 3031 7898 3032 7899
rect 3037 7898 3038 7899
rect 3540 7898 3541 7899
rect 3046 7900 3047 7901
rect 3391 7900 3392 7901
rect 3049 7902 3050 7903
rect 3235 7902 3236 7903
rect 3058 7904 3059 7905
rect 3078 7904 3079 7905
rect 3060 7906 3061 7907
rect 3064 7906 3065 7907
rect 3112 7906 3113 7907
rect 3399 7906 3400 7907
rect 3120 7908 3121 7909
rect 3327 7908 3328 7909
rect 3121 7910 3122 7911
rect 3144 7910 3145 7911
rect 3126 7912 3127 7913
rect 3133 7912 3134 7913
rect 3127 7914 3128 7915
rect 3150 7914 3151 7915
rect 3139 7916 3140 7917
rect 3643 7916 3644 7917
rect 3145 7918 3146 7919
rect 3180 7918 3181 7919
rect 3157 7920 3158 7921
rect 3210 7920 3211 7921
rect 3165 7922 3166 7923
rect 3303 7922 3304 7923
rect 3172 7924 3173 7925
rect 3216 7924 3217 7925
rect 3175 7926 3176 7927
rect 3219 7926 3220 7927
rect 3184 7928 3185 7929
rect 3240 7928 3241 7929
rect 3186 7930 3187 7931
rect 3367 7930 3368 7931
rect 3189 7932 3190 7933
rect 3375 7932 3376 7933
rect 3190 7934 3191 7935
rect 3246 7934 3247 7935
rect 3193 7936 3194 7937
rect 3249 7936 3250 7937
rect 3196 7938 3197 7939
rect 3222 7938 3223 7939
rect 3201 7940 3202 7941
rect 3484 7940 3485 7941
rect 3202 7942 3203 7943
rect 3228 7942 3229 7943
rect 3205 7944 3206 7945
rect 3237 7944 3238 7945
rect 3208 7946 3209 7947
rect 3264 7946 3265 7947
rect 3211 7948 3212 7949
rect 3273 7948 3274 7949
rect 3241 7950 3242 7951
rect 3426 7950 3427 7951
rect 3247 7952 3248 7953
rect 3309 7952 3310 7953
rect 3259 7954 3260 7955
rect 3420 7954 3421 7955
rect 3265 7956 3266 7957
rect 3351 7956 3352 7957
rect 3271 7958 3272 7959
rect 3333 7958 3334 7959
rect 3277 7960 3278 7961
rect 3297 7960 3298 7961
rect 3283 7962 3284 7963
rect 3339 7962 3340 7963
rect 3252 7964 3253 7965
rect 3340 7964 3341 7965
rect 3253 7966 3254 7967
rect 3354 7966 3355 7967
rect 3286 7968 3287 7969
rect 3342 7968 3343 7969
rect 3289 7970 3290 7971
rect 3321 7970 3322 7971
rect 3291 7972 3292 7973
rect 3646 7972 3647 7973
rect 3295 7974 3296 7975
rect 3393 7974 3394 7975
rect 3301 7976 3302 7977
rect 3357 7976 3358 7977
rect 3304 7978 3305 7979
rect 3360 7978 3361 7979
rect 3307 7980 3308 7981
rect 3363 7980 3364 7981
rect 3313 7982 3314 7983
rect 3417 7982 3418 7983
rect 3319 7984 3320 7985
rect 3381 7984 3382 7985
rect 3325 7986 3326 7987
rect 3487 7986 3488 7987
rect 3337 7988 3338 7989
rect 3387 7988 3388 7989
rect 3343 7990 3344 7991
rect 3369 7990 3370 7991
rect 3349 7992 3350 7993
rect 3535 7992 3536 7993
rect 3355 7994 3356 7995
rect 3405 7994 3406 7995
rect 3358 7996 3359 7997
rect 3408 7996 3409 7997
rect 3361 7998 3362 7999
rect 3411 7998 3412 7999
rect 3364 8000 3365 8001
rect 3414 8000 3415 8001
rect 3373 8002 3374 8003
rect 3423 8002 3424 8003
rect 3388 8004 3389 8005
rect 3441 8004 3442 8005
rect 3397 8006 3398 8007
rect 3453 8006 3454 8007
rect 3403 8008 3404 8009
rect 3459 8008 3460 8009
rect 3415 8010 3416 8011
rect 3465 8010 3466 8011
rect 3429 8012 3430 8013
rect 3653 8012 3654 8013
rect 3433 8014 3434 8015
rect 3552 8014 3553 8015
rect 3316 8016 3317 8017
rect 3552 8016 3553 8017
rect 3435 8018 3436 8019
rect 3650 8018 3651 8019
rect 3436 8020 3437 8021
rect 3555 8020 3556 8021
rect 3439 8022 3440 8023
rect 3504 8022 3505 8023
rect 3447 8024 3448 8025
rect 3639 8024 3640 8025
rect 3451 8026 3452 8027
rect 3537 8026 3538 8027
rect 3454 8028 3455 8029
rect 3674 8028 3675 8029
rect 3457 8030 3458 8031
rect 3471 8030 3472 8031
rect 3460 8032 3461 8033
rect 3594 8032 3595 8033
rect 3463 8034 3464 8035
rect 3597 8034 3598 8035
rect 3466 8036 3467 8037
rect 3525 8036 3526 8037
rect 3472 8038 3473 8039
rect 3522 8038 3523 8039
rect 3475 8040 3476 8041
rect 3633 8040 3634 8041
rect 3477 8042 3478 8043
rect 3668 8042 3669 8043
rect 3478 8044 3479 8045
rect 3570 8044 3571 8045
rect 3481 8046 3482 8047
rect 3573 8046 3574 8047
rect 3490 8048 3491 8049
rect 3642 8048 3643 8049
rect 3493 8050 3494 8051
rect 3600 8050 3601 8051
rect 3495 8052 3496 8053
rect 3572 8052 3573 8053
rect 3499 8054 3500 8055
rect 3627 8054 3628 8055
rect 3502 8056 3503 8057
rect 3603 8056 3604 8057
rect 3514 8058 3515 8059
rect 3665 8058 3666 8059
rect 3516 8060 3517 8061
rect 3733 8060 3734 8061
rect 3517 8062 3518 8063
rect 3588 8062 3589 8063
rect 3520 8064 3521 8065
rect 3662 8064 3663 8065
rect 3529 8066 3530 8067
rect 3612 8066 3613 8067
rect 3532 8068 3533 8069
rect 3615 8068 3616 8069
rect 3545 8070 3546 8071
rect 3567 8070 3568 8071
rect 3549 8072 3550 8073
rect 3659 8072 3660 8073
rect 3564 8074 3565 8075
rect 3600 8074 3601 8075
rect 3575 8076 3576 8077
rect 3677 8076 3678 8077
rect 3587 8078 3588 8079
rect 3689 8078 3690 8079
rect 3591 8080 3592 8081
rect 3712 8080 3713 8081
rect 3590 8082 3591 8083
rect 3692 8082 3693 8083
rect 3618 8084 3619 8085
rect 3740 8084 3741 8085
rect 3569 8086 3570 8087
rect 3617 8086 3618 8087
rect 3624 8086 3625 8087
rect 3716 8086 3717 8087
rect 3630 8088 3631 8089
rect 3747 8088 3748 8089
rect 3645 8090 3646 8091
rect 3666 8090 3667 8091
rect 3656 8092 3657 8093
rect 3754 8092 3755 8093
rect 3671 8094 3672 8095
rect 3705 8094 3706 8095
rect 3760 8094 3761 8095
rect 3764 8094 3765 8095
rect 2921 8103 2922 8104
rect 3208 8103 3209 8104
rect 2918 8105 2919 8106
rect 2920 8105 2921 8106
rect 2927 8105 2928 8106
rect 3304 8105 3305 8106
rect 2932 8107 2933 8108
rect 3085 8107 3086 8108
rect 2931 8109 2932 8110
rect 3145 8109 3146 8110
rect 2935 8111 2936 8112
rect 3091 8111 3092 8112
rect 2954 8113 2955 8114
rect 3103 8113 3104 8114
rect 2965 8115 2966 8116
rect 3227 8115 3228 8116
rect 2975 8117 2976 8118
rect 3106 8117 3107 8118
rect 2975 8119 2976 8120
rect 2997 8119 2998 8120
rect 2987 8121 2988 8122
rect 3271 8121 3272 8122
rect 2991 8123 2992 8124
rect 3046 8123 3047 8124
rect 2990 8125 2991 8126
rect 3283 8125 3284 8126
rect 2993 8127 2994 8128
rect 3340 8127 3341 8128
rect 3003 8129 3004 8130
rect 3006 8129 3007 8130
rect 3018 8129 3019 8130
rect 3319 8129 3320 8130
rect 3018 8131 3019 8132
rect 3307 8131 3308 8132
rect 3025 8133 3026 8134
rect 3263 8133 3264 8134
rect 3027 8135 3028 8136
rect 3188 8135 3189 8136
rect 3034 8137 3035 8138
rect 3235 8137 3236 8138
rect 3041 8139 3042 8140
rect 3218 8139 3219 8140
rect 3049 8141 3050 8142
rect 3200 8141 3201 8142
rect 3056 8143 3057 8144
rect 3058 8143 3059 8144
rect 3062 8143 3063 8144
rect 3064 8143 3065 8144
rect 2925 8145 2926 8146
rect 3065 8145 3066 8146
rect 3068 8145 3069 8146
rect 3139 8145 3140 8146
rect 2961 8147 2962 8148
rect 3140 8147 3141 8148
rect 3077 8149 3078 8150
rect 3133 8149 3134 8150
rect 3080 8151 3081 8152
rect 3136 8151 3137 8152
rect 3095 8153 3096 8154
rect 3115 8153 3116 8154
rect 3097 8155 3098 8156
rect 3245 8155 3246 8156
rect 3098 8157 3099 8158
rect 3118 8157 3119 8158
rect 3101 8159 3102 8160
rect 3121 8159 3122 8160
rect 3119 8161 3120 8162
rect 3205 8161 3206 8162
rect 3127 8163 3128 8164
rect 3538 8163 3539 8164
rect 3131 8165 3132 8166
rect 3157 8165 3158 8166
rect 3134 8167 3135 8168
rect 3172 8167 3173 8168
rect 3021 8169 3022 8170
rect 3173 8169 3174 8170
rect 3021 8171 3022 8172
rect 3031 8171 3032 8172
rect 3031 8173 3032 8174
rect 3265 8173 3266 8174
rect 3143 8175 3144 8176
rect 3175 8175 3176 8176
rect 3152 8177 3153 8178
rect 3196 8177 3197 8178
rect 3158 8179 3159 8180
rect 3184 8179 3185 8180
rect 3164 8181 3165 8182
rect 3190 8181 3191 8182
rect 3167 8183 3168 8184
rect 3193 8183 3194 8184
rect 3170 8185 3171 8186
rect 3202 8185 3203 8186
rect 3182 8187 3183 8188
rect 3211 8187 3212 8188
rect 3194 8189 3195 8190
rect 3268 8189 3269 8190
rect 3212 8191 3213 8192
rect 3247 8191 3248 8192
rect 3215 8193 3216 8194
rect 3286 8193 3287 8194
rect 3224 8195 3225 8196
rect 3253 8195 3254 8196
rect 3230 8197 3231 8198
rect 3259 8197 3260 8198
rect 3236 8199 3237 8200
rect 3277 8199 3278 8200
rect 3241 8201 3242 8202
rect 3413 8201 3414 8202
rect 3242 8203 3243 8204
rect 3301 8203 3302 8204
rect 3248 8205 3249 8206
rect 3289 8205 3290 8206
rect 3254 8207 3255 8208
rect 3295 8207 3296 8208
rect 3260 8209 3261 8210
rect 3313 8209 3314 8210
rect 3266 8211 3267 8212
rect 3325 8211 3326 8212
rect 3272 8213 3273 8214
rect 3337 8213 3338 8214
rect 3275 8215 3276 8216
rect 3535 8215 3536 8216
rect 3281 8217 3282 8218
rect 3367 8217 3368 8218
rect 3287 8219 3288 8220
rect 3355 8219 3356 8220
rect 3290 8221 3291 8222
rect 3358 8221 3359 8222
rect 3293 8223 3294 8224
rect 3361 8223 3362 8224
rect 3296 8225 3297 8226
rect 3364 8225 3365 8226
rect 3299 8227 3300 8228
rect 3373 8227 3374 8228
rect 3311 8229 3312 8230
rect 3391 8229 3392 8230
rect 3316 8231 3317 8232
rect 3419 8231 3420 8232
rect 3317 8233 3318 8234
rect 3385 8233 3386 8234
rect 3320 8235 3321 8236
rect 3388 8235 3389 8236
rect 3323 8237 3324 8238
rect 3397 8237 3398 8238
rect 3329 8239 3330 8240
rect 3403 8239 3404 8240
rect 3089 8241 3090 8242
rect 3404 8241 3405 8242
rect 3341 8243 3342 8244
rect 3470 8243 3471 8244
rect 3349 8245 3350 8246
rect 3559 8245 3560 8246
rect 3359 8247 3360 8248
rect 3433 8247 3434 8248
rect 3362 8249 3363 8250
rect 3436 8249 3437 8250
rect 3365 8251 3366 8252
rect 3439 8251 3440 8252
rect 3377 8253 3378 8254
rect 3451 8253 3452 8254
rect 3386 8255 3387 8256
rect 3454 8255 3455 8256
rect 3389 8257 3390 8258
rect 3457 8257 3458 8258
rect 3343 8259 3344 8260
rect 3458 8259 3459 8260
rect 3392 8261 3393 8262
rect 3466 8261 3467 8262
rect 3331 8263 3332 8264
rect 3467 8263 3468 8264
rect 3398 8265 3399 8266
rect 3472 8265 3473 8266
rect 3401 8267 3402 8268
rect 3475 8267 3476 8268
rect 3410 8269 3411 8270
rect 3460 8269 3461 8270
rect 3415 8271 3416 8272
rect 3522 8271 3523 8272
rect 3422 8273 3423 8274
rect 3532 8273 3533 8274
rect 3425 8275 3426 8276
rect 3499 8275 3500 8276
rect 3428 8277 3429 8278
rect 3555 8277 3556 8278
rect 3437 8279 3438 8280
rect 3514 8279 3515 8280
rect 3440 8281 3441 8282
rect 3502 8281 3503 8282
rect 3449 8283 3450 8284
rect 3478 8283 3479 8284
rect 3452 8285 3453 8286
rect 3481 8285 3482 8286
rect 3455 8287 3456 8288
rect 3481 8287 3482 8288
rect 3461 8289 3462 8290
rect 3515 8289 3516 8290
rect 3463 8291 3464 8292
rect 3531 8291 3532 8292
rect 3464 8293 3465 8294
rect 3520 8293 3521 8294
rect 3474 8295 3475 8296
rect 3529 8295 3530 8296
rect 3490 8297 3491 8298
rect 3635 8297 3636 8298
rect 3493 8299 3494 8300
rect 3552 8299 3553 8300
rect 3494 8301 3495 8302
rect 3575 8301 3576 8302
rect 3506 8303 3507 8304
rect 3587 8303 3588 8304
rect 3509 8305 3510 8306
rect 3590 8305 3591 8306
rect 3517 8307 3518 8308
rect 3603 8307 3604 8308
rect 3525 8309 3526 8310
rect 3569 8309 3570 8310
rect 3528 8311 3529 8312
rect 3572 8311 3573 8312
rect 3642 8311 3643 8312
rect 3649 8311 3650 8312
rect 3645 8313 3646 8314
rect 3659 8313 3660 8314
rect 2821 8322 2822 8323
rect 2975 8322 2976 8323
rect 2917 8324 2918 8325
rect 3021 8324 3022 8325
rect 2917 8326 2918 8327
rect 3170 8326 3171 8327
rect 2924 8328 2925 8329
rect 3065 8328 3066 8329
rect 2927 8330 2928 8331
rect 3017 8330 3018 8331
rect 2931 8332 2932 8333
rect 3167 8332 3168 8333
rect 2934 8334 2935 8335
rect 3086 8334 3087 8335
rect 2953 8336 2954 8337
rect 3074 8336 3075 8337
rect 2953 8338 2954 8339
rect 3140 8338 3141 8339
rect 2969 8340 2970 8341
rect 3131 8340 3132 8341
rect 2972 8342 2973 8343
rect 2976 8342 2977 8343
rect 2979 8342 2980 8343
rect 3098 8342 3099 8343
rect 2981 8344 2982 8345
rect 3056 8344 3057 8345
rect 2988 8346 2989 8347
rect 3062 8346 3063 8347
rect 2991 8348 2992 8349
rect 3098 8348 3099 8349
rect 2997 8350 2998 8351
rect 3077 8350 3078 8351
rect 2950 8352 2951 8353
rect 3077 8352 3078 8353
rect 2950 8354 2951 8355
rect 3074 8354 3075 8355
rect 3003 8356 3004 8357
rect 3053 8356 3054 8357
rect 3002 8358 3003 8359
rect 3413 8358 3414 8359
rect 3005 8360 3006 8361
rect 3245 8360 3246 8361
rect 3008 8362 3009 8363
rect 3101 8362 3102 8363
rect 3014 8364 3015 8365
rect 3095 8364 3096 8365
rect 3024 8366 3025 8367
rect 3080 8366 3081 8367
rect 3023 8368 3024 8369
rect 3031 8368 3032 8369
rect 3032 8370 3033 8371
rect 3134 8370 3135 8371
rect 3038 8372 3039 8373
rect 3410 8372 3411 8373
rect 2960 8374 2961 8375
rect 3038 8374 3039 8375
rect 3041 8374 3042 8375
rect 3143 8374 3144 8375
rect 3044 8376 3045 8377
rect 3158 8376 3159 8377
rect 3050 8378 3051 8379
rect 3164 8378 3165 8379
rect 3056 8380 3057 8381
rect 3119 8380 3120 8381
rect 3062 8382 3063 8383
rect 3152 8382 3153 8383
rect 3068 8384 3069 8385
rect 3404 8384 3405 8385
rect 3092 8386 3093 8387
rect 3242 8386 3243 8387
rect 3095 8388 3096 8389
rect 3182 8388 3183 8389
rect 3104 8390 3105 8391
rect 3212 8390 3213 8391
rect 3107 8392 3108 8393
rect 3215 8392 3216 8393
rect 3110 8394 3111 8395
rect 3227 8394 3228 8395
rect 3089 8396 3090 8397
rect 3228 8396 3229 8397
rect 3089 8398 3090 8399
rect 3173 8398 3174 8399
rect 3113 8400 3114 8401
rect 3150 8400 3151 8401
rect 3120 8402 3121 8403
rect 3287 8402 3288 8403
rect 3123 8404 3124 8405
rect 3272 8404 3273 8405
rect 3132 8406 3133 8407
rect 3218 8406 3219 8407
rect 3138 8408 3139 8409
rect 3224 8408 3225 8409
rect 3144 8410 3145 8411
rect 3293 8410 3294 8411
rect 3153 8412 3154 8413
rect 3194 8412 3195 8413
rect 3156 8414 3157 8415
rect 3254 8414 3255 8415
rect 3162 8416 3163 8417
rect 3299 8416 3300 8417
rect 3174 8418 3175 8419
rect 3290 8418 3291 8419
rect 3183 8420 3184 8421
rect 3230 8420 3231 8421
rect 3186 8422 3187 8423
rect 3260 8422 3261 8423
rect 3188 8424 3189 8425
rect 3416 8424 3417 8425
rect 3195 8426 3196 8427
rect 3320 8426 3321 8427
rect 3200 8428 3201 8429
rect 3522 8428 3523 8429
rect 3210 8430 3211 8431
rect 3292 8430 3293 8431
rect 3213 8432 3214 8433
rect 3236 8432 3237 8433
rect 3216 8434 3217 8435
rect 3323 8434 3324 8435
rect 3234 8436 3235 8437
rect 3365 8436 3366 8437
rect 3246 8438 3247 8439
rect 3377 8438 3378 8439
rect 3189 8440 3190 8441
rect 3376 8440 3377 8441
rect 3248 8442 3249 8443
rect 3325 8442 3326 8443
rect 3249 8444 3250 8445
rect 3398 8444 3399 8445
rect 3252 8446 3253 8447
rect 3401 8446 3402 8447
rect 3255 8448 3256 8449
rect 3359 8448 3360 8449
rect 3258 8450 3259 8451
rect 3362 8450 3363 8451
rect 3263 8452 3264 8453
rect 3419 8452 3420 8453
rect 3266 8454 3267 8455
rect 3477 8454 3478 8455
rect 3267 8456 3268 8457
rect 3344 8456 3345 8457
rect 3270 8458 3271 8459
rect 3389 8458 3390 8459
rect 3273 8460 3274 8461
rect 3296 8460 3297 8461
rect 3275 8462 3276 8463
rect 3455 8462 3456 8463
rect 3276 8464 3277 8465
rect 3407 8464 3408 8465
rect 3279 8466 3280 8467
rect 3425 8466 3426 8467
rect 3281 8468 3282 8469
rect 3337 8468 3338 8469
rect 3177 8470 3178 8471
rect 3282 8470 3283 8471
rect 3295 8470 3296 8471
rect 3422 8470 3423 8471
rect 3304 8472 3305 8473
rect 3437 8472 3438 8473
rect 3307 8474 3308 8475
rect 3440 8474 3441 8475
rect 3311 8476 3312 8477
rect 3319 8476 3320 8477
rect 3317 8478 3318 8479
rect 3474 8478 3475 8479
rect 3316 8480 3317 8481
rect 3449 8480 3450 8481
rect 3329 8482 3330 8483
rect 3481 8482 3482 8483
rect 3328 8484 3329 8485
rect 3461 8484 3462 8485
rect 3331 8486 3332 8487
rect 3464 8486 3465 8487
rect 3341 8488 3342 8489
rect 3383 8488 3384 8489
rect 3358 8490 3359 8491
rect 3515 8490 3516 8491
rect 3367 8492 3368 8493
rect 3506 8492 3507 8493
rect 3370 8494 3371 8495
rect 3509 8494 3510 8495
rect 3386 8496 3387 8497
rect 3491 8496 3492 8497
rect 3386 8498 3387 8499
rect 3525 8498 3526 8499
rect 3392 8500 3393 8501
rect 3559 8500 3560 8501
rect 3406 8502 3407 8503
rect 3528 8502 3529 8503
rect 3417 8504 3418 8505
rect 3494 8504 3495 8505
rect 3428 8506 3429 8507
rect 3562 8506 3563 8507
rect 3452 8508 3453 8509
rect 3470 8508 3471 8509
rect 3548 8508 3549 8509
rect 3552 8508 3553 8509
rect 2815 8517 2816 8518
rect 2821 8517 2822 8518
rect 2881 8517 2882 8518
rect 2891 8517 2892 8518
rect 2917 8517 2918 8518
rect 3123 8517 3124 8518
rect 2920 8519 2921 8520
rect 3041 8519 3042 8520
rect 2933 8521 2934 8522
rect 3142 8521 3143 8522
rect 2941 8523 2942 8524
rect 3107 8523 3108 8524
rect 2945 8525 2946 8526
rect 3174 8525 3175 8526
rect 2952 8527 2953 8528
rect 3074 8527 3075 8528
rect 2960 8529 2961 8530
rect 3032 8529 3033 8530
rect 2962 8531 2963 8532
rect 3077 8531 3078 8532
rect 2968 8533 2969 8534
rect 3092 8533 3093 8534
rect 2972 8535 2973 8536
rect 2993 8535 2994 8536
rect 2991 8537 2992 8538
rect 3053 8537 3054 8538
rect 2990 8539 2991 8540
rect 3014 8539 3015 8540
rect 2995 8541 2996 8542
rect 3089 8541 3090 8542
rect 3002 8543 3003 8544
rect 3017 8543 3018 8544
rect 2931 8545 2932 8546
rect 3017 8545 3018 8546
rect 3005 8547 3006 8548
rect 3153 8547 3154 8548
rect 3005 8549 3006 8550
rect 3038 8549 3039 8550
rect 3008 8551 3009 8552
rect 3023 8551 3024 8552
rect 3008 8553 3009 8554
rect 3044 8553 3045 8554
rect 2998 8555 2999 8556
rect 3044 8555 3045 8556
rect 2924 8557 2925 8558
rect 2999 8557 3000 8558
rect 3014 8557 3015 8558
rect 3050 8557 3051 8558
rect 3026 8559 3027 8560
rect 3056 8559 3057 8560
rect 3032 8561 3033 8562
rect 3062 8561 3063 8562
rect 3038 8563 3039 8564
rect 3095 8563 3096 8564
rect 3041 8565 3042 8566
rect 3086 8565 3087 8566
rect 3053 8567 3054 8568
rect 3104 8567 3105 8568
rect 3056 8569 3057 8570
rect 3098 8569 3099 8570
rect 3059 8571 3060 8572
rect 3132 8571 3133 8572
rect 3062 8573 3063 8574
rect 3183 8573 3184 8574
rect 3065 8575 3066 8576
rect 3138 8575 3139 8576
rect 3068 8577 3069 8578
rect 3270 8577 3271 8578
rect 3071 8579 3072 8580
rect 3252 8579 3253 8580
rect 3074 8581 3075 8582
rect 3144 8581 3145 8582
rect 3080 8583 3081 8584
rect 3348 8583 3349 8584
rect 3086 8585 3087 8586
rect 3156 8585 3157 8586
rect 3092 8587 3093 8588
rect 3162 8587 3163 8588
rect 3101 8589 3102 8590
rect 3334 8589 3335 8590
rect 3104 8591 3105 8592
rect 3292 8591 3293 8592
rect 3107 8593 3108 8594
rect 3186 8593 3187 8594
rect 3117 8595 3118 8596
rect 3125 8595 3126 8596
rect 3116 8597 3117 8598
rect 3276 8597 3277 8598
rect 3119 8599 3120 8600
rect 3189 8599 3190 8600
rect 3122 8601 3123 8602
rect 3341 8601 3342 8602
rect 3128 8603 3129 8604
rect 3150 8603 3151 8604
rect 3132 8605 3133 8606
rect 3177 8605 3178 8606
rect 3145 8607 3146 8608
rect 3258 8607 3259 8608
rect 3151 8609 3152 8610
rect 3319 8609 3320 8610
rect 3161 8611 3162 8612
rect 3267 8611 3268 8612
rect 3167 8613 3168 8614
rect 3328 8613 3329 8614
rect 3171 8615 3172 8616
rect 3331 8615 3332 8616
rect 3174 8617 3175 8618
rect 3216 8617 3217 8618
rect 3178 8619 3179 8620
rect 3273 8619 3274 8620
rect 3184 8621 3185 8622
rect 3279 8621 3280 8622
rect 3187 8623 3188 8624
rect 3295 8623 3296 8624
rect 3190 8625 3191 8626
rect 3316 8625 3317 8626
rect 3193 8627 3194 8628
rect 3386 8627 3387 8628
rect 3195 8629 3196 8630
rect 3344 8629 3345 8630
rect 3210 8631 3211 8632
rect 3325 8631 3326 8632
rect 3213 8633 3214 8634
rect 3322 8633 3323 8634
rect 3228 8635 3229 8636
rect 3285 8635 3286 8636
rect 3234 8637 3235 8638
rect 3383 8637 3384 8638
rect 3246 8639 3247 8640
rect 3399 8639 3400 8640
rect 3249 8641 3250 8642
rect 3380 8641 3381 8642
rect 3255 8643 3256 8644
rect 3376 8643 3377 8644
rect 3304 8645 3305 8646
rect 3389 8645 3390 8646
rect 3307 8647 3308 8648
rect 3413 8647 3414 8648
rect 3367 8649 3368 8650
rect 3420 8649 3421 8650
rect 3370 8651 3371 8652
rect 3417 8651 3418 8652
rect 2884 8660 2885 8661
rect 2891 8660 2892 8661
rect 2881 8662 2882 8663
rect 2891 8662 2892 8663
rect 2882 8664 2883 8665
rect 2888 8664 2889 8665
rect 2923 8664 2924 8665
rect 3002 8664 3003 8665
rect 2930 8666 2931 8667
rect 3014 8666 3015 8667
rect 2933 8668 2934 8669
rect 3008 8668 3009 8669
rect 2942 8670 2943 8671
rect 2999 8670 3000 8671
rect 2949 8672 2950 8673
rect 2962 8672 2963 8673
rect 2956 8674 2957 8675
rect 3038 8674 3039 8675
rect 2959 8676 2960 8677
rect 3005 8676 3006 8677
rect 2965 8678 2966 8679
rect 2990 8678 2991 8679
rect 2968 8680 2969 8681
rect 3000 8680 3001 8681
rect 2972 8682 2973 8683
rect 3044 8682 3045 8683
rect 2981 8684 2982 8685
rect 3056 8684 3057 8685
rect 2993 8686 2994 8687
rect 3041 8686 3042 8687
rect 2984 8688 2985 8689
rect 2993 8688 2994 8689
rect 2984 8690 2985 8691
rect 3026 8690 3027 8691
rect 2996 8692 2997 8693
rect 3032 8692 3033 8693
rect 2987 8694 2988 8695
rect 2997 8694 2998 8695
rect 3003 8694 3004 8695
rect 3015 8694 3016 8695
rect 3006 8696 3007 8697
rect 3074 8696 3075 8697
rect 3017 8698 3018 8699
rect 3142 8698 3143 8699
rect 3018 8700 3019 8701
rect 3128 8700 3129 8701
rect 3030 8702 3031 8703
rect 3051 8702 3052 8703
rect 3042 8704 3043 8705
rect 3119 8704 3120 8705
rect 3045 8706 3046 8707
rect 3080 8706 3081 8707
rect 3053 8708 3054 8709
rect 3071 8708 3072 8709
rect 3055 8710 3056 8711
rect 3086 8710 3087 8711
rect 3059 8712 3060 8713
rect 3065 8712 3066 8713
rect 3058 8714 3059 8715
rect 3107 8714 3108 8715
rect 3092 8716 3093 8717
rect 3139 8716 3140 8717
rect 3101 8718 3102 8719
rect 3167 8718 3168 8719
rect 3104 8720 3105 8721
rect 3125 8720 3126 8721
rect 3116 8722 3117 8723
rect 3158 8722 3159 8723
rect 3122 8724 3123 8725
rect 3164 8724 3165 8725
rect 3145 8726 3146 8727
rect 3171 8726 3172 8727
rect 3161 8728 3162 8729
rect 3187 8728 3188 8729
rect 3184 8730 3185 8731
rect 3206 8730 3207 8731
rect 3193 8732 3194 8733
rect 3199 8732 3200 8733
rect 2875 8741 2876 8742
rect 2888 8741 2889 8742
rect 2882 8743 2883 8744
rect 2891 8743 2892 8744
rect 2917 8743 2918 8744
rect 2924 8743 2925 8744
rect 2962 8743 2963 8744
rect 2965 8743 2966 8744
rect 2968 8743 2969 8744
rect 3006 8743 3007 8744
rect 2971 8745 2972 8746
rect 2981 8745 2982 8746
rect 2975 8747 2976 8748
rect 2984 8747 2985 8748
rect 2987 8747 2988 8748
rect 2993 8747 2994 8748
rect 2997 8747 2998 8748
rect 3003 8747 3004 8748
rect 3012 8747 3013 8748
rect 3030 8747 3031 8748
rect 3015 8749 3016 8750
rect 3027 8749 3028 8750
rect 3018 8751 3019 8752
rect 3055 8751 3056 8752
rect 3042 8753 3043 8754
rect 3051 8753 3052 8754
rect 3045 8755 3046 8756
rect 3048 8755 3049 8756
<< end >>
