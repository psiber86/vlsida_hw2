magic
tech scmos
timestamp 1395743075
<< m1p >>
use CELL  1
transform -1 0 605 0 1 851
box 0 0 6 6
use CELL  2
transform -1 0 504 0 1 1069
box 0 0 6 6
use CELL  3
transform -1 0 556 0 1 604
box 0 0 6 6
use CELL  4
transform -1 0 504 0 1 991
box 0 0 6 6
use CELL  5
transform -1 0 540 0 1 604
box 0 0 6 6
use CELL  6
transform -1 0 655 0 -1 369
box 0 0 6 6
use CELL  7
transform -1 0 518 0 1 273
box 0 0 6 6
use CELL  8
transform -1 0 538 0 1 363
box 0 0 6 6
use CELL  9
transform -1 0 487 0 1 604
box 0 0 6 6
use CELL  10
transform -1 0 654 0 1 851
box 0 0 6 6
use CELL  11
transform -1 0 529 0 1 426
box 0 0 6 6
use CELL  12
transform -1 0 738 0 1 705
box 0 0 6 6
use CELL  13
transform 1 0 502 0 -1 857
box 0 0 6 6
use CELL  14
transform -1 0 513 0 1 310
box 0 0 6 6
use CELL  15
transform -1 0 616 0 1 991
box 0 0 6 6
use CELL  16
transform -1 0 691 0 1 604
box 0 0 6 6
use CELL  17
transform -1 0 529 0 1 991
box 0 0 6 6
use CELL  18
transform 1 0 619 0 -1 778
box 0 0 6 6
use CELL  19
transform -1 0 474 0 1 705
box 0 0 6 6
use CELL  20
transform -1 0 542 0 1 705
box 0 0 6 6
use CELL  21
transform 1 0 499 0 -1 1092
box 0 0 6 6
use CELL  22
transform 1 0 540 0 -1 254
box 0 0 6 6
use CELL  23
transform 1 0 622 0 1 991
box 0 0 6 6
use CELL  24
transform 1 0 580 0 1 772
box 0 0 6 6
use CELL  25
transform -1 0 486 0 -1 369
box 0 0 6 6
use CELL  26
transform -1 0 578 0 1 705
box 0 0 6 6
use CELL  27
transform -1 0 668 0 1 851
box 0 0 6 6
use CELL  28
transform 1 0 481 0 1 851
box 0 0 6 6
use CELL  29
transform -1 0 750 0 -1 610
box 0 0 6 6
use CELL  30
transform -1 0 736 0 1 604
box 0 0 6 6
use CELL  31
transform 1 0 703 0 -1 711
box 0 0 6 6
use CELL  32
transform -1 0 530 0 -1 1075
box 0 0 6 6
use CELL  33
transform -1 0 528 0 1 604
box 0 0 6 6
use CELL  34
transform -1 0 746 0 1 515
box 0 0 6 6
use CELL  35
transform 1 0 684 0 1 363
box 0 0 6 6
use CELL  36
transform -1 0 511 0 1 705
box 0 0 6 6
use CELL  37
transform -1 0 515 0 1 851
box 0 0 6 6
use CELL  38
transform -1 0 494 0 1 851
box 0 0 6 6
use CELL  39
transform -1 0 520 0 1 1086
box 0 0 6 6
use CELL  40
transform -1 0 581 0 1 1038
box 0 0 6 6
use CELL  41
transform 1 0 633 0 1 851
box 0 0 6 6
use CELL  42
transform -1 0 510 0 1 772
box 0 0 6 6
use CELL  43
transform -1 0 487 0 1 772
box 0 0 6 6
use CELL  44
transform -1 0 486 0 1 924
box 0 0 6 6
use CELL  45
transform -1 0 480 0 1 515
box 0 0 6 6
use CELL  46
transform -1 0 494 0 1 772
box 0 0 6 6
use CELL  47
transform -1 0 509 0 1 363
box 0 0 6 6
use CELL  48
transform 1 0 535 0 1 310
box 0 0 6 6
use CELL  49
transform -1 0 690 0 1 924
box 0 0 6 6
use CELL  50
transform -1 0 525 0 1 924
box 0 0 6 6
use CELL  51
transform -1 0 589 0 1 310
box 0 0 6 6
use CELL  52
transform -1 0 670 0 -1 930
box 0 0 6 6
use CELL  53
transform -1 0 739 0 1 515
box 0 0 6 6
use CELL  54
transform -1 0 498 0 1 1086
box 0 0 6 6
use CELL  55
transform -1 0 494 0 1 604
box 0 0 6 6
use CELL  56
transform -1 0 661 0 1 851
box 0 0 6 6
use CELL  57
transform -1 0 539 0 1 1038
box 0 0 6 6
use CELL  58
transform 1 0 576 0 1 273
box 0 0 6 6
use CELL  59
transform -1 0 551 0 1 273
box 0 0 6 6
use CELL  60
transform -1 0 487 0 1 515
box 0 0 6 6
use CELL  61
transform -1 0 562 0 1 248
box 0 0 6 6
use CELL  62
transform 1 0 615 0 1 310
box 0 0 6 6
use CELL  63
transform -1 0 532 0 1 1038
box 0 0 6 6
use CELL  64
transform 1 0 706 0 1 426
box 0 0 6 6
use CELL  65
transform -1 0 547 0 1 604
box 0 0 6 6
use CELL  66
transform 1 0 668 0 1 851
box 0 0 6 6
use CELL  67
transform 1 0 720 0 1 426
box 0 0 6 6
use CELL  68
transform -1 0 649 0 1 924
box 0 0 6 6
use CELL  69
transform -1 0 504 0 -1 711
box 0 0 6 6
use CELL  70
transform -1 0 495 0 1 705
box 0 0 6 6
use CELL  71
transform -1 0 523 0 1 1069
box 0 0 6 6
use CELL  72
transform -1 0 596 0 -1 316
box 0 0 6 6
use CELL  73
transform -1 0 517 0 1 772
box 0 0 6 6
use CELL  74
transform 1 0 514 0 1 426
box 0 0 6 6
use CELL  75
transform -1 0 764 0 1 604
box 0 0 6 6
use CELL  76
transform -1 0 516 0 1 1069
box 0 0 6 6
use CELL  77
transform -1 0 705 0 1 426
box 0 0 6 6
use CELL  78
transform -1 0 701 0 1 515
box 0 0 6 6
use CELL  79
transform -1 0 506 0 -1 930
box 0 0 6 6
use CELL  80
transform -1 0 611 0 1 705
box 0 0 6 6
use CELL  81
transform -1 0 607 0 1 426
box 0 0 6 6
use CELL  82
transform -1 0 587 0 1 705
box 0 0 6 6
use CELL  83
transform -1 0 500 0 1 363
box 0 0 6 6
use CELL  84
transform -1 0 557 0 1 1038
box 0 0 6 6
use CELL  85
transform -1 0 498 0 1 1038
box 0 0 6 6
use CELL  86
transform -1 0 533 0 1 705
box 0 0 6 6
use CELL  87
transform -1 0 488 0 1 705
box 0 0 6 6
use CELL  88
transform -1 0 492 0 1 991
box 0 0 6 6
use CELL  89
transform -1 0 642 0 1 924
box 0 0 6 6
use CELL  90
transform -1 0 510 0 1 248
box 0 0 6 6
use CELL  91
transform -1 0 731 0 -1 711
box 0 0 6 6
use CELL  92
transform -1 0 676 0 1 924
box 0 0 6 6
use CELL  93
transform -1 0 480 0 1 851
box 0 0 6 6
use CELL  94
transform 1 0 747 0 1 515
box 0 0 6 6
use CELL  95
transform -1 0 649 0 -1 997
box 0 0 6 6
use CELL  96
transform 1 0 622 0 1 310
box 0 0 6 6
use CELL  97
transform -1 0 716 0 1 705
box 0 0 6 6
use CELL  98
transform -1 0 513 0 1 515
box 0 0 6 6
use CELL  99
transform -1 0 480 0 1 604
box 0 0 6 6
use CELL  100
transform -1 0 492 0 -1 316
box 0 0 6 6
use CELL  101
transform -1 0 522 0 1 991
box 0 0 6 6
use CELL  102
transform -1 0 480 0 1 772
box 0 0 6 6
use CELL  103
transform -1 0 531 0 1 363
box 0 0 6 6
use CELL  104
transform -1 0 513 0 1 426
box 0 0 6 6
use CELL  105
transform -1 0 732 0 1 515
box 0 0 6 6
use CELL  106
transform 1 0 629 0 1 310
box 0 0 6 6
use CELL  107
transform -1 0 607 0 1 363
box 0 0 6 6
use CELL  108
transform 1 0 657 0 1 772
box 0 0 6 6
use CELL  109
transform 1 0 656 0 1 363
box 0 0 6 6
use CELL  110
transform -1 0 468 0 1 426
box 0 0 6 6
use CELL  111
transform -1 0 642 0 1 991
box 0 0 6 6
use CELL  112
transform -1 0 553 0 1 248
box 0 0 6 6
use CELL  113
transform -1 0 676 0 1 363
box 0 0 6 6
use CELL  114
transform 1 0 713 0 -1 432
box 0 0 6 6
use CELL  115
transform -1 0 673 0 -1 432
box 0 0 6 6
use CELL  116
transform -1 0 621 0 1 851
box 0 0 6 6
use CELL  117
transform -1 0 695 0 -1 711
box 0 0 6 6
use CELL  118
transform -1 0 757 0 1 604
box 0 0 6 6
use CELL  119
transform -1 0 501 0 1 604
box 0 0 6 6
use CELL  120
transform -1 0 722 0 -1 711
box 0 0 6 6
use CELL  121
transform -1 0 575 0 1 273
box 0 0 6 6
use CELL  122
transform -1 0 493 0 1 924
box 0 0 6 6
use CELL  123
transform -1 0 632 0 1 772
box 0 0 6 6
use CELL  124
transform -1 0 725 0 1 515
box 0 0 6 6
use CELL  125
transform 1 0 583 0 -1 279
box 0 0 6 6
use CELL  126
transform -1 0 499 0 1 310
box 0 0 6 6
use CELL  127
transform -1 0 518 0 -1 711
box 0 0 6 6
use CELL  128
transform -1 0 616 0 -1 778
box 0 0 6 6
use CELL  129
transform -1 0 504 0 1 273
box 0 0 6 6
use CELL  130
transform -1 0 595 0 1 1038
box 0 0 6 6
use CELL  131
transform -1 0 475 0 1 426
box 0 0 6 6
use CELL  132
transform -1 0 511 0 1 273
box 0 0 6 6
use CELL  133
transform -1 0 635 0 1 991
box 0 0 6 6
use CELL  134
transform -1 0 547 0 1 991
box 0 0 6 6
use CELL  135
transform -1 0 567 0 1 924
box 0 0 6 6
use CELL  136
transform -1 0 520 0 1 515
box 0 0 6 6
use CELL  137
transform -1 0 493 0 1 363
box 0 0 6 6
use CELL  138
transform -1 0 499 0 1 924
box 0 0 6 6
use CELL  139
transform -1 0 554 0 1 1069
box 0 0 6 6
use CELL  140
transform -1 0 743 0 1 604
box 0 0 6 6
use CELL  141
transform -1 0 481 0 1 705
box 0 0 6 6
use CELL  142
transform 1 0 536 0 -1 521
box 0 0 6 6
use CELL  143
transform -1 0 505 0 1 1038
box 0 0 6 6
use CELL  144
transform -1 0 503 0 1 772
box 0 0 6 6
use CELL  145
transform -1 0 698 0 1 426
box 0 0 6 6
use CELL  146
transform -1 0 501 0 1 515
box 0 0 6 6
use CELL  147
transform 1 0 633 0 1 772
box 0 0 6 6
use CELL  148
transform -1 0 670 0 1 772
box 0 0 6 6
use CELL  149
transform -1 0 684 0 1 772
box 0 0 6 6
use CELL  150
transform -1 0 683 0 1 924
box 0 0 6 6
use CELL  151
transform -1 0 518 0 1 924
box 0 0 6 6
use CELL  152
transform -1 0 677 0 1 772
box 0 0 6 6
use CELL  153
transform -1 0 584 0 1 851
box 0 0 6 6
use CELL  154
transform -1 0 529 0 -1 778
box 0 0 6 6
use CELL  155
transform 1 0 677 0 -1 521
box 0 0 6 6
use CELL  156
transform 1 0 685 0 1 426
box 0 0 6 6
use CELL  157
transform 1 0 608 0 1 310
box 0 0 6 6
use CELL  158
transform -1 0 492 0 1 273
box 0 0 6 6
use CELL  159
transform -1 0 495 0 1 426
box 0 0 6 6
use CELL  160
transform -1 0 494 0 1 515
box 0 0 6 6
use CELL  161
transform 1 0 482 0 -1 432
box 0 0 6 6
use CELL  162
transform -1 0 501 0 1 851
box 0 0 6 6
use CELL  163
transform 1 0 696 0 1 705
box 0 0 6 6
use CELL  164
transform 1 0 677 0 -1 369
box 0 0 6 6
use CELL  165
transform -1 0 506 0 1 310
box 0 0 6 6
use CELL  166
transform -1 0 516 0 1 363
box 0 0 6 6
use CELL  167
transform 1 0 582 0 1 1038
box 0 0 6 6
use CELL  168
transform -1 0 641 0 1 705
box 0 0 6 6
use CELL  169
transform -1 0 671 0 1 515
box 0 0 6 6
use CELL  170
transform -1 0 481 0 1 426
box 0 0 6 6
use CELL  171
transform -1 0 612 0 1 851
box 0 0 6 6
use CELL  172
transform -1 0 721 0 1 604
box 0 0 6 6
use CELL  173
transform -1 0 527 0 1 515
box 0 0 6 6
use CELL  174
transform -1 0 519 0 1 248
box 0 0 6 6
use CELL  175
transform 1 0 551 0 -1 279
box 0 0 6 6
use CELL  176
transform -1 0 527 0 1 1086
box 0 0 6 6
use CELL  177
transform -1 0 669 0 1 363
box 0 0 6 6
use CELL  178
transform -1 0 527 0 -1 857
box 0 0 6 6
use CELL  179
transform -1 0 520 0 1 310
box 0 0 6 6
use CELL  180
transform -1 0 679 0 1 604
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 627 0 1 924
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 630 0 1 924
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 610 0 1 604
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 611 0 1 515
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 661 0 1 426
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 523 0 1 1038
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 513 0 1 991
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 527 0 1 515
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 589 0 1 426
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 577 0 1 363
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 547 0 1 604
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 518 0 1 705
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 577 0 1 772
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 575 0 1 851
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 637 0 1 363
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 568 0 1 310
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 542 0 1 273
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 539 0 1 273
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 664 0 1 426
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 592 0 1 363
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 625 0 1 426
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 578 0 1 515
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 613 0 1 604
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 531 0 1 604
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 533 0 1 515
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 504 0 1 426
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 500 0 1 363
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 510 0 1 604
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 516 0 1 604
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 495 0 1 705
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 494 0 1 772
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 642 0 1 851
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 648 0 1 772
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 677 0 1 705
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 727 0 1 604
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 542 0 1 515
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 583 0 1 363
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 556 0 1 310
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 722 0 1 705
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 537 0 1 924
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 510 0 1 991
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 562 0 1 363
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 550 0 1 310
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 566 0 1 1038
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 542 0 1 1069
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 580 0 1 991
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 600 0 1 924
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 646 0 1 604
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 647 0 1 515
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 655 0 1 426
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 640 0 1 363
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 596 0 1 515
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 658 0 1 426
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 602 0 1 515
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 529 0 1 991
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 546 0 1 924
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 587 0 1 851
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 601 0 1 772
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 543 0 1 924
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 507 0 1 604
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 551 0 1 705
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 604 0 1 604
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 590 0 1 515
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 508 0 1 1086
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 507 0 1 1069
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 589 0 1 991
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 604 0 1 772
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 590 0 1 851
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 588 0 1 924
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 559 0 1 991
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 501 0 1 426
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 530 0 1 515
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 528 0 1 604
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 578 0 1 705
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 616 0 1 604
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 607 0 1 772
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 649 0 1 924
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 721 0 1 604
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 713 0 1 515
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 679 0 1 426
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 671 0 1 515
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 679 0 1 604
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 623 0 1 705
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 683 0 1 705
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 595 0 1 604
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 562 0 1 604
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 568 0 1 604
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 707 0 1 515
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 710 0 1 515
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 568 0 1 772
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 527 0 1 851
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 534 0 1 924
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 533 0 1 705
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 586 0 1 604
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 572 0 1 515
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 592 0 1 604
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 563 0 1 515
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 577 0 1 426
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 560 0 1 851
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 574 0 1 772
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 566 0 1 851
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 558 0 1 924
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 538 0 1 991
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 548 0 1 851
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 538 0 1 772
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 545 0 1 705
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 583 0 1 604
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 554 0 1 515
box 0 0 3 6
use FEEDTHRU  F-109
transform 1 0 520 0 1 426
box 0 0 3 6
use FEEDTHRU  F-110
transform 1 0 522 0 1 363
box 0 0 3 6
use FEEDTHRU  F-111
transform 1 0 535 0 1 772
box 0 0 3 6
use FEEDTHRU  F-112
transform 1 0 511 0 1 1086
box 0 0 3 6
use FEEDTHRU  F-113
transform 1 0 569 0 1 1038
box 0 0 3 6
use FEEDTHRU  F-114
transform 1 0 545 0 1 1069
box 0 0 3 6
use FEEDTHRU  F-115
transform 1 0 527 0 1 1086
box 0 0 3 6
use FEEDTHRU  F-116
transform 1 0 621 0 1 851
box 0 0 3 6
use FEEDTHRU  F-117
transform 1 0 633 0 1 924
box 0 0 3 6
use FEEDTHRU  F-118
transform 1 0 616 0 1 991
box 0 0 3 6
use FEEDTHRU  F-119
transform 1 0 565 0 1 772
box 0 0 3 6
use FEEDTHRU  F-120
transform 1 0 545 0 1 851
box 0 0 3 6
use FEEDTHRU  F-121
transform 1 0 525 0 1 924
box 0 0 3 6
use FEEDTHRU  F-122
transform 1 0 536 0 1 851
box 0 0 3 6
use FEEDTHRU  F-123
transform 1 0 542 0 1 851
box 0 0 3 6
use FEEDTHRU  F-124
transform 1 0 545 0 1 515
box 0 0 3 6
use FEEDTHRU  F-125
transform 1 0 538 0 1 426
box 0 0 3 6
use FEEDTHRU  F-126
transform 1 0 553 0 1 363
box 0 0 3 6
use FEEDTHRU  F-127
transform 1 0 550 0 1 426
box 0 0 3 6
use FEEDTHRU  F-128
transform 1 0 569 0 1 515
box 0 0 3 6
use FEEDTHRU  F-129
transform 1 0 544 0 1 310
box 0 0 3 6
use FEEDTHRU  F-130
transform 1 0 658 0 1 924
box 0 0 3 6
use FEEDTHRU  F-131
transform 1 0 661 0 1 924
box 0 0 3 6
use FEEDTHRU  F-132
transform 1 0 619 0 1 363
box 0 0 3 6
use FEEDTHRU  F-133
transform 1 0 565 0 1 310
box 0 0 3 6
use FEEDTHRU  F-134
transform 1 0 607 0 1 363
box 0 0 3 6
use FEEDTHRU  F-135
transform 1 0 716 0 1 515
box 0 0 3 6
use FEEDTHRU  F-136
transform 1 0 724 0 1 604
box 0 0 3 6
use FEEDTHRU  F-137
transform 1 0 659 0 1 705
box 0 0 3 6
use FEEDTHRU  F-138
transform 1 0 505 0 1 1086
box 0 0 3 6
use FEEDTHRU  F-139
transform 1 0 504 0 1 1069
box 0 0 3 6
use FEEDTHRU  F-140
transform 1 0 520 0 1 1038
box 0 0 3 6
use FEEDTHRU  F-141
transform 1 0 580 0 1 604
box 0 0 3 6
use FEEDTHRU  F-142
transform 1 0 639 0 1 851
box 0 0 3 6
use FEEDTHRU  F-143
transform 1 0 580 0 1 310
box 0 0 3 6
use FEEDTHRU  F-144
transform 1 0 553 0 1 248
box 0 0 3 6
use FEEDTHRU  F-145
transform 1 0 563 0 1 273
box 0 0 3 6
use FEEDTHRU  F-146
transform 1 0 602 0 1 310
box 0 0 3 6
use FEEDTHRU  F-147
transform 1 0 643 0 1 363
box 0 0 3 6
use FEEDTHRU  F-148
transform 1 0 682 0 1 426
box 0 0 3 6
use FEEDTHRU  F-149
transform 1 0 683 0 1 515
box 0 0 3 6
use FEEDTHRU  F-150
transform 1 0 691 0 1 604
box 0 0 3 6
use FEEDTHRU  F-151
transform 1 0 662 0 1 705
box 0 0 3 6
use FEEDTHRU  F-152
transform 1 0 569 0 1 705
box 0 0 3 6
use FEEDTHRU  F-153
transform 1 0 586 0 1 772
box 0 0 3 6
use FEEDTHRU  F-154
transform 1 0 560 0 1 705
box 0 0 3 6
use FEEDTHRU  F-155
transform 1 0 621 0 1 924
box 0 0 3 6
use FEEDTHRU  F-156
transform 1 0 624 0 1 924
box 0 0 3 6
use FEEDTHRU  F-157
transform 1 0 595 0 1 991
box 0 0 3 6
use FEEDTHRU  F-158
transform 1 0 548 0 1 705
box 0 0 3 6
use FEEDTHRU  F-159
transform 1 0 571 0 1 772
box 0 0 3 6
use FEEDTHRU  F-160
transform 1 0 557 0 1 851
box 0 0 3 6
use FEEDTHRU  F-161
transform 1 0 540 0 1 924
box 0 0 3 6
use FEEDTHRU  F-162
transform 1 0 542 0 1 705
box 0 0 3 6
use FEEDTHRU  F-163
transform 1 0 577 0 1 310
box 0 0 3 6
use FEEDTHRU  F-164
transform 1 0 613 0 1 363
box 0 0 3 6
use FEEDTHRU  F-165
transform 1 0 646 0 1 426
box 0 0 3 6
use FEEDTHRU  F-166
transform 1 0 653 0 1 515
box 0 0 3 6
use FEEDTHRU  F-167
transform 1 0 670 0 1 604
box 0 0 3 6
use FEEDTHRU  F-168
transform 1 0 572 0 1 851
box 0 0 3 6
use FEEDTHRU  F-169
transform 1 0 555 0 1 924
box 0 0 3 6
use FEEDTHRU  F-170
transform 1 0 671 0 1 705
box 0 0 3 6
use FEEDTHRU  F-171
transform 1 0 703 0 1 604
box 0 0 3 6
use FEEDTHRU  F-172
transform 1 0 674 0 1 705
box 0 0 3 6
use FEEDTHRU  F-173
transform 1 0 652 0 1 426
box 0 0 3 6
use FEEDTHRU  F-174
transform 1 0 674 0 1 515
box 0 0 3 6
use FEEDTHRU  F-175
transform 1 0 631 0 1 604
box 0 0 3 6
use FEEDTHRU  F-176
transform 1 0 599 0 1 705
box 0 0 3 6
use FEEDTHRU  F-177
transform 1 0 616 0 1 772
box 0 0 3 6
use FEEDTHRU  F-178
transform 1 0 650 0 1 515
box 0 0 3 6
use FEEDTHRU  F-179
transform 1 0 637 0 1 604
box 0 0 3 6
use FEEDTHRU  F-180
transform 1 0 667 0 1 604
box 0 0 3 6
use FEEDTHRU  F-181
transform 1 0 643 0 1 604
box 0 0 3 6
use FEEDTHRU  F-182
transform 1 0 644 0 1 515
box 0 0 3 6
use FEEDTHRU  F-183
transform 1 0 559 0 1 363
box 0 0 3 6
use FEEDTHRU  F-184
transform 1 0 571 0 1 426
box 0 0 3 6
use FEEDTHRU  F-185
transform 1 0 539 0 1 1038
box 0 0 3 6
use FEEDTHRU  F-186
transform 1 0 562 0 1 991
box 0 0 3 6
use FEEDTHRU  F-187
transform 1 0 591 0 1 924
box 0 0 3 6
use FEEDTHRU  F-188
transform 1 0 553 0 1 991
box 0 0 3 6
use FEEDTHRU  F-189
transform 1 0 567 0 1 924
box 0 0 3 6
use FEEDTHRU  F-190
transform 1 0 511 0 1 1038
box 0 0 3 6
use FEEDTHRU  F-191
transform 1 0 535 0 1 991
box 0 0 3 6
use FEEDTHRU  F-192
transform 1 0 517 0 1 1038
box 0 0 3 6
use FEEDTHRU  F-193
transform 1 0 566 0 1 705
box 0 0 3 6
use FEEDTHRU  F-194
transform 1 0 592 0 1 772
box 0 0 3 6
use FEEDTHRU  F-195
transform 1 0 532 0 1 991
box 0 0 3 6
use FEEDTHRU  F-196
transform 1 0 592 0 1 991
box 0 0 3 6
use FEEDTHRU  F-197
transform 1 0 510 0 1 248
box 0 0 3 6
use FEEDTHRU  F-198
transform 1 0 536 0 1 273
box 0 0 3 6
use FEEDTHRU  F-199
transform 1 0 706 0 1 604
box 0 0 3 6
use FEEDTHRU  F-200
transform 1 0 653 0 1 705
box 0 0 3 6
use FEEDTHRU  F-201
transform 1 0 612 0 1 924
box 0 0 3 6
use FEEDTHRU  F-202
transform 1 0 645 0 1 851
box 0 0 3 6
use FEEDTHRU  F-203
transform 1 0 605 0 1 310
box 0 0 3 6
use FEEDTHRU  F-204
transform 1 0 646 0 1 363
box 0 0 3 6
use FEEDTHRU  F-205
transform 1 0 647 0 1 705
box 0 0 3 6
use FEEDTHRU  F-206
transform 1 0 651 0 1 772
box 0 0 3 6
use FEEDTHRU  F-207
transform 1 0 556 0 1 426
box 0 0 3 6
use FEEDTHRU  F-208
transform 1 0 550 0 1 363
box 0 0 3 6
use FEEDTHRU  F-209
transform 1 0 562 0 1 772
box 0 0 3 6
use FEEDTHRU  F-210
transform 1 0 559 0 1 772
box 0 0 3 6
use FEEDTHRU  F-211
transform 1 0 580 0 1 363
box 0 0 3 6
use FEEDTHRU  F-212
transform 1 0 553 0 1 310
box 0 0 3 6
use FEEDTHRU  F-213
transform 1 0 592 0 1 426
box 0 0 3 6
use FEEDTHRU  F-214
transform 1 0 574 0 1 426
box 0 0 3 6
use FEEDTHRU  F-215
transform 1 0 598 0 1 363
box 0 0 3 6
use FEEDTHRU  F-216
transform 1 0 619 0 1 426
box 0 0 3 6
use FEEDTHRU  F-217
transform 1 0 620 0 1 515
box 0 0 3 6
use FEEDTHRU  F-218
transform 1 0 529 0 1 426
box 0 0 3 6
use FEEDTHRU  F-219
transform 1 0 619 0 1 991
box 0 0 3 6
use FEEDTHRU  F-220
transform 1 0 604 0 1 991
box 0 0 3 6
use FEEDTHRU  F-221
transform 1 0 572 0 1 1038
box 0 0 3 6
use FEEDTHRU  F-222
transform 1 0 616 0 1 363
box 0 0 3 6
use FEEDTHRU  F-223
transform 1 0 643 0 1 426
box 0 0 3 6
use FEEDTHRU  F-224
transform 1 0 656 0 1 515
box 0 0 3 6
use FEEDTHRU  F-225
transform 1 0 622 0 1 426
box 0 0 3 6
use FEEDTHRU  F-226
transform 1 0 623 0 1 515
box 0 0 3 6
use FEEDTHRU  F-227
transform 1 0 612 0 1 851
box 0 0 3 6
use FEEDTHRU  F-228
transform 1 0 594 0 1 924
box 0 0 3 6
use FEEDTHRU  F-229
transform 1 0 680 0 1 705
box 0 0 3 6
use FEEDTHRU  F-230
transform 1 0 686 0 1 705
box 0 0 3 6
use FEEDTHRU  F-231
transform 1 0 639 0 1 772
box 0 0 3 6
use FEEDTHRU  F-232
transform 1 0 581 0 1 515
box 0 0 3 6
use FEEDTHRU  F-233
transform 1 0 562 0 1 426
box 0 0 3 6
use FEEDTHRU  F-234
transform 1 0 556 0 1 363
box 0 0 3 6
use FEEDTHRU  F-235
transform 1 0 566 0 1 273
box 0 0 3 6
use FEEDTHRU  F-236
transform 1 0 602 0 1 705
box 0 0 3 6
use FEEDTHRU  F-237
transform 1 0 661 0 1 604
box 0 0 3 6
use FEEDTHRU  F-238
transform 1 0 632 0 1 515
box 0 0 3 6
use FEEDTHRU  F-239
transform 1 0 532 0 1 310
box 0 0 3 6
use FEEDTHRU  F-240
transform 1 0 527 0 1 273
box 0 0 3 6
use FEEDTHRU  F-241
transform 1 0 524 0 1 273
box 0 0 3 6
use FEEDTHRU  F-242
transform 1 0 541 0 1 310
box 0 0 3 6
use FEEDTHRU  F-243
transform 1 0 563 0 1 1038
box 0 0 3 6
use FEEDTHRU  F-244
transform 1 0 593 0 1 851
box 0 0 3 6
use FEEDTHRU  F-245
transform 1 0 530 0 1 1069
box 0 0 3 6
use FEEDTHRU  F-246
transform 1 0 542 0 1 1038
box 0 0 3 6
use FEEDTHRU  F-247
transform 1 0 577 0 1 991
box 0 0 3 6
use FEEDTHRU  F-248
transform 1 0 573 0 1 924
box 0 0 3 6
use FEEDTHRU  F-249
transform 1 0 595 0 1 426
box 0 0 3 6
use FEEDTHRU  F-250
transform 1 0 595 0 1 363
box 0 0 3 6
use FEEDTHRU  F-251
transform 1 0 608 0 1 515
box 0 0 3 6
use FEEDTHRU  F-252
transform 1 0 649 0 1 426
box 0 0 3 6
use FEEDTHRU  F-253
transform 1 0 626 0 1 515
box 0 0 3 6
use FEEDTHRU  F-254
transform 1 0 649 0 1 604
box 0 0 3 6
use FEEDTHRU  F-255
transform 1 0 654 0 1 772
box 0 0 3 6
use FEEDTHRU  F-256
transform 1 0 630 0 1 851
box 0 0 3 6
use FEEDTHRU  F-257
transform 1 0 584 0 1 851
box 0 0 3 6
use FEEDTHRU  F-258
transform 1 0 598 0 1 772
box 0 0 3 6
use FEEDTHRU  F-259
transform 1 0 617 0 1 705
box 0 0 3 6
use FEEDTHRU  F-260
transform 1 0 568 0 1 426
box 0 0 3 6
use FEEDTHRU  F-261
transform 1 0 574 0 1 363
box 0 0 3 6
use FEEDTHRU  F-262
transform 1 0 547 0 1 310
box 0 0 3 6
use FEEDTHRU  F-263
transform 1 0 586 0 1 426
box 0 0 3 6
use FEEDTHRU  F-264
transform 1 0 548 0 1 1038
box 0 0 3 6
use FEEDTHRU  F-265
transform 1 0 583 0 1 991
box 0 0 3 6
use FEEDTHRU  F-266
transform 1 0 579 0 1 924
box 0 0 3 6
use FEEDTHRU  F-267
transform 1 0 596 0 1 851
box 0 0 3 6
use FEEDTHRU  F-268
transform 1 0 626 0 1 705
box 0 0 3 6
use FEEDTHRU  F-269
transform 1 0 682 0 1 604
box 0 0 3 6
<< metal1 >>
rect 505 245 512 246
rect 544 245 552 246
rect 554 245 558 246
rect 490 255 529 256
rect 502 257 506 258
rect 506 259 526 260
rect 511 261 538 262
rect 513 263 541 264
rect 517 265 544 266
rect 509 267 517 268
rect 551 267 574 268
rect 552 269 568 270
rect 554 271 565 272
rect 580 271 585 272
rect 487 280 558 281
rect 487 282 505 283
rect 490 284 555 285
rect 494 286 526 287
rect 501 288 552 289
rect 509 290 538 291
rect 516 292 544 293
rect 499 294 543 295
rect 518 296 541 297
rect 528 298 534 299
rect 539 298 546 299
rect 549 298 582 299
rect 515 300 549 301
rect 564 300 604 301
rect 567 302 571 303
rect 566 304 585 305
rect 569 306 588 307
rect 578 308 592 309
rect 606 308 624 309
rect 491 317 543 318
rect 494 319 534 320
rect 495 321 502 322
rect 488 323 502 324
rect 508 323 552 324
rect 511 325 564 326
rect 511 327 552 328
rect 523 329 682 330
rect 533 331 594 332
rect 536 333 546 334
rect 548 333 576 334
rect 557 335 585 336
rect 497 337 558 338
rect 498 339 561 340
rect 566 339 609 340
rect 569 341 639 342
rect 578 343 615 344
rect 515 345 579 346
rect 514 347 597 348
rect 581 349 668 350
rect 554 351 582 352
rect 504 353 555 354
rect 587 353 621 354
rect 603 355 645 356
rect 599 357 603 358
rect 606 357 648 358
rect 617 359 672 360
rect 641 361 675 362
rect 491 370 494 371
rect 490 372 570 373
rect 501 374 506 375
rect 481 376 503 377
rect 507 376 540 377
rect 476 378 509 379
rect 511 378 588 379
rect 514 380 576 381
rect 511 382 576 383
rect 521 384 524 385
rect 529 384 582 385
rect 473 386 531 387
rect 533 386 666 387
rect 560 388 573 389
rect 563 390 603 391
rect 557 392 564 393
rect 551 394 558 395
rect 551 396 555 397
rect 578 396 591 397
rect 488 398 579 399
rect 593 398 627 399
rect 526 400 594 401
rect 527 402 585 403
rect 605 402 609 403
rect 605 404 663 405
rect 620 406 694 407
rect 599 408 621 409
rect 638 408 654 409
rect 641 410 657 411
rect 644 412 684 413
rect 617 414 645 415
rect 647 414 715 415
rect 614 416 648 417
rect 650 416 697 417
rect 653 418 704 419
rect 659 420 701 421
rect 667 422 681 423
rect 623 424 669 425
rect 466 433 531 434
rect 470 435 547 436
rect 475 437 486 438
rect 483 439 570 440
rect 479 441 483 442
rect 490 441 500 442
rect 493 443 573 444
rect 489 445 574 446
rect 496 447 516 448
rect 502 449 532 450
rect 505 451 535 452
rect 508 453 540 454
rect 511 455 558 456
rect 518 457 576 458
rect 521 459 556 460
rect 522 461 588 462
rect 524 463 544 464
rect 525 465 594 466
rect 528 467 591 468
rect 537 469 597 470
rect 540 471 610 472
rect 551 473 571 474
rect 563 475 583 476
rect 564 477 579 478
rect 579 479 627 480
rect 591 481 701 482
rect 597 483 660 484
rect 612 485 663 486
rect 627 487 651 488
rect 633 489 724 490
rect 651 491 700 492
rect 653 493 676 494
rect 647 495 655 496
rect 648 497 657 498
rect 644 499 658 500
rect 645 501 721 502
rect 665 503 690 504
rect 603 505 667 506
rect 672 505 735 506
rect 680 507 715 508
rect 708 509 745 510
rect 711 511 742 512
rect 717 513 738 514
rect 475 522 509 523
rect 478 524 547 525
rect 496 526 622 527
rect 496 528 583 529
rect 489 530 582 531
rect 511 532 571 533
rect 499 534 512 535
rect 523 534 570 535
rect 528 536 539 537
rect 529 538 532 539
rect 532 540 535 541
rect 535 542 549 543
rect 543 544 667 545
rect 545 546 618 547
rect 555 548 585 549
rect 554 550 613 551
rect 518 552 612 553
rect 482 554 518 555
rect 564 554 594 555
rect 526 556 564 557
rect 573 556 588 557
rect 579 558 615 559
rect 591 560 606 561
rect 597 562 690 563
rect 515 564 597 565
rect 603 564 687 565
rect 624 566 670 567
rect 633 568 663 569
rect 632 570 700 571
rect 638 572 652 573
rect 627 574 651 575
rect 668 576 724 577
rect 672 578 735 579
rect 654 580 672 581
rect 675 580 721 581
rect 678 582 728 583
rect 609 584 678 585
rect 684 584 693 585
rect 683 586 720 587
rect 704 588 760 589
rect 708 590 756 591
rect 707 592 749 593
rect 711 594 738 595
rect 657 596 739 597
rect 714 598 723 599
rect 717 600 726 601
rect 728 600 731 601
rect 680 602 732 603
rect 472 611 509 612
rect 482 613 512 614
rect 483 615 497 616
rect 485 617 533 618
rect 486 619 570 620
rect 492 621 582 622
rect 493 623 564 624
rect 496 625 518 626
rect 499 627 530 628
rect 506 629 594 630
rect 519 631 549 632
rect 499 633 550 634
rect 526 635 597 636
rect 528 637 539 638
rect 531 639 568 640
rect 534 641 588 642
rect 540 643 606 644
rect 542 645 562 646
rect 545 647 571 648
rect 546 649 585 650
rect 551 651 612 652
rect 489 653 553 654
rect 490 655 544 656
rect 579 655 618 656
rect 585 657 645 658
rect 600 659 633 660
rect 603 661 663 662
rect 609 663 669 664
rect 614 665 735 666
rect 618 667 701 668
rect 624 669 681 670
rect 627 671 684 672
rect 638 673 678 674
rect 647 675 687 676
rect 648 677 712 678
rect 650 679 717 680
rect 654 681 708 682
rect 660 683 726 684
rect 663 685 693 686
rect 671 687 698 688
rect 672 689 760 690
rect 675 691 705 692
rect 678 693 729 694
rect 681 695 739 696
rect 684 697 753 698
rect 687 699 756 700
rect 722 701 749 702
rect 723 703 737 704
rect 469 712 480 713
rect 476 714 564 715
rect 486 716 550 717
rect 490 718 544 719
rect 493 720 514 721
rect 506 722 535 723
rect 537 722 553 723
rect 561 722 583 723
rect 478 724 561 725
rect 567 724 594 725
rect 483 726 567 727
rect 570 726 588 727
rect 509 728 570 729
rect 573 728 609 729
rect 499 730 573 731
rect 498 732 537 733
rect 576 732 580 733
rect 505 734 576 735
rect 519 736 579 737
rect 603 736 631 737
rect 540 738 603 739
rect 539 740 547 741
rect 606 740 625 741
rect 581 742 606 743
rect 611 742 664 743
rect 627 744 640 745
rect 640 746 688 747
rect 648 748 653 749
rect 649 750 679 751
rect 654 752 712 753
rect 655 754 680 755
rect 660 756 715 757
rect 665 758 676 759
rect 672 760 676 761
rect 618 762 673 763
rect 600 764 618 765
rect 599 766 637 767
rect 681 766 691 767
rect 684 768 708 769
rect 720 768 734 769
rect 723 770 730 771
rect 475 779 564 780
rect 482 781 547 782
rect 485 783 496 784
rect 475 785 486 786
rect 489 785 537 786
rect 478 787 538 788
rect 492 789 550 790
rect 492 791 540 792
rect 496 793 561 794
rect 498 795 509 796
rect 499 797 544 798
rect 505 799 567 800
rect 515 801 609 802
rect 527 803 588 804
rect 528 805 570 806
rect 558 807 573 808
rect 512 809 574 810
rect 513 811 568 812
rect 561 813 576 814
rect 576 815 579 816
rect 579 817 594 818
rect 522 819 595 820
rect 582 821 618 822
rect 585 823 600 824
rect 588 825 603 826
rect 591 827 606 828
rect 597 829 608 830
rect 610 829 624 830
rect 613 831 620 832
rect 616 833 628 834
rect 622 835 638 836
rect 631 837 656 838
rect 640 839 680 840
rect 640 841 676 842
rect 643 843 650 844
rect 646 845 673 846
rect 652 847 669 848
rect 656 849 664 850
rect 475 858 547 859
rect 481 860 544 861
rect 492 862 550 863
rect 484 864 492 865
rect 496 864 577 865
rect 497 866 511 867
rect 513 866 562 867
rect 513 868 545 869
rect 516 870 586 871
rect 520 872 583 873
rect 526 874 538 875
rect 503 876 539 877
rect 528 878 536 879
rect 541 878 559 879
rect 547 880 589 881
rect 556 882 574 883
rect 559 884 568 885
rect 565 886 595 887
rect 568 888 617 889
rect 574 890 580 891
rect 580 892 598 893
rect 589 894 592 895
rect 592 896 611 897
rect 595 898 614 899
rect 603 900 629 901
rect 613 902 647 903
rect 622 904 635 905
rect 622 906 675 907
rect 631 908 679 909
rect 600 910 632 911
rect 523 912 602 913
rect 640 912 657 913
rect 643 914 653 915
rect 625 916 645 917
rect 650 916 667 917
rect 659 918 673 919
rect 662 920 689 921
rect 665 922 672 923
rect 484 931 527 932
rect 491 933 534 934
rect 494 935 542 936
rect 497 937 502 938
rect 502 939 515 940
rect 511 941 539 942
rect 517 943 632 944
rect 527 945 545 946
rect 530 947 548 948
rect 535 949 546 950
rect 490 951 537 952
rect 539 951 560 952
rect 554 953 569 954
rect 556 955 563 956
rect 560 957 590 958
rect 520 959 591 960
rect 563 961 593 962
rect 565 963 645 964
rect 574 965 579 966
rect 580 965 585 966
rect 581 967 602 968
rect 593 969 641 970
rect 595 971 631 972
rect 596 973 626 974
rect 605 975 641 976
rect 613 977 645 978
rect 617 979 635 980
rect 620 981 634 982
rect 622 983 648 984
rect 628 985 638 986
rect 650 985 682 986
rect 659 987 689 988
rect 662 989 675 990
rect 487 998 534 999
rect 511 1000 543 1001
rect 512 1002 537 1003
rect 517 1004 561 1005
rect 496 1006 519 1007
rect 520 1006 540 1007
rect 500 1008 522 1009
rect 524 1008 531 1009
rect 502 1010 525 1011
rect 503 1012 515 1013
rect 527 1012 538 1013
rect 540 1012 564 1013
rect 543 1014 579 1015
rect 545 1016 553 1017
rect 549 1018 585 1019
rect 567 1020 615 1021
rect 570 1022 580 1023
rect 573 1024 606 1025
rect 581 1026 612 1027
rect 590 1028 627 1029
rect 593 1030 645 1031
rect 564 1032 594 1033
rect 596 1032 631 1033
rect 617 1034 634 1035
rect 620 1036 638 1037
rect 496 1045 513 1046
rect 500 1047 519 1048
rect 505 1049 522 1050
rect 508 1051 522 1052
rect 518 1053 538 1054
rect 524 1055 528 1056
rect 531 1055 544 1056
rect 540 1057 556 1058
rect 543 1059 568 1060
rect 546 1061 571 1062
rect 549 1063 584 1064
rect 552 1065 580 1066
rect 552 1067 565 1068
rect 573 1067 594 1068
rect 493 1076 500 1077
rect 511 1076 544 1077
rect 512 1078 523 1079
rect 514 1080 529 1081
rect 496 1082 516 1083
rect 528 1082 547 1083
rect 531 1084 550 1085
rect 496 1093 507 1094
rect 503 1095 510 1096
rect 512 1095 519 1096
rect 522 1095 529 1096
<< metal2 >>
rect 505 245 506 249
rect 511 245 512 249
rect 544 245 545 249
rect 551 245 552 249
rect 554 245 555 249
rect 557 245 558 249
rect 490 255 491 274
rect 528 255 529 274
rect 502 257 503 274
rect 505 253 506 258
rect 506 259 507 274
rect 525 259 526 274
rect 511 253 512 262
rect 537 261 538 274
rect 513 263 514 274
rect 540 263 541 274
rect 517 253 518 266
rect 543 265 544 274
rect 509 267 510 274
rect 516 267 517 274
rect 551 253 552 268
rect 573 267 574 274
rect 552 269 553 274
rect 567 269 568 274
rect 554 253 555 272
rect 564 271 565 274
rect 580 271 581 274
rect 584 271 585 274
rect 487 278 488 281
rect 557 280 558 311
rect 487 282 488 311
rect 504 282 505 311
rect 490 278 491 285
rect 554 284 555 311
rect 494 286 495 311
rect 525 278 526 287
rect 501 288 502 311
rect 551 288 552 311
rect 509 278 510 291
rect 537 278 538 291
rect 516 278 517 293
rect 543 278 544 293
rect 499 278 500 295
rect 542 294 543 311
rect 518 296 519 311
rect 540 278 541 297
rect 528 278 529 299
rect 533 298 534 311
rect 539 298 540 311
rect 545 298 546 311
rect 549 278 550 299
rect 581 298 582 311
rect 515 300 516 311
rect 548 300 549 311
rect 564 278 565 301
rect 603 300 604 311
rect 567 278 568 303
rect 570 278 571 303
rect 566 304 567 311
rect 584 304 585 311
rect 569 306 570 311
rect 587 306 588 311
rect 578 308 579 311
rect 591 308 592 311
rect 606 308 607 311
rect 623 308 624 311
rect 491 317 492 364
rect 542 315 543 318
rect 494 315 495 320
rect 533 315 534 320
rect 495 321 496 364
rect 501 315 502 322
rect 488 323 489 364
rect 501 323 502 364
rect 508 315 509 324
rect 551 315 552 324
rect 511 315 512 326
rect 563 325 564 364
rect 511 327 512 364
rect 551 327 552 364
rect 523 329 524 364
rect 681 329 682 364
rect 533 331 534 364
rect 593 331 594 364
rect 536 315 537 334
rect 545 315 546 334
rect 548 315 549 334
rect 575 333 576 364
rect 557 315 558 336
rect 584 335 585 364
rect 497 315 498 338
rect 557 337 558 364
rect 498 339 499 364
rect 560 339 561 364
rect 566 315 567 340
rect 608 339 609 364
rect 569 315 570 342
rect 638 341 639 364
rect 578 315 579 344
rect 614 343 615 364
rect 515 315 516 346
rect 578 345 579 364
rect 514 347 515 364
rect 596 347 597 364
rect 581 315 582 350
rect 667 349 668 364
rect 554 315 555 352
rect 581 351 582 364
rect 504 353 505 364
rect 554 353 555 364
rect 587 315 588 354
rect 620 353 621 364
rect 603 315 604 356
rect 644 355 645 364
rect 599 357 600 364
rect 602 357 603 364
rect 606 315 607 358
rect 647 357 648 364
rect 617 359 618 364
rect 671 359 672 364
rect 641 361 642 364
rect 674 361 675 364
rect 491 368 492 371
rect 493 370 494 427
rect 490 372 491 427
rect 569 372 570 427
rect 501 368 502 375
rect 505 374 506 427
rect 481 368 482 377
rect 502 376 503 427
rect 507 368 508 377
rect 539 376 540 427
rect 476 378 477 427
rect 508 378 509 427
rect 511 368 512 379
rect 587 378 588 427
rect 514 368 515 381
rect 575 368 576 381
rect 511 382 512 427
rect 575 382 576 427
rect 521 384 522 427
rect 523 368 524 385
rect 529 368 530 385
rect 581 368 582 385
rect 473 386 474 427
rect 530 386 531 427
rect 533 368 534 387
rect 665 386 666 427
rect 560 368 561 389
rect 572 388 573 427
rect 563 368 564 391
rect 602 390 603 427
rect 557 368 558 393
rect 563 392 564 427
rect 551 368 552 395
rect 557 394 558 427
rect 551 396 552 427
rect 554 368 555 397
rect 578 368 579 397
rect 590 396 591 427
rect 488 368 489 399
rect 578 398 579 427
rect 593 368 594 399
rect 626 398 627 427
rect 526 368 527 401
rect 593 400 594 427
rect 527 402 528 427
rect 584 368 585 403
rect 596 402 597 427
rect 596 368 597 403
rect 605 368 606 403
rect 608 368 609 403
rect 605 404 606 427
rect 662 404 663 427
rect 620 368 621 407
rect 693 406 694 427
rect 599 368 600 409
rect 620 408 621 427
rect 638 368 639 409
rect 653 368 654 409
rect 641 368 642 411
rect 656 410 657 427
rect 644 368 645 413
rect 683 412 684 427
rect 617 368 618 415
rect 644 414 645 427
rect 647 368 648 415
rect 714 414 715 427
rect 614 368 615 417
rect 647 416 648 427
rect 650 416 651 427
rect 696 416 697 427
rect 653 418 654 427
rect 703 418 704 427
rect 659 420 660 427
rect 700 420 701 427
rect 667 368 668 423
rect 680 422 681 427
rect 623 424 624 427
rect 668 424 669 427
rect 466 431 467 434
rect 530 431 531 434
rect 470 431 471 436
rect 546 435 547 516
rect 475 437 476 516
rect 485 437 486 516
rect 483 431 484 440
rect 569 431 570 440
rect 479 431 480 442
rect 482 441 483 516
rect 490 431 491 442
rect 499 441 500 516
rect 493 431 494 444
rect 572 431 573 444
rect 489 445 490 516
rect 573 445 574 516
rect 496 447 497 516
rect 515 431 516 448
rect 502 431 503 450
rect 531 449 532 516
rect 505 431 506 452
rect 534 451 535 516
rect 508 431 509 454
rect 539 431 540 454
rect 511 455 512 516
rect 557 431 558 456
rect 518 457 519 516
rect 575 431 576 458
rect 521 431 522 460
rect 555 459 556 516
rect 522 461 523 516
rect 587 431 588 462
rect 524 431 525 464
rect 543 463 544 516
rect 525 465 526 516
rect 593 431 594 466
rect 528 467 529 516
rect 590 431 591 468
rect 537 469 538 516
rect 596 431 597 470
rect 540 471 541 516
rect 609 471 610 516
rect 551 431 552 474
rect 570 473 571 516
rect 563 431 564 476
rect 582 475 583 516
rect 564 477 565 516
rect 578 431 579 478
rect 579 479 580 516
rect 626 431 627 480
rect 591 481 592 516
rect 700 431 701 482
rect 597 483 598 516
rect 659 431 660 484
rect 612 485 613 516
rect 662 431 663 486
rect 620 431 621 488
rect 621 487 622 516
rect 623 431 624 488
rect 624 487 625 516
rect 627 487 628 516
rect 650 431 651 488
rect 633 489 634 516
rect 723 489 724 516
rect 651 491 652 516
rect 699 491 700 516
rect 653 431 654 494
rect 675 493 676 516
rect 647 431 648 496
rect 654 495 655 516
rect 648 497 649 516
rect 656 431 657 498
rect 644 431 645 500
rect 657 499 658 516
rect 645 501 646 516
rect 720 501 721 516
rect 665 431 666 504
rect 689 431 690 504
rect 603 505 604 516
rect 666 505 667 516
rect 672 505 673 516
rect 734 505 735 516
rect 680 431 681 508
rect 714 507 715 516
rect 683 431 684 510
rect 684 509 685 516
rect 708 509 709 516
rect 744 509 745 516
rect 711 511 712 516
rect 741 511 742 516
rect 717 513 718 516
rect 737 513 738 516
rect 475 522 476 605
rect 508 522 509 605
rect 478 520 479 525
rect 546 520 547 525
rect 485 524 486 605
rect 485 520 486 525
rect 496 520 497 527
rect 621 520 622 527
rect 496 528 497 605
rect 582 520 583 529
rect 489 520 490 531
rect 581 530 582 605
rect 511 520 512 533
rect 570 520 571 533
rect 499 520 500 535
rect 511 534 512 605
rect 523 534 524 605
rect 569 534 570 605
rect 528 520 529 537
rect 538 536 539 605
rect 529 538 530 605
rect 531 520 532 539
rect 532 540 533 605
rect 534 520 535 541
rect 535 542 536 605
rect 548 542 549 605
rect 543 520 544 545
rect 666 520 667 545
rect 545 546 546 605
rect 617 546 618 605
rect 555 520 556 549
rect 584 548 585 605
rect 554 550 555 605
rect 612 520 613 551
rect 518 520 519 553
rect 611 552 612 605
rect 482 554 483 605
rect 517 554 518 605
rect 564 520 565 555
rect 593 554 594 605
rect 526 556 527 605
rect 563 556 564 605
rect 573 520 574 557
rect 587 556 588 605
rect 579 520 580 559
rect 614 558 615 605
rect 591 520 592 561
rect 605 560 606 605
rect 597 520 598 563
rect 689 562 690 605
rect 515 520 516 565
rect 596 564 597 605
rect 603 520 604 565
rect 686 564 687 605
rect 624 520 625 567
rect 669 520 670 567
rect 633 520 634 569
rect 662 568 663 605
rect 632 570 633 605
rect 699 520 700 571
rect 638 572 639 605
rect 651 520 652 573
rect 627 520 628 575
rect 650 574 651 605
rect 644 576 645 605
rect 645 520 646 577
rect 647 576 648 605
rect 648 520 649 577
rect 668 576 669 605
rect 723 520 724 577
rect 672 520 673 579
rect 734 578 735 605
rect 654 520 655 581
rect 671 580 672 605
rect 675 520 676 581
rect 720 520 721 581
rect 678 520 679 583
rect 727 520 728 583
rect 609 520 610 585
rect 677 584 678 605
rect 684 520 685 585
rect 692 584 693 605
rect 683 586 684 605
rect 719 586 720 605
rect 704 588 705 605
rect 759 588 760 605
rect 708 520 709 591
rect 755 590 756 605
rect 707 592 708 605
rect 748 520 749 593
rect 711 520 712 595
rect 737 520 738 595
rect 657 520 658 597
rect 738 596 739 605
rect 714 520 715 599
rect 722 598 723 605
rect 717 520 718 601
rect 725 600 726 605
rect 728 600 729 605
rect 730 520 731 601
rect 680 602 681 605
rect 731 602 732 605
rect 472 611 473 706
rect 508 609 509 612
rect 482 609 483 614
rect 511 609 512 614
rect 483 615 484 706
rect 496 609 497 616
rect 485 609 486 618
rect 532 609 533 618
rect 486 619 487 706
rect 569 609 570 620
rect 492 609 493 622
rect 581 609 582 622
rect 493 623 494 706
rect 563 609 564 624
rect 496 625 497 706
rect 517 609 518 626
rect 499 609 500 628
rect 529 609 530 628
rect 506 629 507 706
rect 593 609 594 630
rect 519 631 520 706
rect 548 609 549 632
rect 499 633 500 706
rect 549 633 550 706
rect 526 609 527 636
rect 596 609 597 636
rect 528 637 529 706
rect 538 609 539 638
rect 531 639 532 706
rect 567 639 568 706
rect 534 641 535 706
rect 587 609 588 642
rect 540 643 541 706
rect 605 609 606 644
rect 542 609 543 646
rect 561 645 562 706
rect 545 609 546 648
rect 570 647 571 706
rect 546 649 547 706
rect 584 609 585 650
rect 551 609 552 652
rect 611 609 612 652
rect 489 609 490 654
rect 552 653 553 706
rect 490 655 491 706
rect 543 655 544 706
rect 579 655 580 706
rect 617 609 618 656
rect 585 657 586 706
rect 644 609 645 658
rect 600 659 601 706
rect 632 609 633 660
rect 603 661 604 706
rect 662 609 663 662
rect 609 663 610 706
rect 668 609 669 664
rect 614 609 615 666
rect 734 609 735 666
rect 618 667 619 706
rect 700 667 701 706
rect 624 669 625 706
rect 680 609 681 670
rect 627 671 628 706
rect 683 609 684 672
rect 638 609 639 674
rect 677 609 678 674
rect 647 609 648 676
rect 686 609 687 676
rect 648 677 649 706
rect 711 677 712 706
rect 650 609 651 680
rect 716 609 717 680
rect 654 681 655 706
rect 707 609 708 682
rect 660 683 661 706
rect 725 609 726 684
rect 663 685 664 706
rect 692 609 693 686
rect 671 609 672 688
rect 697 687 698 706
rect 672 689 673 706
rect 759 609 760 690
rect 675 691 676 706
rect 704 609 705 692
rect 678 693 679 706
rect 728 609 729 694
rect 681 695 682 706
rect 738 609 739 696
rect 684 697 685 706
rect 752 609 753 698
rect 687 699 688 706
rect 755 609 756 700
rect 722 609 723 702
rect 748 609 749 702
rect 723 703 724 706
rect 736 703 737 706
rect 469 710 470 713
rect 479 710 480 713
rect 476 710 477 715
rect 563 714 564 773
rect 486 710 487 717
rect 549 710 550 717
rect 490 710 491 719
rect 543 710 544 719
rect 493 710 494 721
rect 513 710 514 721
rect 495 722 496 773
rect 496 710 497 723
rect 506 710 507 723
rect 534 710 535 723
rect 537 710 538 723
rect 552 710 553 723
rect 561 710 562 723
rect 582 710 583 723
rect 478 724 479 773
rect 560 724 561 773
rect 567 710 568 725
rect 593 724 594 773
rect 483 710 484 727
rect 566 726 567 773
rect 570 710 571 727
rect 587 726 588 773
rect 509 710 510 729
rect 569 728 570 773
rect 573 710 574 729
rect 608 728 609 773
rect 499 710 500 731
rect 572 730 573 773
rect 498 732 499 773
rect 536 732 537 773
rect 576 710 577 733
rect 579 710 580 733
rect 505 734 506 773
rect 575 734 576 773
rect 519 710 520 737
rect 578 736 579 773
rect 603 710 604 737
rect 630 736 631 773
rect 540 710 541 739
rect 602 738 603 773
rect 539 740 540 773
rect 546 710 547 741
rect 606 710 607 741
rect 624 710 625 741
rect 581 742 582 773
rect 605 742 606 773
rect 611 742 612 773
rect 663 710 664 743
rect 627 710 628 745
rect 639 710 640 745
rect 640 746 641 773
rect 687 710 688 747
rect 648 710 649 749
rect 652 748 653 773
rect 649 750 650 773
rect 678 710 679 751
rect 654 710 655 753
rect 711 710 712 753
rect 655 754 656 773
rect 679 754 680 773
rect 660 710 661 757
rect 714 710 715 757
rect 665 758 666 773
rect 675 710 676 759
rect 672 710 673 761
rect 675 760 676 773
rect 618 710 619 763
rect 672 762 673 773
rect 600 710 601 765
rect 617 764 618 773
rect 599 766 600 773
rect 636 710 637 767
rect 681 710 682 767
rect 690 710 691 767
rect 684 710 685 769
rect 707 710 708 769
rect 720 710 721 769
rect 733 710 734 769
rect 723 710 724 771
rect 729 710 730 771
rect 475 777 476 780
rect 563 777 564 780
rect 482 777 483 782
rect 546 781 547 852
rect 485 777 486 784
rect 495 777 496 784
rect 475 785 476 852
rect 485 785 486 852
rect 489 785 490 852
rect 536 777 537 786
rect 478 787 479 852
rect 537 787 538 852
rect 492 777 493 790
rect 549 789 550 852
rect 492 791 493 852
rect 539 777 540 792
rect 496 793 497 852
rect 560 777 561 794
rect 498 777 499 796
rect 508 777 509 796
rect 499 797 500 852
rect 543 797 544 852
rect 505 777 506 800
rect 566 777 567 800
rect 515 777 516 802
rect 608 777 609 802
rect 527 777 528 804
rect 587 777 588 804
rect 528 805 529 852
rect 569 777 570 806
rect 558 807 559 852
rect 572 777 573 808
rect 512 777 513 810
rect 573 809 574 852
rect 513 811 514 852
rect 567 811 568 852
rect 561 813 562 852
rect 575 777 576 814
rect 576 815 577 852
rect 578 777 579 816
rect 579 817 580 852
rect 593 777 594 818
rect 522 819 523 852
rect 594 819 595 852
rect 582 821 583 852
rect 617 777 618 822
rect 585 823 586 852
rect 599 777 600 824
rect 588 825 589 852
rect 602 777 603 826
rect 591 827 592 852
rect 605 777 606 828
rect 597 829 598 852
rect 607 829 608 852
rect 610 829 611 852
rect 623 777 624 830
rect 613 831 614 852
rect 619 831 620 852
rect 616 833 617 852
rect 627 777 628 834
rect 622 835 623 852
rect 637 835 638 852
rect 631 837 632 852
rect 655 777 656 838
rect 640 777 641 840
rect 679 777 680 840
rect 640 841 641 852
rect 675 777 676 842
rect 643 843 644 852
rect 649 777 650 844
rect 646 845 647 852
rect 672 777 673 846
rect 652 777 653 848
rect 668 777 669 848
rect 656 849 657 852
rect 663 849 664 852
rect 475 856 476 859
rect 546 856 547 859
rect 481 860 482 925
rect 543 856 544 861
rect 492 856 493 863
rect 549 856 550 863
rect 484 864 485 925
rect 491 864 492 925
rect 496 856 497 865
rect 576 856 577 865
rect 497 866 498 925
rect 510 856 511 867
rect 513 856 514 867
rect 561 856 562 867
rect 513 868 514 925
rect 544 868 545 925
rect 516 870 517 925
rect 585 856 586 871
rect 520 872 521 925
rect 582 856 583 873
rect 526 874 527 925
rect 537 856 538 875
rect 503 856 504 877
rect 538 876 539 925
rect 528 856 529 879
rect 535 878 536 925
rect 541 878 542 925
rect 558 856 559 879
rect 547 880 548 925
rect 588 856 589 881
rect 556 882 557 925
rect 573 856 574 883
rect 559 884 560 925
rect 567 856 568 885
rect 565 886 566 925
rect 594 856 595 887
rect 568 888 569 925
rect 616 856 617 889
rect 574 890 575 925
rect 579 856 580 891
rect 580 892 581 925
rect 597 856 598 893
rect 589 894 590 925
rect 591 856 592 895
rect 592 896 593 925
rect 610 856 611 897
rect 595 898 596 925
rect 613 856 614 899
rect 603 856 604 901
rect 628 900 629 925
rect 613 902 614 925
rect 646 856 647 903
rect 622 856 623 905
rect 634 904 635 925
rect 622 906 623 925
rect 674 906 675 925
rect 631 856 632 909
rect 678 908 679 925
rect 600 856 601 911
rect 631 910 632 925
rect 523 912 524 925
rect 601 912 602 925
rect 640 856 641 913
rect 656 856 657 913
rect 643 856 644 915
rect 652 856 653 915
rect 625 916 626 925
rect 644 916 645 925
rect 650 916 651 925
rect 666 856 667 917
rect 659 918 660 925
rect 672 856 673 919
rect 662 920 663 925
rect 688 920 689 925
rect 665 922 666 925
rect 671 922 672 925
rect 484 929 485 932
rect 526 929 527 932
rect 491 929 492 934
rect 533 933 534 992
rect 494 929 495 936
rect 541 929 542 936
rect 497 929 498 938
rect 501 929 502 938
rect 502 939 503 992
rect 514 939 515 992
rect 511 941 512 992
rect 538 929 539 942
rect 517 943 518 992
rect 631 929 632 944
rect 527 945 528 992
rect 544 929 545 946
rect 530 947 531 992
rect 547 929 548 948
rect 535 929 536 950
rect 545 949 546 992
rect 490 951 491 992
rect 536 951 537 992
rect 539 951 540 992
rect 559 929 560 952
rect 554 953 555 992
rect 568 929 569 954
rect 556 929 557 956
rect 562 929 563 956
rect 560 957 561 992
rect 589 929 590 958
rect 520 959 521 992
rect 590 959 591 992
rect 563 961 564 992
rect 592 929 593 962
rect 565 929 566 964
rect 644 929 645 964
rect 574 929 575 966
rect 578 965 579 992
rect 580 929 581 966
rect 584 965 585 992
rect 581 967 582 992
rect 601 929 602 968
rect 593 969 594 992
rect 640 929 641 970
rect 595 929 596 972
rect 630 971 631 992
rect 596 973 597 992
rect 625 929 626 974
rect 605 975 606 992
rect 640 975 641 992
rect 613 929 614 978
rect 644 977 645 992
rect 617 979 618 992
rect 634 929 635 980
rect 620 981 621 992
rect 633 981 634 992
rect 622 929 623 984
rect 647 929 648 984
rect 628 929 629 986
rect 637 929 638 986
rect 650 929 651 986
rect 681 929 682 986
rect 659 929 660 988
rect 688 929 689 988
rect 662 929 663 990
rect 674 929 675 990
rect 487 996 488 999
rect 533 996 534 999
rect 511 996 512 1001
rect 542 996 543 1001
rect 512 1002 513 1039
rect 536 996 537 1003
rect 517 996 518 1005
rect 560 996 561 1005
rect 496 1006 497 1039
rect 518 1006 519 1039
rect 520 996 521 1007
rect 539 996 540 1007
rect 500 1008 501 1039
rect 521 1008 522 1039
rect 524 996 525 1009
rect 530 996 531 1009
rect 502 996 503 1011
rect 524 1010 525 1039
rect 503 1012 504 1039
rect 514 996 515 1013
rect 527 996 528 1013
rect 537 1012 538 1039
rect 540 1012 541 1039
rect 563 996 564 1013
rect 543 1014 544 1039
rect 578 996 579 1015
rect 545 996 546 1017
rect 552 1016 553 1039
rect 549 1018 550 1039
rect 584 996 585 1019
rect 554 996 555 1021
rect 555 1020 556 1039
rect 567 1020 568 1039
rect 614 996 615 1021
rect 570 1022 571 1039
rect 579 1022 580 1039
rect 573 1024 574 1039
rect 605 996 606 1025
rect 581 996 582 1027
rect 611 996 612 1027
rect 590 996 591 1029
rect 626 996 627 1029
rect 593 996 594 1031
rect 644 996 645 1031
rect 564 1032 565 1039
rect 593 1032 594 1039
rect 596 996 597 1033
rect 630 996 631 1033
rect 617 996 618 1035
rect 633 996 634 1035
rect 620 996 621 1037
rect 637 996 638 1037
rect 496 1043 497 1046
rect 512 1043 513 1046
rect 500 1043 501 1048
rect 518 1043 519 1048
rect 505 1049 506 1070
rect 521 1043 522 1050
rect 508 1051 509 1070
rect 521 1051 522 1070
rect 518 1053 519 1070
rect 537 1043 538 1054
rect 524 1043 525 1056
rect 527 1043 528 1056
rect 531 1055 532 1070
rect 543 1043 544 1056
rect 540 1043 541 1058
rect 555 1043 556 1058
rect 543 1059 544 1070
rect 567 1043 568 1060
rect 546 1061 547 1070
rect 570 1043 571 1062
rect 549 1043 550 1064
rect 583 1043 584 1064
rect 552 1043 553 1066
rect 579 1043 580 1066
rect 552 1067 553 1070
rect 564 1043 565 1068
rect 573 1043 574 1068
rect 593 1043 594 1068
rect 493 1076 494 1087
rect 499 1074 500 1077
rect 505 1074 506 1077
rect 506 1076 507 1087
rect 508 1074 509 1077
rect 509 1076 510 1087
rect 511 1074 512 1077
rect 543 1074 544 1077
rect 512 1078 513 1087
rect 522 1078 523 1087
rect 514 1074 515 1081
rect 528 1074 529 1081
rect 496 1082 497 1087
rect 515 1082 516 1087
rect 528 1082 529 1087
rect 546 1074 547 1083
rect 531 1074 532 1085
rect 549 1074 550 1085
rect 496 1091 497 1094
rect 506 1091 507 1094
rect 503 1091 504 1096
rect 509 1091 510 1096
rect 512 1091 513 1096
rect 518 1091 519 1096
rect 522 1091 523 1096
rect 528 1091 529 1096
<< via >>
rect 505 245 506 246
rect 511 245 512 246
rect 544 245 545 246
rect 551 245 552 246
rect 554 245 555 246
rect 557 245 558 246
rect 490 255 491 256
rect 528 255 529 256
rect 502 257 503 258
rect 505 257 506 258
rect 506 259 507 260
rect 525 259 526 260
rect 511 261 512 262
rect 537 261 538 262
rect 513 263 514 264
rect 540 263 541 264
rect 517 265 518 266
rect 543 265 544 266
rect 509 267 510 268
rect 516 267 517 268
rect 551 267 552 268
rect 573 267 574 268
rect 552 269 553 270
rect 567 269 568 270
rect 554 271 555 272
rect 564 271 565 272
rect 580 271 581 272
rect 584 271 585 272
rect 487 280 488 281
rect 557 280 558 281
rect 487 282 488 283
rect 504 282 505 283
rect 490 284 491 285
rect 554 284 555 285
rect 494 286 495 287
rect 525 286 526 287
rect 501 288 502 289
rect 551 288 552 289
rect 509 290 510 291
rect 537 290 538 291
rect 516 292 517 293
rect 543 292 544 293
rect 499 294 500 295
rect 542 294 543 295
rect 518 296 519 297
rect 540 296 541 297
rect 528 298 529 299
rect 533 298 534 299
rect 539 298 540 299
rect 545 298 546 299
rect 549 298 550 299
rect 581 298 582 299
rect 515 300 516 301
rect 548 300 549 301
rect 564 300 565 301
rect 603 300 604 301
rect 567 302 568 303
rect 570 302 571 303
rect 566 304 567 305
rect 584 304 585 305
rect 569 306 570 307
rect 587 306 588 307
rect 578 308 579 309
rect 591 308 592 309
rect 606 308 607 309
rect 623 308 624 309
rect 491 317 492 318
rect 542 317 543 318
rect 494 319 495 320
rect 533 319 534 320
rect 495 321 496 322
rect 501 321 502 322
rect 488 323 489 324
rect 501 323 502 324
rect 508 323 509 324
rect 551 323 552 324
rect 511 325 512 326
rect 563 325 564 326
rect 511 327 512 328
rect 551 327 552 328
rect 523 329 524 330
rect 681 329 682 330
rect 533 331 534 332
rect 593 331 594 332
rect 536 333 537 334
rect 545 333 546 334
rect 548 333 549 334
rect 575 333 576 334
rect 557 335 558 336
rect 584 335 585 336
rect 497 337 498 338
rect 557 337 558 338
rect 498 339 499 340
rect 560 339 561 340
rect 566 339 567 340
rect 608 339 609 340
rect 569 341 570 342
rect 638 341 639 342
rect 578 343 579 344
rect 614 343 615 344
rect 515 345 516 346
rect 578 345 579 346
rect 514 347 515 348
rect 596 347 597 348
rect 581 349 582 350
rect 667 349 668 350
rect 554 351 555 352
rect 581 351 582 352
rect 504 353 505 354
rect 554 353 555 354
rect 587 353 588 354
rect 620 353 621 354
rect 603 355 604 356
rect 644 355 645 356
rect 599 357 600 358
rect 602 357 603 358
rect 606 357 607 358
rect 647 357 648 358
rect 617 359 618 360
rect 671 359 672 360
rect 641 361 642 362
rect 674 361 675 362
rect 491 370 492 371
rect 493 370 494 371
rect 490 372 491 373
rect 569 372 570 373
rect 501 374 502 375
rect 505 374 506 375
rect 481 376 482 377
rect 502 376 503 377
rect 507 376 508 377
rect 539 376 540 377
rect 476 378 477 379
rect 508 378 509 379
rect 511 378 512 379
rect 587 378 588 379
rect 514 380 515 381
rect 575 380 576 381
rect 511 382 512 383
rect 575 382 576 383
rect 521 384 522 385
rect 523 384 524 385
rect 529 384 530 385
rect 581 384 582 385
rect 473 386 474 387
rect 530 386 531 387
rect 533 386 534 387
rect 665 386 666 387
rect 560 388 561 389
rect 572 388 573 389
rect 563 390 564 391
rect 602 390 603 391
rect 557 392 558 393
rect 563 392 564 393
rect 551 394 552 395
rect 557 394 558 395
rect 551 396 552 397
rect 554 396 555 397
rect 578 396 579 397
rect 590 396 591 397
rect 488 398 489 399
rect 578 398 579 399
rect 593 398 594 399
rect 626 398 627 399
rect 526 400 527 401
rect 593 400 594 401
rect 527 402 528 403
rect 584 402 585 403
rect 605 402 606 403
rect 608 402 609 403
rect 605 404 606 405
rect 662 404 663 405
rect 620 406 621 407
rect 693 406 694 407
rect 599 408 600 409
rect 620 408 621 409
rect 638 408 639 409
rect 653 408 654 409
rect 641 410 642 411
rect 656 410 657 411
rect 644 412 645 413
rect 683 412 684 413
rect 617 414 618 415
rect 644 414 645 415
rect 647 414 648 415
rect 714 414 715 415
rect 614 416 615 417
rect 647 416 648 417
rect 650 416 651 417
rect 696 416 697 417
rect 653 418 654 419
rect 703 418 704 419
rect 659 420 660 421
rect 700 420 701 421
rect 667 422 668 423
rect 680 422 681 423
rect 623 424 624 425
rect 668 424 669 425
rect 466 433 467 434
rect 530 433 531 434
rect 470 435 471 436
rect 546 435 547 436
rect 475 437 476 438
rect 485 437 486 438
rect 483 439 484 440
rect 569 439 570 440
rect 479 441 480 442
rect 482 441 483 442
rect 490 441 491 442
rect 499 441 500 442
rect 493 443 494 444
rect 572 443 573 444
rect 489 445 490 446
rect 573 445 574 446
rect 496 447 497 448
rect 515 447 516 448
rect 502 449 503 450
rect 531 449 532 450
rect 505 451 506 452
rect 534 451 535 452
rect 508 453 509 454
rect 539 453 540 454
rect 511 455 512 456
rect 557 455 558 456
rect 518 457 519 458
rect 575 457 576 458
rect 521 459 522 460
rect 555 459 556 460
rect 522 461 523 462
rect 587 461 588 462
rect 524 463 525 464
rect 543 463 544 464
rect 525 465 526 466
rect 593 465 594 466
rect 528 467 529 468
rect 590 467 591 468
rect 537 469 538 470
rect 596 469 597 470
rect 540 471 541 472
rect 609 471 610 472
rect 551 473 552 474
rect 570 473 571 474
rect 563 475 564 476
rect 582 475 583 476
rect 564 477 565 478
rect 578 477 579 478
rect 579 479 580 480
rect 626 479 627 480
rect 591 481 592 482
rect 700 481 701 482
rect 597 483 598 484
rect 659 483 660 484
rect 612 485 613 486
rect 662 485 663 486
rect 627 487 628 488
rect 650 487 651 488
rect 633 489 634 490
rect 723 489 724 490
rect 651 491 652 492
rect 699 491 700 492
rect 653 493 654 494
rect 675 493 676 494
rect 647 495 648 496
rect 654 495 655 496
rect 648 497 649 498
rect 656 497 657 498
rect 644 499 645 500
rect 657 499 658 500
rect 645 501 646 502
rect 720 501 721 502
rect 665 503 666 504
rect 689 503 690 504
rect 603 505 604 506
rect 666 505 667 506
rect 672 505 673 506
rect 734 505 735 506
rect 680 507 681 508
rect 714 507 715 508
rect 708 509 709 510
rect 744 509 745 510
rect 711 511 712 512
rect 741 511 742 512
rect 717 513 718 514
rect 737 513 738 514
rect 475 522 476 523
rect 508 522 509 523
rect 478 524 479 525
rect 546 524 547 525
rect 496 526 497 527
rect 621 526 622 527
rect 496 528 497 529
rect 582 528 583 529
rect 489 530 490 531
rect 581 530 582 531
rect 511 532 512 533
rect 570 532 571 533
rect 499 534 500 535
rect 511 534 512 535
rect 523 534 524 535
rect 569 534 570 535
rect 528 536 529 537
rect 538 536 539 537
rect 529 538 530 539
rect 531 538 532 539
rect 532 540 533 541
rect 534 540 535 541
rect 535 542 536 543
rect 548 542 549 543
rect 543 544 544 545
rect 666 544 667 545
rect 545 546 546 547
rect 617 546 618 547
rect 555 548 556 549
rect 584 548 585 549
rect 554 550 555 551
rect 612 550 613 551
rect 518 552 519 553
rect 611 552 612 553
rect 482 554 483 555
rect 517 554 518 555
rect 564 554 565 555
rect 593 554 594 555
rect 526 556 527 557
rect 563 556 564 557
rect 573 556 574 557
rect 587 556 588 557
rect 579 558 580 559
rect 614 558 615 559
rect 591 560 592 561
rect 605 560 606 561
rect 597 562 598 563
rect 689 562 690 563
rect 515 564 516 565
rect 596 564 597 565
rect 603 564 604 565
rect 686 564 687 565
rect 624 566 625 567
rect 669 566 670 567
rect 633 568 634 569
rect 662 568 663 569
rect 632 570 633 571
rect 699 570 700 571
rect 638 572 639 573
rect 651 572 652 573
rect 627 574 628 575
rect 650 574 651 575
rect 668 576 669 577
rect 723 576 724 577
rect 672 578 673 579
rect 734 578 735 579
rect 654 580 655 581
rect 671 580 672 581
rect 675 580 676 581
rect 720 580 721 581
rect 678 582 679 583
rect 727 582 728 583
rect 609 584 610 585
rect 677 584 678 585
rect 684 584 685 585
rect 692 584 693 585
rect 683 586 684 587
rect 719 586 720 587
rect 704 588 705 589
rect 759 588 760 589
rect 708 590 709 591
rect 755 590 756 591
rect 707 592 708 593
rect 748 592 749 593
rect 711 594 712 595
rect 737 594 738 595
rect 657 596 658 597
rect 738 596 739 597
rect 714 598 715 599
rect 722 598 723 599
rect 717 600 718 601
rect 725 600 726 601
rect 728 600 729 601
rect 730 600 731 601
rect 680 602 681 603
rect 731 602 732 603
rect 472 611 473 612
rect 508 611 509 612
rect 482 613 483 614
rect 511 613 512 614
rect 483 615 484 616
rect 496 615 497 616
rect 485 617 486 618
rect 532 617 533 618
rect 486 619 487 620
rect 569 619 570 620
rect 492 621 493 622
rect 581 621 582 622
rect 493 623 494 624
rect 563 623 564 624
rect 496 625 497 626
rect 517 625 518 626
rect 499 627 500 628
rect 529 627 530 628
rect 506 629 507 630
rect 593 629 594 630
rect 519 631 520 632
rect 548 631 549 632
rect 499 633 500 634
rect 549 633 550 634
rect 526 635 527 636
rect 596 635 597 636
rect 528 637 529 638
rect 538 637 539 638
rect 531 639 532 640
rect 567 639 568 640
rect 534 641 535 642
rect 587 641 588 642
rect 540 643 541 644
rect 605 643 606 644
rect 542 645 543 646
rect 561 645 562 646
rect 545 647 546 648
rect 570 647 571 648
rect 546 649 547 650
rect 584 649 585 650
rect 551 651 552 652
rect 611 651 612 652
rect 489 653 490 654
rect 552 653 553 654
rect 490 655 491 656
rect 543 655 544 656
rect 579 655 580 656
rect 617 655 618 656
rect 585 657 586 658
rect 644 657 645 658
rect 600 659 601 660
rect 632 659 633 660
rect 603 661 604 662
rect 662 661 663 662
rect 609 663 610 664
rect 668 663 669 664
rect 614 665 615 666
rect 734 665 735 666
rect 618 667 619 668
rect 700 667 701 668
rect 624 669 625 670
rect 680 669 681 670
rect 627 671 628 672
rect 683 671 684 672
rect 638 673 639 674
rect 677 673 678 674
rect 647 675 648 676
rect 686 675 687 676
rect 648 677 649 678
rect 711 677 712 678
rect 650 679 651 680
rect 716 679 717 680
rect 654 681 655 682
rect 707 681 708 682
rect 660 683 661 684
rect 725 683 726 684
rect 663 685 664 686
rect 692 685 693 686
rect 671 687 672 688
rect 697 687 698 688
rect 672 689 673 690
rect 759 689 760 690
rect 675 691 676 692
rect 704 691 705 692
rect 678 693 679 694
rect 728 693 729 694
rect 681 695 682 696
rect 738 695 739 696
rect 684 697 685 698
rect 752 697 753 698
rect 687 699 688 700
rect 755 699 756 700
rect 722 701 723 702
rect 748 701 749 702
rect 723 703 724 704
rect 736 703 737 704
rect 469 712 470 713
rect 479 712 480 713
rect 476 714 477 715
rect 563 714 564 715
rect 486 716 487 717
rect 549 716 550 717
rect 490 718 491 719
rect 543 718 544 719
rect 493 720 494 721
rect 513 720 514 721
rect 506 722 507 723
rect 534 722 535 723
rect 537 722 538 723
rect 552 722 553 723
rect 561 722 562 723
rect 582 722 583 723
rect 478 724 479 725
rect 560 724 561 725
rect 567 724 568 725
rect 593 724 594 725
rect 483 726 484 727
rect 566 726 567 727
rect 570 726 571 727
rect 587 726 588 727
rect 509 728 510 729
rect 569 728 570 729
rect 573 728 574 729
rect 608 728 609 729
rect 499 730 500 731
rect 572 730 573 731
rect 498 732 499 733
rect 536 732 537 733
rect 576 732 577 733
rect 579 732 580 733
rect 505 734 506 735
rect 575 734 576 735
rect 519 736 520 737
rect 578 736 579 737
rect 603 736 604 737
rect 630 736 631 737
rect 540 738 541 739
rect 602 738 603 739
rect 539 740 540 741
rect 546 740 547 741
rect 606 740 607 741
rect 624 740 625 741
rect 581 742 582 743
rect 605 742 606 743
rect 611 742 612 743
rect 663 742 664 743
rect 627 744 628 745
rect 639 744 640 745
rect 640 746 641 747
rect 687 746 688 747
rect 648 748 649 749
rect 652 748 653 749
rect 649 750 650 751
rect 678 750 679 751
rect 654 752 655 753
rect 711 752 712 753
rect 655 754 656 755
rect 679 754 680 755
rect 660 756 661 757
rect 714 756 715 757
rect 665 758 666 759
rect 675 758 676 759
rect 672 760 673 761
rect 675 760 676 761
rect 618 762 619 763
rect 672 762 673 763
rect 600 764 601 765
rect 617 764 618 765
rect 599 766 600 767
rect 636 766 637 767
rect 681 766 682 767
rect 690 766 691 767
rect 684 768 685 769
rect 707 768 708 769
rect 720 768 721 769
rect 733 768 734 769
rect 723 770 724 771
rect 729 770 730 771
rect 475 779 476 780
rect 563 779 564 780
rect 482 781 483 782
rect 546 781 547 782
rect 485 783 486 784
rect 495 783 496 784
rect 475 785 476 786
rect 485 785 486 786
rect 489 785 490 786
rect 536 785 537 786
rect 478 787 479 788
rect 537 787 538 788
rect 492 789 493 790
rect 549 789 550 790
rect 492 791 493 792
rect 539 791 540 792
rect 496 793 497 794
rect 560 793 561 794
rect 498 795 499 796
rect 508 795 509 796
rect 499 797 500 798
rect 543 797 544 798
rect 505 799 506 800
rect 566 799 567 800
rect 515 801 516 802
rect 608 801 609 802
rect 527 803 528 804
rect 587 803 588 804
rect 528 805 529 806
rect 569 805 570 806
rect 558 807 559 808
rect 572 807 573 808
rect 512 809 513 810
rect 573 809 574 810
rect 513 811 514 812
rect 567 811 568 812
rect 561 813 562 814
rect 575 813 576 814
rect 576 815 577 816
rect 578 815 579 816
rect 579 817 580 818
rect 593 817 594 818
rect 522 819 523 820
rect 594 819 595 820
rect 582 821 583 822
rect 617 821 618 822
rect 585 823 586 824
rect 599 823 600 824
rect 588 825 589 826
rect 602 825 603 826
rect 591 827 592 828
rect 605 827 606 828
rect 597 829 598 830
rect 607 829 608 830
rect 610 829 611 830
rect 623 829 624 830
rect 613 831 614 832
rect 619 831 620 832
rect 616 833 617 834
rect 627 833 628 834
rect 622 835 623 836
rect 637 835 638 836
rect 631 837 632 838
rect 655 837 656 838
rect 640 839 641 840
rect 679 839 680 840
rect 640 841 641 842
rect 675 841 676 842
rect 643 843 644 844
rect 649 843 650 844
rect 646 845 647 846
rect 672 845 673 846
rect 652 847 653 848
rect 668 847 669 848
rect 656 849 657 850
rect 663 849 664 850
rect 475 858 476 859
rect 546 858 547 859
rect 481 860 482 861
rect 543 860 544 861
rect 492 862 493 863
rect 549 862 550 863
rect 484 864 485 865
rect 491 864 492 865
rect 496 864 497 865
rect 576 864 577 865
rect 497 866 498 867
rect 510 866 511 867
rect 513 866 514 867
rect 561 866 562 867
rect 513 868 514 869
rect 544 868 545 869
rect 516 870 517 871
rect 585 870 586 871
rect 520 872 521 873
rect 582 872 583 873
rect 526 874 527 875
rect 537 874 538 875
rect 503 876 504 877
rect 538 876 539 877
rect 528 878 529 879
rect 535 878 536 879
rect 541 878 542 879
rect 558 878 559 879
rect 547 880 548 881
rect 588 880 589 881
rect 556 882 557 883
rect 573 882 574 883
rect 559 884 560 885
rect 567 884 568 885
rect 565 886 566 887
rect 594 886 595 887
rect 568 888 569 889
rect 616 888 617 889
rect 574 890 575 891
rect 579 890 580 891
rect 580 892 581 893
rect 597 892 598 893
rect 589 894 590 895
rect 591 894 592 895
rect 592 896 593 897
rect 610 896 611 897
rect 595 898 596 899
rect 613 898 614 899
rect 603 900 604 901
rect 628 900 629 901
rect 613 902 614 903
rect 646 902 647 903
rect 622 904 623 905
rect 634 904 635 905
rect 622 906 623 907
rect 674 906 675 907
rect 631 908 632 909
rect 678 908 679 909
rect 600 910 601 911
rect 631 910 632 911
rect 523 912 524 913
rect 601 912 602 913
rect 640 912 641 913
rect 656 912 657 913
rect 643 914 644 915
rect 652 914 653 915
rect 625 916 626 917
rect 644 916 645 917
rect 650 916 651 917
rect 666 916 667 917
rect 659 918 660 919
rect 672 918 673 919
rect 662 920 663 921
rect 688 920 689 921
rect 665 922 666 923
rect 671 922 672 923
rect 484 931 485 932
rect 526 931 527 932
rect 491 933 492 934
rect 533 933 534 934
rect 494 935 495 936
rect 541 935 542 936
rect 497 937 498 938
rect 501 937 502 938
rect 502 939 503 940
rect 514 939 515 940
rect 511 941 512 942
rect 538 941 539 942
rect 517 943 518 944
rect 631 943 632 944
rect 527 945 528 946
rect 544 945 545 946
rect 530 947 531 948
rect 547 947 548 948
rect 535 949 536 950
rect 545 949 546 950
rect 490 951 491 952
rect 536 951 537 952
rect 539 951 540 952
rect 559 951 560 952
rect 554 953 555 954
rect 568 953 569 954
rect 556 955 557 956
rect 562 955 563 956
rect 560 957 561 958
rect 589 957 590 958
rect 520 959 521 960
rect 590 959 591 960
rect 563 961 564 962
rect 592 961 593 962
rect 565 963 566 964
rect 644 963 645 964
rect 574 965 575 966
rect 578 965 579 966
rect 580 965 581 966
rect 584 965 585 966
rect 581 967 582 968
rect 601 967 602 968
rect 593 969 594 970
rect 640 969 641 970
rect 595 971 596 972
rect 630 971 631 972
rect 596 973 597 974
rect 625 973 626 974
rect 605 975 606 976
rect 640 975 641 976
rect 613 977 614 978
rect 644 977 645 978
rect 617 979 618 980
rect 634 979 635 980
rect 620 981 621 982
rect 633 981 634 982
rect 622 983 623 984
rect 647 983 648 984
rect 628 985 629 986
rect 637 985 638 986
rect 650 985 651 986
rect 681 985 682 986
rect 659 987 660 988
rect 688 987 689 988
rect 662 989 663 990
rect 674 989 675 990
rect 487 998 488 999
rect 533 998 534 999
rect 511 1000 512 1001
rect 542 1000 543 1001
rect 512 1002 513 1003
rect 536 1002 537 1003
rect 517 1004 518 1005
rect 560 1004 561 1005
rect 496 1006 497 1007
rect 518 1006 519 1007
rect 520 1006 521 1007
rect 539 1006 540 1007
rect 500 1008 501 1009
rect 521 1008 522 1009
rect 524 1008 525 1009
rect 530 1008 531 1009
rect 502 1010 503 1011
rect 524 1010 525 1011
rect 503 1012 504 1013
rect 514 1012 515 1013
rect 527 1012 528 1013
rect 537 1012 538 1013
rect 540 1012 541 1013
rect 563 1012 564 1013
rect 543 1014 544 1015
rect 578 1014 579 1015
rect 545 1016 546 1017
rect 552 1016 553 1017
rect 549 1018 550 1019
rect 584 1018 585 1019
rect 567 1020 568 1021
rect 614 1020 615 1021
rect 570 1022 571 1023
rect 579 1022 580 1023
rect 573 1024 574 1025
rect 605 1024 606 1025
rect 581 1026 582 1027
rect 611 1026 612 1027
rect 590 1028 591 1029
rect 626 1028 627 1029
rect 593 1030 594 1031
rect 644 1030 645 1031
rect 564 1032 565 1033
rect 593 1032 594 1033
rect 596 1032 597 1033
rect 630 1032 631 1033
rect 617 1034 618 1035
rect 633 1034 634 1035
rect 620 1036 621 1037
rect 637 1036 638 1037
rect 496 1045 497 1046
rect 512 1045 513 1046
rect 500 1047 501 1048
rect 518 1047 519 1048
rect 505 1049 506 1050
rect 521 1049 522 1050
rect 508 1051 509 1052
rect 521 1051 522 1052
rect 518 1053 519 1054
rect 537 1053 538 1054
rect 524 1055 525 1056
rect 527 1055 528 1056
rect 531 1055 532 1056
rect 543 1055 544 1056
rect 540 1057 541 1058
rect 555 1057 556 1058
rect 543 1059 544 1060
rect 567 1059 568 1060
rect 546 1061 547 1062
rect 570 1061 571 1062
rect 549 1063 550 1064
rect 583 1063 584 1064
rect 552 1065 553 1066
rect 579 1065 580 1066
rect 552 1067 553 1068
rect 564 1067 565 1068
rect 573 1067 574 1068
rect 593 1067 594 1068
rect 493 1076 494 1077
rect 499 1076 500 1077
rect 511 1076 512 1077
rect 543 1076 544 1077
rect 512 1078 513 1079
rect 522 1078 523 1079
rect 514 1080 515 1081
rect 528 1080 529 1081
rect 496 1082 497 1083
rect 515 1082 516 1083
rect 528 1082 529 1083
rect 546 1082 547 1083
rect 531 1084 532 1085
rect 549 1084 550 1085
rect 496 1093 497 1094
rect 506 1093 507 1094
rect 503 1095 504 1096
rect 509 1095 510 1096
rect 512 1095 513 1096
rect 518 1095 519 1096
rect 522 1095 523 1096
rect 528 1095 529 1096
<< end >>
