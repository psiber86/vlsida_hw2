magic
tech scmos
timestamp 1395741038
<< m1p >>
use CELL  1
transform -1 0 2912 0 1 1485
box 0 0 6 6
use CELL  2
transform 1 0 2924 0 1 1485
box 0 0 6 6
use CELL  3
transform -1 0 2912 0 1 1530
box 0 0 6 6
use CELL  4
transform -1 0 2949 0 1 1512
box 0 0 6 6
use CELL  5
transform -1 0 3198 0 1 1548
box 0 0 6 6
use CELL  6
transform -1 0 2923 0 1 1422
box 0 0 6 6
use CELL  7
transform 1 0 3797 0 -1 1554
box 0 0 6 6
use CELL  8
transform 1 0 3551 0 1 1440
box 0 0 6 6
use CELL  9
transform -1 0 3168 0 1 1548
box 0 0 6 6
use CELL  10
transform -1 0 3677 0 1 1647
box 0 0 6 6
use CELL  11
transform -1 0 3042 0 1 1620
box 0 0 6 6
use CELL  12
transform -1 0 3139 0 1 1629
box 0 0 6 6
use CELL  13
transform -1 0 3698 0 1 1602
box 0 0 6 6
use CELL  14
transform 1 0 3099 0 -1 1689
box 0 0 6 6
use CELL  15
transform -1 0 3799 0 1 1476
box 0 0 6 6
use CELL  16
transform 1 0 3800 0 1 1476
box 0 0 6 6
use CELL  17
transform -1 0 2911 0 1 1602
box 0 0 6 6
use CELL  18
transform -1 0 3654 0 1 1638
box 0 0 6 6
use CELL  19
transform -1 0 3703 0 1 1629
box 0 0 6 6
use CELL  20
transform -1 0 2913 0 1 1566
box 0 0 6 6
use CELL  21
transform -1 0 3144 0 1 1422
box 0 0 6 6
use CELL  22
transform -1 0 2944 0 1 1638
box 0 0 6 6
use CELL  23
transform 1 0 3471 0 -1 1437
box 0 0 6 6
use CELL  24
transform -1 0 3092 0 1 1467
box 0 0 6 6
use CELL  25
transform -1 0 2952 0 1 1539
box 0 0 6 6
use CELL  26
transform 1 0 3755 0 -1 1617
box 0 0 6 6
use CELL  27
transform -1 0 3564 0 1 1656
box 0 0 6 6
use CELL  28
transform -1 0 3675 0 1 1638
box 0 0 6 6
use CELL  29
transform -1 0 3892 0 1 1530
box 0 0 6 6
use CELL  30
transform -1 0 3806 0 1 1557
box 0 0 6 6
use CELL  31
transform -1 0 3021 0 1 1521
box 0 0 6 6
use CELL  32
transform -1 0 2948 0 1 1665
box 0 0 6 6
use CELL  33
transform -1 0 3424 0 1 1665
box 0 0 6 6
use CELL  34
transform -1 0 3105 0 1 1422
box 0 0 6 6
use CELL  35
transform -1 0 3313 0 1 1674
box 0 0 6 6
use CELL  36
transform -1 0 3834 0 1 1557
box 0 0 6 6
use CELL  37
transform -1 0 2906 0 1 1494
box 0 0 6 6
use CELL  38
transform -1 0 2951 0 1 1575
box 0 0 6 6
use CELL  39
transform -1 0 3848 0 1 1467
box 0 0 6 6
use CELL  40
transform -1 0 2944 0 1 1647
box 0 0 6 6
use CELL  41
transform -1 0 2911 0 1 1476
box 0 0 6 6
use CELL  42
transform -1 0 3684 0 1 1647
box 0 0 6 6
use CELL  43
transform -1 0 2958 0 1 1449
box 0 0 6 6
use CELL  44
transform -1 0 2892 0 -1 1617
box 0 0 6 6
use CELL  45
transform -1 0 2924 0 1 1521
box 0 0 6 6
use CELL  46
transform -1 0 2989 0 1 1503
box 0 0 6 6
use CELL  47
transform -1 0 3818 0 1 1575
box 0 0 6 6
use CELL  48
transform 1 0 3697 0 1 1593
box 0 0 6 6
use CELL  49
transform -1 0 3710 0 1 1494
box 0 0 6 6
use CELL  50
transform -1 0 2986 0 1 1449
box 0 0 6 6
use CELL  51
transform -1 0 3084 0 1 1683
box 0 0 6 6
use CELL  52
transform 1 0 2944 0 1 1431
box 0 0 6 6
use CELL  53
transform -1 0 3893 0 1 1503
box 0 0 6 6
use CELL  54
transform 1 0 3836 0 -1 1464
box 0 0 6 6
use CELL  55
transform 1 0 2945 0 1 1449
box 0 0 6 6
use CELL  56
transform 1 0 3041 0 -1 1653
box 0 0 6 6
use CELL  57
transform -1 0 3074 0 1 1566
box 0 0 6 6
use CELL  58
transform -1 0 3500 0 1 1656
box 0 0 6 6
use CELL  59
transform -1 0 3860 0 -1 1590
box 0 0 6 6
use CELL  60
transform 1 0 2950 0 1 1611
box 0 0 6 6
use CELL  61
transform -1 0 3054 0 1 1647
box 0 0 6 6
use CELL  62
transform -1 0 2938 0 1 1521
box 0 0 6 6
use CELL  63
transform -1 0 3278 0 -1 1428
box 0 0 6 6
use CELL  64
transform -1 0 2960 0 1 1566
box 0 0 6 6
use CELL  65
transform 1 0 2920 0 -1 1563
box 0 0 6 6
use CELL  66
transform -1 0 3834 0 1 1602
box 0 0 6 6
use CELL  67
transform -1 0 2982 0 1 1503
box 0 0 6 6
use CELL  68
transform 1 0 3711 0 1 1629
box 0 0 6 6
use CELL  69
transform -1 0 3735 0 1 1548
box 0 0 6 6
use CELL  70
transform 1 0 3039 0 1 1593
box 0 0 6 6
use CELL  71
transform -1 0 3839 0 1 1584
box 0 0 6 6
use CELL  72
transform -1 0 2959 0 1 1656
box 0 0 6 6
use CELL  73
transform -1 0 3236 0 1 1494
box 0 0 6 6
use CELL  74
transform -1 0 3847 0 1 1593
box 0 0 6 6
use CELL  75
transform -1 0 2922 0 1 1674
box 0 0 6 6
use CELL  76
transform -1 0 2946 0 1 1476
box 0 0 6 6
use CELL  77
transform -1 0 3030 0 1 1683
box 0 0 6 6
use CELL  78
transform -1 0 3491 0 1 1431
box 0 0 6 6
use CELL  79
transform -1 0 2983 0 1 1530
box 0 0 6 6
use CELL  80
transform -1 0 3069 0 1 1647
box 0 0 6 6
use CELL  81
transform -1 0 2953 0 1 1566
box 0 0 6 6
use CELL  82
transform -1 0 2911 0 -1 1626
box 0 0 6 6
use CELL  83
transform -1 0 3804 0 1 1539
box 0 0 6 6
use CELL  84
transform -1 0 3583 0 1 1629
box 0 0 6 6
use CELL  85
transform -1 0 3708 0 1 1566
box 0 0 6 6
use CELL  86
transform -1 0 2990 0 1 1539
box 0 0 6 6
use CELL  87
transform -1 0 3696 0 1 1566
box 0 0 6 6
use CELL  88
transform -1 0 3886 0 1 1503
box 0 0 6 6
use CELL  89
transform -1 0 3910 0 1 1521
box 0 0 6 6
use CELL  90
transform 1 0 2947 0 1 1476
box 0 0 6 6
use CELL  91
transform -1 0 2876 0 1 1611
box 0 0 6 6
use CELL  92
transform -1 0 3512 0 1 1431
box 0 0 6 6
use CELL  93
transform 1 0 3734 0 -1 1581
box 0 0 6 6
use CELL  94
transform 1 0 3810 0 1 1539
box 0 0 6 6
use CELL  95
transform 1 0 3560 0 1 1638
box 0 0 6 6
use CELL  96
transform -1 0 2964 0 1 1629
box 0 0 6 6
use CELL  97
transform -1 0 3271 0 1 1422
box 0 0 6 6
use CELL  98
transform -1 0 3928 0 1 1503
box 0 0 6 6
use CELL  99
transform -1 0 2952 0 1 1629
box 0 0 6 6
use CELL  100
transform 1 0 3821 0 1 1602
box 0 0 6 6
use CELL  101
transform 1 0 3288 0 1 1503
box 0 0 6 6
use CELL  102
transform -1 0 2951 0 1 1647
box 0 0 6 6
use CELL  103
transform -1 0 2958 0 1 1575
box 0 0 6 6
use CELL  104
transform -1 0 3820 0 1 1476
box 0 0 6 6
use CELL  105
transform -1 0 3152 0 1 1494
box 0 0 6 6
use CELL  106
transform 1 0 3778 0 -1 1527
box 0 0 6 6
use CELL  107
transform -1 0 3855 0 -1 1608
box 0 0 6 6
use CELL  108
transform -1 0 3076 0 1 1647
box 0 0 6 6
use CELL  109
transform 1 0 3699 0 1 1647
box 0 0 6 6
use CELL  110
transform 1 0 2994 0 1 1449
box 0 0 6 6
use CELL  111
transform -1 0 2930 0 1 1530
box 0 0 6 6
use CELL  112
transform -1 0 3645 0 1 1656
box 0 0 6 6
use CELL  113
transform -1 0 3144 0 1 1476
box 0 0 6 6
use CELL  114
transform -1 0 2944 0 1 1494
box 0 0 6 6
use CELL  115
transform -1 0 2929 0 1 1512
box 0 0 6 6
use CELL  116
transform -1 0 2989 0 1 1521
box 0 0 6 6
use CELL  117
transform 1 0 2821 0 -1 1644
box 0 0 6 6
use CELL  118
transform 1 0 2814 0 -1 1662
box 0 0 6 6
use CELL  119
transform -1 0 3111 0 1 1521
box 0 0 6 6
use CELL  120
transform -1 0 2952 0 1 1674
box 0 0 6 6
use CELL  121
transform -1 0 3939 0 1 1530
box 0 0 6 6
use CELL  122
transform -1 0 3869 0 1 1539
box 0 0 6 6
use CELL  123
transform -1 0 2972 0 1 1683
box 0 0 6 6
use CELL  124
transform -1 0 2984 0 1 1674
box 0 0 6 6
use CELL  125
transform -1 0 3285 0 1 1422
box 0 0 6 6
use CELL  126
transform -1 0 3088 0 1 1593
box 0 0 6 6
use CELL  127
transform -1 0 3826 0 1 1593
box 0 0 6 6
use CELL  128
transform -1 0 2898 0 1 1467
box 0 0 6 6
use CELL  129
transform -1 0 3496 0 -1 1671
box 0 0 6 6
use CELL  130
transform -1 0 3802 0 1 1566
box 0 0 6 6
use CELL  131
transform -1 0 2943 0 1 1656
box 0 0 6 6
use CELL  132
transform -1 0 2898 0 1 1530
box 0 0 6 6
use CELL  133
transform -1 0 3759 0 1 1584
box 0 0 6 6
use CELL  134
transform -1 0 2972 0 1 1476
box 0 0 6 6
use CELL  135
transform -1 0 2905 0 1 1503
box 0 0 6 6
use CELL  136
transform -1 0 2939 0 1 1476
box 0 0 6 6
use CELL  137
transform -1 0 3909 0 1 1584
box 0 0 6 6
use CELL  138
transform -1 0 2970 0 1 1503
box 0 0 6 6
use CELL  139
transform -1 0 2945 0 -1 1635
box 0 0 6 6
use CELL  140
transform 1 0 3878 0 -1 1500
box 0 0 6 6
use CELL  141
transform -1 0 3654 0 1 1485
box 0 0 6 6
use CELL  142
transform -1 0 2913 0 1 1494
box 0 0 6 6
use CELL  143
transform -1 0 3784 0 1 1512
box 0 0 6 6
use CELL  144
transform -1 0 3825 0 1 1575
box 0 0 6 6
use CELL  145
transform 1 0 2925 0 -1 1590
box 0 0 6 6
use CELL  146
transform -1 0 2935 0 1 1512
box 0 0 6 6
use CELL  147
transform -1 0 3533 0 -1 1437
box 0 0 6 6
use CELL  148
transform -1 0 3653 0 1 1647
box 0 0 6 6
use CELL  149
transform -1 0 3698 0 1 1647
box 0 0 6 6
use CELL  150
transform -1 0 3799 0 1 1602
box 0 0 6 6
use CELL  151
transform 1 0 3902 0 1 1485
box 0 0 6 6
use CELL  152
transform -1 0 3868 0 1 1512
box 0 0 6 6
use CELL  153
transform -1 0 3827 0 1 1557
box 0 0 6 6
use CELL  154
transform -1 0 2944 0 1 1458
box 0 0 6 6
use CELL  155
transform -1 0 3078 0 1 1458
box 0 0 6 6
use CELL  156
transform 1 0 3741 0 -1 1617
box 0 0 6 6
use CELL  157
transform -1 0 3431 0 1 1440
box 0 0 6 6
use CELL  158
transform -1 0 2940 0 1 1557
box 0 0 6 6
use CELL  159
transform -1 0 3854 0 1 1512
box 0 0 6 6
use CELL  160
transform -1 0 3861 0 1 1593
box 0 0 6 6
use CELL  161
transform 1 0 3833 0 1 1575
box 0 0 6 6
use CELL  162
transform -1 0 3094 0 1 1575
box 0 0 6 6
use CELL  163
transform 1 0 3432 0 1 1665
box 0 0 6 6
use CELL  164
transform -1 0 3602 0 1 1611
box 0 0 6 6
use CELL  165
transform -1 0 3739 0 -1 1653
box 0 0 6 6
use CELL  166
transform -1 0 2960 0 1 1620
box 0 0 6 6
use CELL  167
transform -1 0 2967 0 1 1620
box 0 0 6 6
use CELL  168
transform 1 0 3040 0 1 1476
box 0 0 6 6
use CELL  169
transform -1 0 3573 0 1 1503
box 0 0 6 6
use CELL  170
transform -1 0 3875 0 1 1521
box 0 0 6 6
use CELL  171
transform -1 0 2977 0 -1 1419
box 0 0 6 6
use CELL  172
transform -1 0 2898 0 1 1557
box 0 0 6 6
use CELL  173
transform -1 0 2993 0 1 1602
box 0 0 6 6
use CELL  174
transform -1 0 2937 0 1 1458
box 0 0 6 6
use CELL  175
transform -1 0 2972 0 1 1458
box 0 0 6 6
use CELL  176
transform -1 0 2970 0 1 1494
box 0 0 6 6
use CELL  177
transform 1 0 3818 0 -1 1554
box 0 0 6 6
use CELL  178
transform -1 0 3789 0 1 1575
box 0 0 6 6
use CELL  179
transform -1 0 3081 0 1 1674
box 0 0 6 6
use CELL  180
transform 1 0 3835 0 1 1557
box 0 0 6 6
use CELL  181
transform -1 0 2978 0 1 1440
box 0 0 6 6
use CELL  182
transform 1 0 3956 0 1 1503
box 0 0 6 6
use CELL  183
transform -1 0 2924 0 1 1584
box 0 0 6 6
use CELL  184
transform -1 0 2925 0 1 1566
box 0 0 6 6
use CELL  185
transform -1 0 3072 0 1 1665
box 0 0 6 6
use CELL  186
transform 1 0 3732 0 1 1602
box 0 0 6 6
use CELL  187
transform 1 0 3285 0 1 1674
box 0 0 6 6
use CELL  188
transform -1 0 2944 0 1 1449
box 0 0 6 6
use CELL  189
transform -1 0 2970 0 -1 1671
box 0 0 6 6
use CELL  190
transform -1 0 3874 0 1 1503
box 0 0 6 6
use CELL  191
transform -1 0 3689 0 1 1638
box 0 0 6 6
use CELL  192
transform -1 0 3248 0 1 1422
box 0 0 6 6
use CELL  193
transform -1 0 2912 0 1 1584
box 0 0 6 6
use CELL  194
transform -1 0 2919 0 1 1557
box 0 0 6 6
use CELL  195
transform -1 0 3845 0 -1 1554
box 0 0 6 6
use CELL  196
transform -1 0 3033 0 1 1413
box 0 0 6 6
use CELL  197
transform -1 0 3056 0 1 1494
box 0 0 6 6
use CELL  198
transform -1 0 3578 0 1 1539
box 0 0 6 6
use CELL  199
transform -1 0 3876 0 1 1467
box 0 0 6 6
use CELL  200
transform 1 0 3897 0 1 1521
box 0 0 6 6
use CELL  201
transform -1 0 2910 0 1 1629
box 0 0 6 6
use CELL  202
transform -1 0 3921 0 1 1503
box 0 0 6 6
use CELL  203
transform -1 0 3686 0 1 1602
box 0 0 6 6
use CELL  204
transform 1 0 2946 0 1 1467
box 0 0 6 6
use CELL  205
transform -1 0 3188 0 1 1512
box 0 0 6 6
use CELL  206
transform -1 0 2930 0 1 1575
box 0 0 6 6
use CELL  207
transform 1 0 3762 0 1 1611
box 0 0 6 6
use CELL  208
transform -1 0 3020 0 1 1557
box 0 0 6 6
use CELL  209
transform -1 0 2951 0 1 1638
box 0 0 6 6
use CELL  210
transform -1 0 3802 0 -1 1518
box 0 0 6 6
use CELL  211
transform -1 0 3900 0 1 1503
box 0 0 6 6
use CELL  212
transform -1 0 2892 0 1 1512
box 0 0 6 6
use CELL  213
transform 1 0 3605 0 1 1656
box 0 0 6 6
use CELL  214
transform -1 0 2982 0 1 1494
box 0 0 6 6
use CELL  215
transform 1 0 3321 0 -1 1680
box 0 0 6 6
use CELL  216
transform 1 0 3912 0 1 1530
box 0 0 6 6
use CELL  217
transform -1 0 2971 0 1 1440
box 0 0 6 6
use CELL  218
transform -1 0 3841 0 1 1467
box 0 0 6 6
use CELL  219
transform -1 0 2932 0 1 1620
box 0 0 6 6
use CELL  220
transform -1 0 3564 0 1 1440
box 0 0 6 6
use CELL  221
transform 1 0 3840 0 -1 1581
box 0 0 6 6
use CELL  222
transform -1 0 2959 0 1 1539
box 0 0 6 6
use CELL  223
transform -1 0 2992 0 1 1611
box 0 0 6 6
use CELL  224
transform -1 0 3752 0 1 1629
box 0 0 6 6
use CELL  225
transform -1 0 2992 0 1 1512
box 0 0 6 6
use CELL  226
transform -1 0 3020 0 1 1467
box 0 0 6 6
use CELL  227
transform -1 0 3102 0 1 1674
box 0 0 6 6
use CELL  228
transform -1 0 2904 0 1 1449
box 0 0 6 6
use CELL  229
transform -1 0 3069 0 -1 1455
box 0 0 6 6
use CELL  230
transform -1 0 3661 0 1 1611
box 0 0 6 6
use CELL  231
transform -1 0 2972 0 1 1566
box 0 0 6 6
use CELL  232
transform 1 0 3084 0 -1 1590
box 0 0 6 6
use CELL  233
transform -1 0 2919 0 1 1467
box 0 0 6 6
use CELL  234
transform -1 0 3260 0 1 1674
box 0 0 6 6
use CELL  235
transform 1 0 3395 0 1 1431
box 0 0 6 6
use CELL  236
transform -1 0 3042 0 1 1584
box 0 0 6 6
use CELL  237
transform -1 0 3858 0 -1 1572
box 0 0 6 6
use CELL  238
transform -1 0 3775 0 1 1611
box 0 0 6 6
use CELL  239
transform -1 0 3813 0 1 1602
box 0 0 6 6
use CELL  240
transform -1 0 2936 0 1 1602
box 0 0 6 6
use CELL  241
transform -1 0 3832 0 1 1575
box 0 0 6 6
use CELL  242
transform -1 0 3733 0 -1 1617
box 0 0 6 6
use CELL  243
transform -1 0 2838 0 -1 1689
box 0 0 6 6
use CELL  244
transform -1 0 3613 0 1 1620
box 0 0 6 6
use CELL  245
transform 1 0 3720 0 1 1647
box 0 0 6 6
use CELL  246
transform -1 0 2958 0 1 1458
box 0 0 6 6
use CELL  247
transform 1 0 3286 0 -1 1428
box 0 0 6 6
use CELL  248
transform -1 0 3810 0 1 1548
box 0 0 6 6
use CELL  249
transform -1 0 3792 0 1 1557
box 0 0 6 6
use CELL  250
transform 1 0 3327 0 1 1674
box 0 0 6 6
use CELL  251
transform -1 0 3024 0 1 1458
box 0 0 6 6
use CELL  252
transform -1 0 3904 0 1 1467
box 0 0 6 6
use CELL  253
transform -1 0 3078 0 1 1584
box 0 0 6 6
use CELL  254
transform -1 0 2820 0 1 1638
box 0 0 6 6
use CELL  255
transform -1 0 3383 0 1 1431
box 0 0 6 6
use CELL  256
transform 1 0 3871 0 -1 1500
box 0 0 6 6
use CELL  257
transform -1 0 3060 0 1 1476
box 0 0 6 6
use CELL  258
transform -1 0 2970 0 1 1575
box 0 0 6 6
use CELL  259
transform -1 0 3063 0 1 1575
box 0 0 6 6
use CELL  260
transform -1 0 3116 0 1 1656
box 0 0 6 6
use CELL  261
transform -1 0 3848 0 -1 1563
box 0 0 6 6
use CELL  262
transform -1 0 2949 0 1 1422
box 0 0 6 6
use CELL  263
transform -1 0 3789 0 1 1611
box 0 0 6 6
use CELL  264
transform 1 0 3122 0 -1 1500
box 0 0 6 6
use CELL  265
transform -1 0 3792 0 1 1602
box 0 0 6 6
use CELL  266
transform -1 0 3894 0 1 1485
box 0 0 6 6
use CELL  267
transform -1 0 2959 0 1 1584
box 0 0 6 6
use CELL  268
transform -1 0 3627 0 -1 1635
box 0 0 6 6
use CELL  269
transform -1 0 3649 0 1 1620
box 0 0 6 6
use CELL  270
transform -1 0 2931 0 1 1629
box 0 0 6 6
use CELL  271
transform -1 0 3020 0 1 1566
box 0 0 6 6
use CELL  272
transform -1 0 2918 0 1 1449
box 0 0 6 6
use CELL  273
transform 1 0 2822 0 1 1566
box 0 0 6 6
use CELL  274
transform 1 0 2959 0 1 1683
box 0 0 6 6
use CELL  275
transform 1 0 2839 0 -1 1689
box 0 0 6 6
use CELL  276
transform -1 0 2946 0 1 1566
box 0 0 6 6
use CELL  277
transform -1 0 3662 0 1 1494
box 0 0 6 6
use CELL  278
transform -1 0 2925 0 1 1449
box 0 0 6 6
use CELL  279
transform -1 0 3569 0 1 1647
box 0 0 6 6
use CELL  280
transform 1 0 2951 0 -1 1599
box 0 0 6 6
use CELL  281
transform 1 0 2893 0 1 1566
box 0 0 6 6
use CELL  282
transform -1 0 3630 0 1 1467
box 0 0 6 6
use CELL  283
transform 1 0 2892 0 -1 1671
box 0 0 6 6
use CELL  284
transform -1 0 3737 0 1 1620
box 0 0 6 6
use CELL  285
transform 1 0 3821 0 -1 1482
box 0 0 6 6
use CELL  286
transform -1 0 2899 0 1 1512
box 0 0 6 6
use CELL  287
transform 1 0 3052 0 1 1638
box 0 0 6 6
use CELL  288
transform 1 0 3428 0 -1 1545
box 0 0 6 6
use CELL  289
transform 1 0 3813 0 1 1593
box 0 0 6 6
use CELL  290
transform -1 0 3613 0 1 1512
box 0 0 6 6
use CELL  291
transform -1 0 2964 0 1 1440
box 0 0 6 6
use CELL  292
transform 1 0 3141 0 1 1503
box 0 0 6 6
use CELL  293
transform -1 0 2929 0 1 1674
box 0 0 6 6
use CELL  294
transform 1 0 3825 0 1 1548
box 0 0 6 6
use CELL  295
transform 1 0 3918 0 1 1467
box 0 0 6 6
use CELL  296
transform -1 0 3753 0 1 1485
box 0 0 6 6
use CELL  297
transform -1 0 3197 0 1 1431
box 0 0 6 6
use CELL  298
transform -1 0 3008 0 1 1422
box 0 0 6 6
use CELL  299
transform 1 0 3021 0 1 1548
box 0 0 6 6
use CELL  300
transform -1 0 3942 0 -1 1509
box 0 0 6 6
use CELL  301
transform 1 0 3673 0 1 1449
box 0 0 6 6
use CELL  302
transform -1 0 2960 0 1 1476
box 0 0 6 6
use CELL  303
transform 1 0 3834 0 1 1512
box 0 0 6 6
use CELL  304
transform -1 0 2898 0 1 1539
box 0 0 6 6
use CELL  305
transform -1 0 2972 0 1 1449
box 0 0 6 6
use CELL  306
transform -1 0 3848 0 1 1539
box 0 0 6 6
use CELL  307
transform -1 0 3779 0 1 1593
box 0 0 6 6
use CELL  308
transform -1 0 3881 0 1 1584
box 0 0 6 6
use CELL  309
transform -1 0 3081 0 1 1566
box 0 0 6 6
use CELL  310
transform 1 0 3828 0 1 1476
box 0 0 6 6
use CELL  311
transform -1 0 2910 0 1 1593
box 0 0 6 6
use CELL  312
transform -1 0 3925 0 1 1530
box 0 0 6 6
use CELL  313
transform 1 0 3849 0 1 1485
box 0 0 6 6
use CELL  314
transform -1 0 2955 0 1 1665
box 0 0 6 6
use CELL  315
transform 1 0 2930 0 1 1656
box 0 0 6 6
use CELL  316
transform 1 0 3341 0 -1 1680
box 0 0 6 6
use CELL  317
transform -1 0 3741 0 1 1449
box 0 0 6 6
use CELL  318
transform -1 0 2932 0 1 1566
box 0 0 6 6
use CELL  319
transform -1 0 3147 0 1 1521
box 0 0 6 6
use CELL  320
transform 1 0 2907 0 1 1512
box 0 0 6 6
use CELL  321
transform 1 0 2856 0 1 1611
box 0 0 6 6
use CELL  322
transform -1 0 2952 0 1 1521
box 0 0 6 6
use CELL  323
transform -1 0 3799 0 1 1557
box 0 0 6 6
use CELL  324
transform -1 0 3072 0 1 1674
box 0 0 6 6
use CELL  325
transform -1 0 3874 0 1 1584
box 0 0 6 6
use CELL  326
transform -1 0 3833 0 1 1512
box 0 0 6 6
use CELL  327
transform -1 0 2963 0 1 1494
box 0 0 6 6
use CELL  328
transform 1 0 3597 0 1 1440
box 0 0 6 6
use CELL  329
transform -1 0 3732 0 1 1566
box 0 0 6 6
use CELL  330
transform -1 0 3711 0 -1 1554
box 0 0 6 6
use CELL  331
transform 1 0 3724 0 -1 1626
box 0 0 6 6
use CELL  332
transform -1 0 3680 0 1 1539
box 0 0 6 6
use CELL  333
transform -1 0 3016 0 1 1665
box 0 0 6 6
use CELL  334
transform -1 0 3216 0 1 1566
box 0 0 6 6
use CELL  335
transform -1 0 2944 0 1 1575
box 0 0 6 6
use CELL  336
transform -1 0 3236 0 1 1512
box 0 0 6 6
use CELL  337
transform -1 0 2912 0 1 1467
box 0 0 6 6
use CELL  338
transform -1 0 3862 0 1 1557
box 0 0 6 6
use CELL  339
transform 1 0 3633 0 1 1656
box 0 0 6 6
use CELL  340
transform 1 0 2874 0 1 1458
box 0 0 6 6
use CELL  341
transform -1 0 3189 0 1 1422
box 0 0 6 6
use CELL  342
transform 1 0 3811 0 -1 1554
box 0 0 6 6
use CELL  343
transform -1 0 3853 0 1 1584
box 0 0 6 6
use CELL  344
transform -1 0 3320 0 1 1674
box 0 0 6 6
use CELL  345
transform 1 0 3877 0 -1 1473
box 0 0 6 6
use CELL  346
transform -1 0 3076 0 1 1593
box 0 0 6 6
use CELL  347
transform -1 0 3686 0 -1 1455
box 0 0 6 6
use CELL  348
transform -1 0 3609 0 1 1611
box 0 0 6 6
use CELL  349
transform -1 0 3132 0 1 1584
box 0 0 6 6
use CELL  350
transform -1 0 3038 0 1 1539
box 0 0 6 6
use CELL  351
transform 1 0 2944 0 1 1440
box 0 0 6 6
use CELL  352
transform -1 0 3734 0 -1 1545
box 0 0 6 6
use CELL  353
transform -1 0 3652 0 1 1629
box 0 0 6 6
use CELL  354
transform -1 0 3700 0 1 1521
box 0 0 6 6
use CELL  355
transform -1 0 3591 0 -1 1464
box 0 0 6 6
use CELL  356
transform -1 0 2977 0 1 1665
box 0 0 6 6
use CELL  357
transform 1 0 3734 0 1 1494
box 0 0 6 6
use CELL  358
transform 1 0 3414 0 -1 1437
box 0 0 6 6
use CELL  359
transform 1 0 3846 0 1 1548
box 0 0 6 6
use CELL  360
transform -1 0 2930 0 -1 1644
box 0 0 6 6
use CELL  361
transform -1 0 3716 0 1 1620
box 0 0 6 6
use CELL  362
transform 1 0 3831 0 -1 1572
box 0 0 6 6
use CELL  363
transform -1 0 3651 0 1 1584
box 0 0 6 6
use CELL  364
transform 1 0 3810 0 -1 1617
box 0 0 6 6
use CELL  365
transform -1 0 3551 0 1 1647
box 0 0 6 6
use CELL  366
transform -1 0 3809 0 1 1566
box 0 0 6 6
use CELL  367
transform -1 0 3354 0 1 1665
box 0 0 6 6
use CELL  368
transform -1 0 3170 0 1 1539
box 0 0 6 6
use CELL  369
transform -1 0 2985 0 1 1512
box 0 0 6 6
use CELL  370
transform 1 0 2953 0 1 1674
box 0 0 6 6
use CELL  371
transform -1 0 3738 0 1 1503
box 0 0 6 6
use CELL  372
transform 1 0 3848 0 1 1593
box 0 0 6 6
use CELL  373
transform -1 0 2973 0 1 1512
box 0 0 6 6
use CELL  374
transform -1 0 2929 0 1 1593
box 0 0 6 6
use CELL  375
transform -1 0 3008 0 1 1584
box 0 0 6 6
use CELL  376
transform 1 0 2874 0 -1 1473
box 0 0 6 6
use CELL  377
transform 1 0 3038 0 1 1557
box 0 0 6 6
use CELL  378
transform -1 0 3885 0 1 1530
box 0 0 6 6
use CELL  379
transform 1 0 3859 0 -1 1554
box 0 0 6 6
use CELL  380
transform -1 0 2945 0 1 1584
box 0 0 6 6
use CELL  381
transform 1 0 3739 0 -1 1635
box 0 0 6 6
use CELL  382
transform -1 0 3841 0 1 1476
box 0 0 6 6
use CELL  383
transform -1 0 2892 0 1 1575
box 0 0 6 6
use CELL  384
transform 1 0 3703 0 1 1620
box 0 0 6 6
use CELL  385
transform 1 0 3612 0 1 1656
box 0 0 6 6
use CELL  386
transform -1 0 2991 0 1 1674
box 0 0 6 6
use CELL  387
transform -1 0 3636 0 -1 1572
box 0 0 6 6
use CELL  388
transform 1 0 2973 0 1 1449
box 0 0 6 6
use CELL  389
transform -1 0 3915 0 1 1485
box 0 0 6 6
use CELL  390
transform -1 0 3813 0 1 1557
box 0 0 6 6
use CELL  391
transform -1 0 2939 0 1 1566
box 0 0 6 6
use CELL  392
transform -1 0 2931 0 1 1521
box 0 0 6 6
use CELL  393
transform -1 0 3848 0 1 1476
box 0 0 6 6
use CELL  394
transform 1 0 2951 0 1 1440
box 0 0 6 6
use CELL  395
transform -1 0 2930 0 1 1503
box 0 0 6 6
use CELL  396
transform -1 0 2933 0 1 1557
box 0 0 6 6
use CELL  397
transform -1 0 3768 0 1 1566
box 0 0 6 6
use CELL  398
transform -1 0 2898 0 1 1521
box 0 0 6 6
use CELL  399
transform -1 0 3445 0 1 1665
box 0 0 6 6
use CELL  400
transform -1 0 3062 0 1 1485
box 0 0 6 6
use CELL  401
transform -1 0 2953 0 1 1548
box 0 0 6 6
use CELL  402
transform -1 0 2905 0 1 1665
box 0 0 6 6
use CELL  403
transform -1 0 3786 0 1 1584
box 0 0 6 6
use CELL  404
transform -1 0 3766 0 1 1629
box 0 0 6 6
use CELL  405
transform -1 0 3683 0 1 1557
box 0 0 6 6
use CELL  406
transform -1 0 2939 0 1 1548
box 0 0 6 6
use CELL  407
transform 1 0 3584 0 1 1656
box 0 0 6 6
use CELL  408
transform -1 0 3114 0 1 1620
box 0 0 6 6
use CELL  409
transform -1 0 3086 0 1 1494
box 0 0 6 6
use CELL  410
transform -1 0 3710 0 1 1593
box 0 0 6 6
use CELL  411
transform -1 0 2995 0 1 1665
box 0 0 6 6
use CELL  412
transform 1 0 2932 0 -1 1590
box 0 0 6 6
use CELL  413
transform -1 0 3484 0 1 1431
box 0 0 6 6
use CELL  414
transform -1 0 2959 0 1 1521
box 0 0 6 6
use CELL  415
transform 1 0 3911 0 1 1521
box 0 0 6 6
use CELL  416
transform 1 0 2919 0 -1 1446
box 0 0 6 6
use CELL  417
transform -1 0 3051 0 1 1638
box 0 0 6 6
use CELL  418
transform 1 0 3725 0 1 1629
box 0 0 6 6
use CELL  419
transform -1 0 2986 0 1 1602
box 0 0 6 6
use CELL  420
transform -1 0 3615 0 1 1548
box 0 0 6 6
use CELL  421
transform -1 0 3093 0 1 1665
box 0 0 6 6
use CELL  422
transform -1 0 3899 0 1 1530
box 0 0 6 6
use CELL  423
transform -1 0 2905 0 1 1530
box 0 0 6 6
use CELL  424
transform -1 0 2904 0 1 1458
box 0 0 6 6
use CELL  425
transform -1 0 2950 0 1 1656
box 0 0 6 6
use CELL  426
transform -1 0 2937 0 1 1638
box 0 0 6 6
use CELL  427
transform -1 0 3765 0 1 1485
box 0 0 6 6
use CELL  428
transform -1 0 2950 0 1 1593
box 0 0 6 6
use CELL  429
transform -1 0 2953 0 1 1620
box 0 0 6 6
use CELL  430
transform -1 0 3040 0 1 1647
box 0 0 6 6
use CELL  431
transform -1 0 3604 0 1 1656
box 0 0 6 6
use CELL  432
transform -1 0 3081 0 1 1485
box 0 0 6 6
use CELL  433
transform 1 0 3929 0 -1 1509
box 0 0 6 6
use CELL  434
transform -1 0 3482 0 1 1665
box 0 0 6 6
use CELL  435
transform -1 0 3902 0 1 1584
box 0 0 6 6
use CELL  436
transform -1 0 3106 0 1 1638
box 0 0 6 6
use CELL  437
transform -1 0 3006 0 -1 1473
box 0 0 6 6
use CELL  438
transform 1 0 3165 0 1 1449
box 0 0 6 6
use CELL  439
transform 1 0 2809 0 -1 1635
box 0 0 6 6
use CELL  440
transform -1 0 2918 0 1 1548
box 0 0 6 6
use CELL  441
transform -1 0 3929 0 1 1485
box 0 0 6 6
use CELL  442
transform -1 0 3045 0 1 1683
box 0 0 6 6
use CELL  443
transform -1 0 2926 0 1 1467
box 0 0 6 6
use CELL  444
transform 1 0 3835 0 1 1602
box 0 0 6 6
use CELL  445
transform -1 0 2904 0 1 1620
box 0 0 6 6
use CELL  446
transform -1 0 2993 0 1 1449
box 0 0 6 6
use CELL  447
transform -1 0 3128 0 1 1503
box 0 0 6 6
use CELL  448
transform -1 0 3035 0 1 1656
box 0 0 6 6
use CELL  449
transform -1 0 3844 0 1 1521
box 0 0 6 6
use CELL  450
transform -1 0 3123 0 1 1530
box 0 0 6 6
use CELL  451
transform 1 0 2937 0 -1 1599
box 0 0 6 6
use CELL  452
transform -1 0 3817 0 1 1467
box 0 0 6 6
use CELL  453
transform -1 0 3782 0 1 1575
box 0 0 6 6
use CELL  454
transform -1 0 2917 0 1 1629
box 0 0 6 6
use CELL  455
transform -1 0 3519 0 -1 1437
box 0 0 6 6
use CELL  456
transform 1 0 3071 0 1 1656
box 0 0 6 6
use CELL  457
transform 1 0 3817 0 -1 1617
box 0 0 6 6
use CELL  458
transform 1 0 3604 0 1 1440
box 0 0 6 6
use CELL  459
transform -1 0 2923 0 1 1647
box 0 0 6 6
use CELL  460
transform -1 0 2963 0 1 1503
box 0 0 6 6
use CELL  461
transform -1 0 3176 0 1 1467
box 0 0 6 6
use CELL  462
transform -1 0 3135 0 1 1503
box 0 0 6 6
use CELL  463
transform -1 0 2999 0 1 1512
box 0 0 6 6
use CELL  464
transform 1 0 3611 0 1 1440
box 0 0 6 6
use CELL  465
transform -1 0 2932 0 1 1548
box 0 0 6 6
use CELL  466
transform 1 0 3849 0 -1 1563
box 0 0 6 6
use CELL  467
transform 1 0 3772 0 1 1548
box 0 0 6 6
use CELL  468
transform -1 0 3212 0 1 1557
box 0 0 6 6
use CELL  469
transform -1 0 3153 0 1 1530
box 0 0 6 6
use CELL  470
transform 1 0 3908 0 1 1503
box 0 0 6 6
use CELL  471
transform -1 0 2949 0 1 1485
box 0 0 6 6
use CELL  472
transform -1 0 2911 0 1 1440
box 0 0 6 6
use CELL  473
transform 1 0 2990 0 1 1485
box 0 0 6 6
use CELL  474
transform -1 0 2905 0 1 1521
box 0 0 6 6
use CELL  475
transform -1 0 3816 0 1 1566
box 0 0 6 6
use CELL  476
transform -1 0 3590 0 1 1629
box 0 0 6 6
use CELL  477
transform -1 0 2951 0 1 1530
box 0 0 6 6
use CELL  478
transform -1 0 2868 0 1 1602
box 0 0 6 6
use CELL  479
transform -1 0 3087 0 1 1548
box 0 0 6 6
use CELL  480
transform -1 0 3103 0 1 1629
box 0 0 6 6
use CELL  481
transform -1 0 3666 0 1 1485
box 0 0 6 6
use CELL  482
transform -1 0 2898 0 1 1485
box 0 0 6 6
use CELL  483
transform -1 0 3722 0 1 1494
box 0 0 6 6
use CELL  484
transform 1 0 3734 0 -1 1599
box 0 0 6 6
use CELL  485
transform 1 0 2939 0 1 1467
box 0 0 6 6
use CELL  486
transform 1 0 3217 0 1 1422
box 0 0 6 6
use CELL  487
transform 1 0 3745 0 1 1620
box 0 0 6 6
use CELL  488
transform -1 0 3069 0 1 1485
box 0 0 6 6
use CELL  489
transform -1 0 2925 0 -1 1554
box 0 0 6 6
use CELL  490
transform -1 0 3695 0 1 1557
box 0 0 6 6
use CELL  491
transform 1 0 3687 0 -1 1464
box 0 0 6 6
use CELL  492
transform 1 0 3011 0 -1 1464
box 0 0 6 6
use CELL  493
transform -1 0 3862 0 1 1539
box 0 0 6 6
use CELL  494
transform -1 0 3896 0 1 1521
box 0 0 6 6
use CELL  495
transform -1 0 3062 0 1 1512
box 0 0 6 6
use CELL  496
transform 1 0 3618 0 1 1440
box 0 0 6 6
use CELL  497
transform -1 0 3023 0 -1 1671
box 0 0 6 6
use CELL  498
transform 1 0 2951 0 1 1431
box 0 0 6 6
use CELL  499
transform -1 0 2868 0 1 1620
box 0 0 6 6
use CELL  500
transform -1 0 3840 0 1 1593
box 0 0 6 6
use CELL  501
transform -1 0 3705 0 1 1602
box 0 0 6 6
use CELL  502
transform -1 0 3834 0 1 1539
box 0 0 6 6
use CELL  503
transform -1 0 3015 0 1 1584
box 0 0 6 6
use CELL  504
transform -1 0 3804 0 1 1575
box 0 0 6 6
use CELL  505
transform -1 0 2931 0 1 1539
box 0 0 6 6
use CELL  506
transform 1 0 2931 0 1 1647
box 0 0 6 6
use CELL  507
transform -1 0 3740 0 1 1611
box 0 0 6 6
use CELL  508
transform -1 0 3889 0 1 1521
box 0 0 6 6
use CELL  509
transform -1 0 3676 0 1 1521
box 0 0 6 6
use CELL  510
transform -1 0 3732 0 1 1647
box 0 0 6 6
use CELL  511
transform 1 0 3453 0 1 1665
box 0 0 6 6
use CELL  512
transform -1 0 3637 0 1 1620
box 0 0 6 6
use CELL  513
transform -1 0 3879 0 1 1566
box 0 0 6 6
use CELL  514
transform -1 0 3654 0 1 1611
box 0 0 6 6
use CELL  515
transform -1 0 2924 0 1 1539
box 0 0 6 6
use CELL  516
transform -1 0 3049 0 1 1629
box 0 0 6 6
use CELL  517
transform -1 0 2943 0 1 1440
box 0 0 6 6
use CELL  518
transform 1 0 3849 0 1 1467
box 0 0 6 6
use CELL  519
transform -1 0 3392 0 1 1512
box 0 0 6 6
use CELL  520
transform -1 0 3000 0 1 1593
box 0 0 6 6
use CELL  521
transform -1 0 2918 0 1 1620
box 0 0 6 6
use CELL  522
transform 1 0 3676 0 -1 1644
box 0 0 6 6
use CELL  523
transform -1 0 3798 0 1 1458
box 0 0 6 6
use CELL  524
transform -1 0 3724 0 -1 1635
box 0 0 6 6
use CELL  525
transform -1 0 3075 0 1 1575
box 0 0 6 6
use CELL  526
transform -1 0 3549 0 1 1449
box 0 0 6 6
use CELL  527
transform -1 0 3571 0 1 1620
box 0 0 6 6
use CELL  528
transform 1 0 3790 0 -1 1617
box 0 0 6 6
use CELL  529
transform -1 0 2912 0 1 1557
box 0 0 6 6
use CELL  530
transform -1 0 2904 0 1 1575
box 0 0 6 6
use CELL  531
transform 1 0 3824 0 1 1566
box 0 0 6 6
use CELL  532
transform -1 0 2983 0 1 1539
box 0 0 6 6
use CELL  533
transform -1 0 3837 0 1 1494
box 0 0 6 6
use CELL  534
transform -1 0 3039 0 1 1575
box 0 0 6 6
use CELL  535
transform -1 0 3720 0 1 1476
box 0 0 6 6
use CELL  536
transform -1 0 3033 0 1 1422
box 0 0 6 6
use CELL  537
transform -1 0 3010 0 1 1458
box 0 0 6 6
use CELL  538
transform -1 0 2820 0 1 1521
box 0 0 6 6
use CELL  539
transform 1 0 3748 0 1 1611
box 0 0 6 6
use CELL  540
transform -1 0 3589 0 1 1620
box 0 0 6 6
use CELL  541
transform -1 0 2930 0 1 1647
box 0 0 6 6
use CELL  542
transform -1 0 2958 0 1 1530
box 0 0 6 6
use CELL  543
transform -1 0 2938 0 1 1539
box 0 0 6 6
use CELL  544
transform -1 0 3114 0 1 1584
box 0 0 6 6
use CELL  545
transform -1 0 3856 0 1 1458
box 0 0 6 6
use CELL  546
transform -1 0 3618 0 1 1638
box 0 0 6 6
use CELL  547
transform -1 0 3901 0 1 1485
box 0 0 6 6
use CELL  548
transform -1 0 3801 0 1 1584
box 0 0 6 6
use CELL  549
transform -1 0 2996 0 1 1422
box 0 0 6 6
use CELL  550
transform -1 0 3039 0 1 1548
box 0 0 6 6
use CELL  551
transform -1 0 2935 0 -1 1428
box 0 0 6 6
use CELL  552
transform -1 0 3558 0 1 1476
box 0 0 6 6
use CELL  553
transform -1 0 2972 0 1 1422
box 0 0 6 6
use CELL  554
transform -1 0 2821 0 1 1566
box 0 0 6 6
use CELL  555
transform -1 0 3874 0 1 1575
box 0 0 6 6
use CELL  556
transform -1 0 3594 0 1 1584
box 0 0 6 6
use CELL  557
transform 1 0 2938 0 1 1530
box 0 0 6 6
use CELL  558
transform -1 0 3488 0 1 1656
box 0 0 6 6
use CELL  559
transform -1 0 2993 0 1 1593
box 0 0 6 6
use CELL  560
transform -1 0 2986 0 1 1476
box 0 0 6 6
use CELL  561
transform -1 0 2912 0 1 1521
box 0 0 6 6
use CELL  562
transform -1 0 3853 0 1 1575
box 0 0 6 6
use CELL  563
transform -1 0 2971 0 1 1431
box 0 0 6 6
use CELL  564
transform -1 0 2986 0 1 1458
box 0 0 6 6
use CELL  565
transform -1 0 2939 0 1 1620
box 0 0 6 6
use CELL  566
transform -1 0 2979 0 1 1476
box 0 0 6 6
use CELL  567
transform -1 0 2906 0 1 1566
box 0 0 6 6
use CELL  568
transform -1 0 3846 0 1 1530
box 0 0 6 6
use CELL  569
transform -1 0 3703 0 1 1638
box 0 0 6 6
use CELL  570
transform -1 0 2922 0 1 1512
box 0 0 6 6
use CELL  571
transform -1 0 2921 0 1 1611
box 0 0 6 6
use CELL  572
transform -1 0 3013 0 1 1467
box 0 0 6 6
use CELL  573
transform -1 0 3748 0 -1 1518
box 0 0 6 6
use CELL  574
transform -1 0 2965 0 1 1530
box 0 0 6 6
use CELL  575
transform 1 0 2862 0 1 1557
box 0 0 6 6
use CELL  576
transform -1 0 2991 0 1 1647
box 0 0 6 6
use CELL  577
transform -1 0 2862 0 1 1566
box 0 0 6 6
use CELL  578
transform -1 0 3849 0 1 1494
box 0 0 6 6
use CELL  579
transform -1 0 2868 0 1 1593
box 0 0 6 6
use CELL  580
transform -1 0 2880 0 -1 1581
box 0 0 6 6
use CELL  581
transform -1 0 2953 0 1 1683
box 0 0 6 6
use CELL  582
transform 1 0 3874 0 1 1485
box 0 0 6 6
use CELL  583
transform -1 0 3820 0 1 1557
box 0 0 6 6
use CELL  584
transform 1 0 2995 0 1 1584
box 0 0 6 6
use CELL  585
transform 1 0 2993 0 1 1440
box 0 0 6 6
use CELL  586
transform 1 0 3663 0 1 1521
box 0 0 6 6
use CELL  587
transform -1 0 3074 0 1 1467
box 0 0 6 6
use CELL  588
transform -1 0 2983 0 1 1656
box 0 0 6 6
use CELL  589
transform -1 0 3306 0 1 1674
box 0 0 6 6
use CELL  590
transform -1 0 3587 0 1 1647
box 0 0 6 6
use CELL  591
transform -1 0 2946 0 1 1413
box 0 0 6 6
use CELL  592
transform -1 0 3645 0 1 1440
box 0 0 6 6
use CELL  593
transform -1 0 2905 0 1 1584
box 0 0 6 6
use CELL  594
transform -1 0 3744 0 1 1620
box 0 0 6 6
use CELL  595
transform -1 0 2965 0 1 1548
box 0 0 6 6
use CELL  596
transform -1 0 3564 0 1 1620
box 0 0 6 6
use CELL  597
transform -1 0 2814 0 1 1566
box 0 0 6 6
use CELL  598
transform -1 0 3935 0 -1 1491
box 0 0 6 6
use CELL  599
transform -1 0 3129 0 1 1485
box 0 0 6 6
use CELL  600
transform -1 0 3051 0 1 1530
box 0 0 6 6
use CELL  601
transform -1 0 3863 0 1 1521
box 0 0 6 6
use CELL  602
transform -1 0 3863 0 1 1494
box 0 0 6 6
use CELL  603
transform 1 0 3702 0 1 1476
box 0 0 6 6
use CELL  604
transform -1 0 3015 0 1 1674
box 0 0 6 6
use CELL  605
transform 1 0 3171 0 -1 1428
box 0 0 6 6
use CELL  606
transform -1 0 3585 0 1 1449
box 0 0 6 6
use CELL  607
transform -1 0 3766 0 1 1458
box 0 0 6 6
use CELL  608
transform -1 0 3895 0 1 1584
box 0 0 6 6
use CELL  609
transform -1 0 3191 0 1 1557
box 0 0 6 6
use CELL  610
transform 1 0 3850 0 1 1521
box 0 0 6 6
use CELL  611
transform -1 0 3417 0 1 1665
box 0 0 6 6
use CELL  612
transform -1 0 3720 0 1 1467
box 0 0 6 6
use CELL  613
transform -1 0 2978 0 1 1431
box 0 0 6 6
use CELL  614
transform -1 0 3606 0 1 1476
box 0 0 6 6
use CELL  615
transform -1 0 3888 0 1 1584
box 0 0 6 6
use CELL  616
transform -1 0 3660 0 1 1530
box 0 0 6 6
use CELL  617
transform -1 0 2905 0 1 1485
box 0 0 6 6
use CELL  618
transform -1 0 3501 0 1 1521
box 0 0 6 6
use CELL  619
transform -1 0 3855 0 1 1476
box 0 0 6 6
use CELL  620
transform -1 0 3408 0 1 1431
box 0 0 6 6
use CELL  621
transform -1 0 2916 0 1 1647
box 0 0 6 6
use CELL  622
transform -1 0 3844 0 1 1566
box 0 0 6 6
use CELL  623
transform -1 0 2936 0 1 1674
box 0 0 6 6
use CELL  624
transform -1 0 2904 0 1 1602
box 0 0 6 6
use CELL  625
transform 1 0 2802 0 1 1629
box 0 0 6 6
use CELL  626
transform -1 0 2922 0 1 1656
box 0 0 6 6
use CELL  627
transform -1 0 3027 0 1 1593
box 0 0 6 6
use CELL  628
transform -1 0 3775 0 1 1566
box 0 0 6 6
use CELL  629
transform -1 0 2834 0 1 1656
box 0 0 6 6
use CELL  630
transform -1 0 3324 0 1 1620
box 0 0 6 6
use CELL  631
transform 1 0 3805 0 1 1575
box 0 0 6 6
use CELL  632
transform -1 0 2944 0 1 1503
box 0 0 6 6
use CELL  633
transform 1 0 3713 0 1 1647
box 0 0 6 6
use CELL  634
transform 1 0 3799 0 -1 1599
box 0 0 6 6
use CELL  635
transform -1 0 2899 0 1 1611
box 0 0 6 6
use CELL  636
transform -1 0 3459 0 1 1431
box 0 0 6 6
use CELL  637
transform -1 0 3029 0 1 1602
box 0 0 6 6
use CELL  638
transform -1 0 2985 0 1 1440
box 0 0 6 6
use CELL  639
transform -1 0 3609 0 1 1458
box 0 0 6 6
use CELL  640
transform -1 0 2935 0 1 1611
box 0 0 6 6
use CELL  641
transform -1 0 3791 0 1 1458
box 0 0 6 6
use CELL  642
transform 1 0 3603 0 1 1449
box 0 0 6 6
use CELL  643
transform 1 0 3708 0 1 1449
box 0 0 6 6
use CELL  644
transform -1 0 3797 0 1 1539
box 0 0 6 6
use CELL  645
transform -1 0 2946 0 1 1683
box 0 0 6 6
use CELL  646
transform -1 0 3327 0 1 1665
box 0 0 6 6
use CELL  647
transform -1 0 3867 0 1 1530
box 0 0 6 6
use CELL  648
transform -1 0 3830 0 1 1494
box 0 0 6 6
use CELL  649
transform -1 0 2911 0 1 1458
box 0 0 6 6
use CELL  650
transform 1 0 3752 0 1 1620
box 0 0 6 6
use CELL  651
transform -1 0 3907 0 1 1503
box 0 0 6 6
use CELL  652
transform -1 0 2938 0 1 1467
box 0 0 6 6
use CELL  653
transform 1 0 2973 0 -1 1464
box 0 0 6 6
use CELL  654
transform -1 0 3832 0 1 1584
box 0 0 6 6
use CELL  655
transform -1 0 3001 0 1 1413
box 0 0 6 6
use CELL  656
transform -1 0 3034 0 1 1611
box 0 0 6 6
use CELL  657
transform -1 0 3248 0 1 1557
box 0 0 6 6
use CELL  658
transform -1 0 3216 0 1 1422
box 0 0 6 6
use CELL  659
transform -1 0 3773 0 -1 1563
box 0 0 6 6
use CELL  660
transform 1 0 3942 0 1 1503
box 0 0 6 6
use CELL  661
transform 1 0 3499 0 -1 1437
box 0 0 6 6
use CELL  662
transform -1 0 3068 0 1 1557
box 0 0 6 6
use CELL  663
transform -1 0 2997 0 1 1620
box 0 0 6 6
use CELL  664
transform -1 0 3623 0 -1 1473
box 0 0 6 6
use CELL  665
transform -1 0 2820 0 1 1512
box 0 0 6 6
use CELL  666
transform -1 0 2997 0 1 1692
box 0 0 6 6
use CELL  667
transform -1 0 3759 0 1 1458
box 0 0 6 6
use CELL  668
transform 1 0 3892 0 1 1494
box 0 0 6 6
use CELL  669
transform -1 0 3285 0 1 1476
box 0 0 6 6
use CELL  670
transform 1 0 3002 0 1 1656
box 0 0 6 6
use CELL  671
transform -1 0 2869 0 1 1566
box 0 0 6 6
use CELL  672
transform -1 0 3102 0 1 1620
box 0 0 6 6
use CELL  673
transform -1 0 3806 0 1 1602
box 0 0 6 6
use CELL  674
transform -1 0 2992 0 1 1440
box 0 0 6 6
use CELL  675
transform -1 0 3738 0 1 1629
box 0 0 6 6
use CELL  676
transform -1 0 3678 0 1 1530
box 0 0 6 6
use CELL  677
transform 1 0 2930 0 1 1593
box 0 0 6 6
use CELL  678
transform -1 0 3137 0 1 1602
box 0 0 6 6
use CELL  679
transform -1 0 3867 0 1 1584
box 0 0 6 6
use CELL  680
transform -1 0 3771 0 1 1548
box 0 0 6 6
use CELL  681
transform -1 0 3237 0 1 1485
box 0 0 6 6
use CELL  682
transform -1 0 3885 0 -1 1572
box 0 0 6 6
use CELL  683
transform -1 0 2905 0 1 1611
box 0 0 6 6
use CELL  684
transform -1 0 2963 0 -1 1428
box 0 0 6 6
use CELL  685
transform -1 0 3122 0 1 1611
box 0 0 6 6
use CELL  686
transform -1 0 2929 0 1 1656
box 0 0 6 6
use CELL  687
transform 1 0 3646 0 1 1656
box 0 0 6 6
use CELL  688
transform -1 0 3583 0 -1 1662
box 0 0 6 6
use CELL  689
transform -1 0 2943 0 1 1431
box 0 0 6 6
use CELL  690
transform -1 0 3851 0 1 1566
box 0 0 6 6
use CELL  691
transform -1 0 3798 0 1 1593
box 0 0 6 6
use CELL  692
transform -1 0 2959 0 1 1467
box 0 0 6 6
use CELL  693
transform 1 0 3884 0 1 1467
box 0 0 6 6
use CELL  694
transform 1 0 3799 0 1 1458
box 0 0 6 6
use CELL  695
transform -1 0 2979 0 1 1548
box 0 0 6 6
use CELL  696
transform -1 0 2943 0 1 1674
box 0 0 6 6
use CELL  697
transform 1 0 2986 0 1 1431
box 0 0 6 6
use CELL  698
transform -1 0 3053 0 1 1476
box 0 0 6 6
use CELL  699
transform -1 0 2925 0 1 1476
box 0 0 6 6
use CELL  700
transform -1 0 3862 0 1 1602
box 0 0 6 6
use CELL  701
transform 1 0 3882 0 1 1575
box 0 0 6 6
use CELL  702
transform 1 0 3251 0 -1 1428
box 0 0 6 6
use CELL  703
transform 1 0 3866 0 -1 1572
box 0 0 6 6
use CELL  704
transform 1 0 3701 0 1 1449
box 0 0 6 6
use CELL  705
transform -1 0 3015 0 1 1422
box 0 0 6 6
use CELL  706
transform -1 0 2956 0 1 1503
box 0 0 6 6
use CELL  707
transform -1 0 2942 0 1 1422
box 0 0 6 6
use CELL  708
transform -1 0 2946 0 -1 1626
box 0 0 6 6
use CELL  709
transform -1 0 3264 0 -1 1428
box 0 0 6 6
use CELL  710
transform -1 0 2918 0 1 1440
box 0 0 6 6
use CELL  711
transform -1 0 3783 0 1 1485
box 0 0 6 6
use CELL  712
transform -1 0 3897 0 1 1467
box 0 0 6 6
use CELL  713
transform -1 0 3503 0 1 1440
box 0 0 6 6
use CELL  714
transform -1 0 2911 0 1 1548
box 0 0 6 6
use CELL  715
transform -1 0 3614 0 1 1557
box 0 0 6 6
use CELL  716
transform -1 0 2918 0 1 1476
box 0 0 6 6
use CELL  717
transform -1 0 2985 0 1 1431
box 0 0 6 6
use CELL  718
transform 1 0 3655 0 -1 1644
box 0 0 6 6
use CELL  719
transform -1 0 2906 0 1 1512
box 0 0 6 6
use CELL  720
transform -1 0 2924 0 1 1629
box 0 0 6 6
use CELL  721
transform -1 0 2904 0 -1 1437
box 0 0 6 6
use CELL  722
transform -1 0 3033 0 1 1530
box 0 0 6 6
use CELL  723
transform 1 0 2983 0 1 1485
box 0 0 6 6
use CELL  724
transform 1 0 3235 0 1 1422
box 0 0 6 6
use CELL  725
transform 1 0 3481 0 1 1638
box 0 0 6 6
use CELL  726
transform -1 0 2965 0 1 1458
box 0 0 6 6
use CELL  727
transform -1 0 3719 0 -1 1563
box 0 0 6 6
use CELL  728
transform -1 0 3066 0 1 1683
box 0 0 6 6
use CELL  729
transform -1 0 3814 0 1 1512
box 0 0 6 6
use CELL  730
transform -1 0 2937 0 1 1503
box 0 0 6 6
use CELL  731
transform 1 0 3626 0 1 1656
box 0 0 6 6
use CELL  732
transform -1 0 3691 0 1 1512
box 0 0 6 6
use CELL  733
transform -1 0 3019 0 1 1629
box 0 0 6 6
use CELL  734
transform 1 0 3602 0 1 1602
box 0 0 6 6
use CELL  735
transform 1 0 3035 0 -1 1617
box 0 0 6 6
use CELL  736
transform -1 0 3044 0 1 1503
box 0 0 6 6
use CELL  737
transform -1 0 2984 0 1 1647
box 0 0 6 6
use CELL  738
transform 1 0 2922 0 -1 1617
box 0 0 6 6
use CELL  739
transform -1 0 3865 0 1 1566
box 0 0 6 6
use CELL  740
transform 1 0 2898 0 -1 1446
box 0 0 6 6
use CELL  741
transform 1 0 3437 0 1 1440
box 0 0 6 6
use CELL  742
transform -1 0 2942 0 1 1611
box 0 0 6 6
use CELL  743
transform 1 0 2926 0 -1 1482
box 0 0 6 6
use CELL  744
transform -1 0 2923 0 1 1638
box 0 0 6 6
use CELL  745
transform -1 0 2925 0 1 1431
box 0 0 6 6
use CELL  746
transform -1 0 2998 0 1 1647
box 0 0 6 6
use CELL  747
transform -1 0 3155 0 1 1602
box 0 0 6 6
use CELL  748
transform -1 0 3057 0 1 1422
box 0 0 6 6
use CELL  749
transform -1 0 2934 0 1 1665
box 0 0 6 6
use CELL  750
transform -1 0 3946 0 -1 1536
box 0 0 6 6
use CELL  751
transform -1 0 3960 0 1 1530
box 0 0 6 6
use CELL  752
transform -1 0 3820 0 1 1602
box 0 0 6 6
use CELL  753
transform -1 0 3060 0 1 1620
box 0 0 6 6
use CELL  754
transform -1 0 3018 0 1 1638
box 0 0 6 6
use CELL  755
transform -1 0 3402 0 1 1665
box 0 0 6 6
use CELL  756
transform -1 0 3086 0 1 1440
box 0 0 6 6
use CELL  757
transform -1 0 3855 0 1 1503
box 0 0 6 6
use CELL  758
transform 1 0 3479 0 1 1440
box 0 0 6 6
use CELL  759
transform 1 0 3881 0 -1 1491
box 0 0 6 6
use CELL  760
transform -1 0 3573 0 1 1638
box 0 0 6 6
use CELL  761
transform 1 0 3837 0 1 1485
box 0 0 6 6
use CELL  762
transform -1 0 3693 0 1 1449
box 0 0 6 6
use CELL  763
transform -1 0 3673 0 1 1611
box 0 0 6 6
use CELL  764
transform -1 0 2943 0 1 1602
box 0 0 6 6
use CELL  765
transform -1 0 3823 0 1 1566
box 0 0 6 6
use CELL  766
transform -1 0 2938 0 1 1629
box 0 0 6 6
use CELL  767
transform -1 0 2990 0 1 1530
box 0 0 6 6
use CELL  768
transform -1 0 3723 0 -1 1626
box 0 0 6 6
use CELL  769
transform -1 0 3668 0 1 1638
box 0 0 6 6
use CELL  770
transform 1 0 3051 0 1 1593
box 0 0 6 6
use CELL  771
transform -1 0 3810 0 1 1467
box 0 0 6 6
use CELL  772
transform -1 0 3846 0 -1 1590
box 0 0 6 6
use CELL  773
transform -1 0 3647 0 1 1494
box 0 0 6 6
use CELL  774
transform -1 0 3809 0 1 1611
box 0 0 6 6
use CELL  775
transform -1 0 3870 0 1 1494
box 0 0 6 6
use CELL  776
transform -1 0 2892 0 1 1566
box 0 0 6 6
use CELL  777
transform -1 0 3821 0 1 1458
box 0 0 6 6
use CELL  778
transform -1 0 3069 0 1 1593
box 0 0 6 6
use CELL  779
transform -1 0 3862 0 1 1503
box 0 0 6 6
use CELL  780
transform -1 0 3847 0 1 1512
box 0 0 6 6
use CELL  781
transform -1 0 3738 0 1 1467
box 0 0 6 6
use CELL  782
transform -1 0 3507 0 1 1656
box 0 0 6 6
use CELL  783
transform -1 0 3632 0 1 1539
box 0 0 6 6
use CELL  784
transform -1 0 2934 0 1 1413
box 0 0 6 6
use CELL  785
transform -1 0 3712 0 -1 1653
box 0 0 6 6
use CELL  786
transform -1 0 2996 0 1 1521
box 0 0 6 6
use CELL  787
transform -1 0 3589 0 1 1440
box 0 0 6 6
use CELL  788
transform -1 0 3710 0 -1 1635
box 0 0 6 6
use CELL  789
transform -1 0 3750 0 1 1503
box 0 0 6 6
use CELL  790
transform -1 0 3858 0 1 1548
box 0 0 6 6
use CELL  791
transform -1 0 2945 0 1 1521
box 0 0 6 6
use CELL  792
transform -1 0 3932 0 1 1530
box 0 0 6 6
use CELL  793
transform -1 0 3826 0 1 1521
box 0 0 6 6
use CELL  794
transform 1 0 2910 0 -1 1644
box 0 0 6 6
use CELL  795
transform -1 0 2966 0 1 1674
box 0 0 6 6
use CELL  796
transform -1 0 3883 0 1 1539
box 0 0 6 6
use CELL  797
transform 1 0 3856 0 1 1485
box 0 0 6 6
use CELL  798
transform 1 0 3492 0 -1 1437
box 0 0 6 6
use CELL  799
transform -1 0 3955 0 1 1503
box 0 0 6 6
use CELL  800
transform -1 0 2912 0 1 1611
box 0 0 6 6
use CELL  801
transform -1 0 3625 0 1 1593
box 0 0 6 6
use CELL  802
transform -1 0 3017 0 1 1431
box 0 0 6 6
use CELL  803
transform -1 0 3881 0 1 1575
box 0 0 6 6
use CELL  804
transform -1 0 3696 0 1 1638
box 0 0 6 6
use CELL  805
transform -1 0 2966 0 1 1557
box 0 0 6 6
use CELL  806
transform -1 0 3867 0 -1 1581
box 0 0 6 6
use CELL  807
transform 1 0 3590 0 1 1440
box 0 0 6 6
use CELL  808
transform -1 0 3424 0 1 1575
box 0 0 6 6
use CELL  809
transform -1 0 2814 0 -1 1455
box 0 0 6 6
use CELL  810
transform -1 0 3917 0 1 1467
box 0 0 6 6
use CELL  811
transform -1 0 3838 0 1 1548
box 0 0 6 6
use CELL  812
transform -1 0 2950 0 1 1602
box 0 0 6 6
use CELL  813
transform -1 0 2930 0 1 1602
box 0 0 6 6
use CELL  814
transform -1 0 2949 0 1 1611
box 0 0 6 6
use CELL  815
transform -1 0 3098 0 1 1656
box 0 0 6 6
use CELL  816
transform -1 0 2911 0 1 1431
box 0 0 6 6
use CELL  817
transform 1 0 2935 0 -1 1671
box 0 0 6 6
use CELL  818
transform 1 0 3855 0 -1 1518
box 0 0 6 6
use CELL  819
transform -1 0 3862 0 1 1467
box 0 0 6 6
use CELL  820
transform -1 0 3284 0 1 1674
box 0 0 6 6
use CELL  821
transform -1 0 3285 0 1 1665
box 0 0 6 6
use CELL  822
transform -1 0 2999 0 1 1638
box 0 0 6 6
use CELL  823
transform -1 0 3760 0 1 1521
box 0 0 6 6
use CELL  824
transform -1 0 2925 0 1 1494
box 0 0 6 6
use CELL  825
transform -1 0 3788 0 1 1494
box 0 0 6 6
use CELL  826
transform -1 0 2905 0 1 1539
box 0 0 6 6
use CELL  827
transform -1 0 3875 0 1 1512
box 0 0 6 6
use CELL  828
transform -1 0 3691 0 1 1647
box 0 0 6 6
use CELL  829
transform -1 0 3119 0 1 1602
box 0 0 6 6
use CELL  830
transform -1 0 3077 0 -1 1437
box 0 0 6 6
use CELL  831
transform -1 0 3091 0 1 1683
box 0 0 6 6
use CELL  832
transform -1 0 2963 0 1 1485
box 0 0 6 6
use CELL  833
transform -1 0 3784 0 1 1458
box 0 0 6 6
use CELL  834
transform 1 0 3663 0 1 1548
box 0 0 6 6
use CELL  835
transform -1 0 3654 0 1 1449
box 0 0 6 6
use CELL  836
transform -1 0 3803 0 1 1611
box 0 0 6 6
use CELL  837
transform -1 0 3855 0 1 1539
box 0 0 6 6
use CELL  838
transform -1 0 2942 0 1 1512
box 0 0 6 6
use CELL  839
transform -1 0 3062 0 1 1503
box 0 0 6 6
use CELL  840
transform -1 0 3855 0 1 1530
box 0 0 6 6
use CELL  841
transform -1 0 2925 0 1 1620
box 0 0 6 6
use CELL  842
transform -1 0 3808 0 1 1584
box 0 0 6 6
use CELL  843
transform -1 0 2956 0 1 1494
box 0 0 6 6
use CELL  844
transform -1 0 3001 0 1 1656
box 0 0 6 6
use CELL  845
transform -1 0 3812 0 1 1593
box 0 0 6 6
use CELL  846
transform -1 0 2911 0 1 1449
box 0 0 6 6
use CELL  847
transform -1 0 3218 0 1 1539
box 0 0 6 6
use CELL  848
transform -1 0 3041 0 1 1602
box 0 0 6 6
use CELL  849
transform 1 0 2964 0 -1 1419
box 0 0 6 6
use CELL  850
transform -1 0 2904 0 1 1548
box 0 0 6 6
use CELL  851
transform -1 0 3531 0 1 1449
box 0 0 6 6
use CELL  852
transform -1 0 3535 0 1 1638
box 0 0 6 6
use CELL  853
transform -1 0 3780 0 1 1557
box 0 0 6 6
use CELL  854
transform -1 0 2862 0 1 1575
box 0 0 6 6
use CELL  855
transform 1 0 3778 0 1 1476
box 0 0 6 6
use CELL  856
transform -1 0 3792 0 1 1530
box 0 0 6 6
use CELL  857
transform -1 0 2922 0 1 1593
box 0 0 6 6
use CELL  858
transform -1 0 3351 0 1 1485
box 0 0 6 6
use CELL  859
transform -1 0 3523 0 1 1638
box 0 0 6 6
use CELL  860
transform 1 0 3625 0 1 1440
box 0 0 6 6
use CELL  861
transform -1 0 3911 0 1 1530
box 0 0 6 6
use CELL  862
transform -1 0 2932 0 1 1494
box 0 0 6 6
use CELL  863
transform -1 0 3198 0 1 1566
box 0 0 6 6
use CELL  864
transform -1 0 2947 0 1 1557
box 0 0 6 6
use CELL  865
transform 1 0 2954 0 1 1647
box 0 0 6 6
use CELL  866
transform -1 0 3597 0 1 1629
box 0 0 6 6
use CELL  867
transform -1 0 3026 0 1 1539
box 0 0 6 6
use CELL  868
transform -1 0 3813 0 1 1476
box 0 0 6 6
use CELL  869
transform -1 0 3735 0 1 1449
box 0 0 6 6
use CELL  870
transform -1 0 2925 0 -1 1464
box 0 0 6 6
use CELL  871
transform -1 0 2827 0 1 1656
box 0 0 6 6
use CELL  872
transform -1 0 3661 0 1 1449
box 0 0 6 6
use CELL  873
transform 1 0 3591 0 -1 1662
box 0 0 6 6
use CELL  874
transform -1 0 3431 0 1 1665
box 0 0 6 6
use CELL  875
transform -1 0 3876 0 1 1539
box 0 0 6 6
use CELL  876
transform -1 0 3255 0 1 1521
box 0 0 6 6
use CELL  877
transform 1 0 3534 0 1 1431
box 0 0 6 6
use CELL  878
transform -1 0 3098 0 1 1683
box 0 0 6 6
use CELL  879
transform -1 0 2899 0 1 1494
box 0 0 6 6
use CELL  880
transform -1 0 2954 0 1 1557
box 0 0 6 6
use CELL  881
transform -1 0 2979 0 1 1683
box 0 0 6 6
use CELL  882
transform -1 0 3953 0 -1 1536
box 0 0 6 6
use CELL  883
transform -1 0 3814 0 1 1458
box 0 0 6 6
use CELL  884
transform -1 0 3634 0 1 1629
box 0 0 6 6
use CELL  885
transform -1 0 3110 0 1 1440
box 0 0 6 6
use CELL  886
transform 1 0 3790 0 1 1548
box 0 0 6 6
use CELL  887
transform -1 0 2956 0 1 1485
box 0 0 6 6
use CELL  888
transform -1 0 3777 0 -1 1482
box 0 0 6 6
use CELL  889
transform -1 0 3260 0 1 1611
box 0 0 6 6
use CELL  890
transform -1 0 2922 0 -1 1671
box 0 0 6 6
use CELL  891
transform -1 0 2918 0 -1 1464
box 0 0 6 6
use CELL  892
transform -1 0 3782 0 -1 1617
box 0 0 6 6
use CELL  893
transform -1 0 2923 0 1 1602
box 0 0 6 6
use CELL  894
transform -1 0 3696 0 1 1476
box 0 0 6 6
use CELL  895
transform -1 0 2937 0 1 1485
box 0 0 6 6
use CELL  896
transform -1 0 3349 0 1 1629
box 0 0 6 6
use CELL  897
transform 1 0 3715 0 1 1449
box 0 0 6 6
use CELL  898
transform -1 0 2997 0 1 1530
box 0 0 6 6
use CELL  899
transform 1 0 2958 0 -1 1437
box 0 0 6 6
use CELL  900
transform -1 0 2994 0 1 1629
box 0 0 6 6
use CELL  901
transform -1 0 3764 0 1 1620
box 0 0 6 6
use CELL  902
transform 1 0 2928 0 1 1683
box 0 0 6 6
use CELL  903
transform -1 0 3253 0 1 1674
box 0 0 6 6
use CELL  904
transform 1 0 2898 0 1 1656
box 0 0 6 6
use CELL  905
transform -1 0 3452 0 1 1665
box 0 0 6 6
use CELL  906
transform -1 0 3860 0 1 1575
box 0 0 6 6
use CELL  907
transform -1 0 3065 0 1 1665
box 0 0 6 6
use CELL  908
transform -1 0 3733 0 1 1575
box 0 0 6 6
use CELL  909
transform -1 0 3849 0 1 1458
box 0 0 6 6
use CELL  910
transform -1 0 2869 0 1 1611
box 0 0 6 6
use CELL  911
transform -1 0 3765 0 1 1476
box 0 0 6 6
use CELL  912
transform -1 0 3246 0 1 1674
box 0 0 6 6
use CELL  913
transform -1 0 3176 0 1 1611
box 0 0 6 6
use CELL  914
transform -1 0 3606 0 1 1512
box 0 0 6 6
use CELL  915
transform -1 0 2923 0 1 1575
box 0 0 6 6
use CELL  916
transform 1 0 3758 0 -1 1581
box 0 0 6 6
use CELL  917
transform -1 0 2991 0 1 1548
box 0 0 6 6
use CELL  918
transform -1 0 3473 0 1 1665
box 0 0 6 6
use CELL  919
transform -1 0 3582 0 1 1440
box 0 0 6 6
use CELL  920
transform -1 0 3790 0 1 1566
box 0 0 6 6
use CELL  921
transform -1 0 3340 0 -1 1680
box 0 0 6 6
use CELL  922
transform -1 0 3890 0 1 1539
box 0 0 6 6
use CELL  923
transform -1 0 3922 0 1 1485
box 0 0 6 6
use CELL  924
transform -1 0 3599 0 -1 1518
box 0 0 6 6
use CELL  925
transform -1 0 3638 0 1 1440
box 0 0 6 6
use CELL  926
transform 1 0 3051 0 1 1683
box 0 0 6 6
use CELL  927
transform -1 0 3848 0 1 1602
box 0 0 6 6
use CELL  928
transform -1 0 2966 0 1 1467
box 0 0 6 6
use CELL  929
transform -1 0 3759 0 1 1629
box 0 0 6 6
use CELL  930
transform -1 0 2937 0 -1 1581
box 0 0 6 6
use CELL  931
transform -1 0 3625 0 1 1656
box 0 0 6 6
use CELL  932
transform -1 0 2918 0 1 1431
box 0 0 6 6
use CELL  933
transform -1 0 3050 0 1 1539
box 0 0 6 6
use CELL  934
transform 1 0 3288 0 1 1566
box 0 0 6 6
use CELL  935
transform -1 0 3654 0 1 1503
box 0 0 6 6
use CELL  936
transform -1 0 3489 0 1 1665
box 0 0 6 6
use CELL  937
transform 1 0 2899 0 1 1467
box 0 0 6 6
use CELL  938
transform -1 0 2969 0 1 1638
box 0 0 6 6
use CELL  939
transform -1 0 3053 0 1 1602
box 0 0 6 6
use CELL  940
transform -1 0 2916 0 1 1422
box 0 0 6 6
use CELL  941
transform -1 0 2898 0 1 1503
box 0 0 6 6
use CELL  942
transform -1 0 2951 0 1 1458
box 0 0 6 6
use CELL  943
transform 1 0 3020 0 1 1440
box 0 0 6 6
use CELL  944
transform -1 0 3542 0 1 1638
box 0 0 6 6
use CELL  945
transform -1 0 3134 0 1 1611
box 0 0 6 6
use CELL  946
transform -1 0 2892 0 -1 1500
box 0 0 6 6
use CELL  947
transform 1 0 3829 0 1 1458
box 0 0 6 6
use CELL  948
transform -1 0 3833 0 1 1593
box 0 0 6 6
use CELL  949
transform -1 0 3711 0 1 1458
box 0 0 6 6
use CELL  950
transform 1 0 2964 0 1 1485
box 0 0 6 6
use CELL  951
transform 1 0 3863 0 1 1467
box 0 0 6 6
use CELL  952
transform -1 0 2973 0 1 1467
box 0 0 6 6
use CELL  953
transform 1 0 3835 0 -1 1545
box 0 0 6 6
use CELL  954
transform -1 0 2912 0 1 1503
box 0 0 6 6
use CELL  955
transform -1 0 3087 0 1 1575
box 0 0 6 6
use CELL  956
transform -1 0 2945 0 1 1539
box 0 0 6 6
use CELL  957
transform 1 0 2976 0 1 1485
box 0 0 6 6
use CELL  958
transform -1 0 3014 0 1 1521
box 0 0 6 6
use CELL  959
transform -1 0 2989 0 1 1494
box 0 0 6 6
use CELL  960
transform -1 0 3571 0 1 1656
box 0 0 6 6
use CELL  961
transform -1 0 3040 0 1 1413
box 0 0 6 6
use CELL  962
transform -1 0 2898 0 1 1584
box 0 0 6 6
use CELL  963
transform -1 0 3882 0 1 1521
box 0 0 6 6
use CELL  964
transform -1 0 3752 0 1 1539
box 0 0 6 6
use CELL  965
transform -1 0 3911 0 1 1467
box 0 0 6 6
use CELL  966
transform -1 0 3924 0 1 1521
box 0 0 6 6
use CELL  967
transform -1 0 3001 0 1 1629
box 0 0 6 6
use CELL  968
transform -1 0 2972 0 1 1548
box 0 0 6 6
use CELL  969
transform -1 0 3466 0 -1 1671
box 0 0 6 6
use CELL  970
transform -1 0 2956 0 1 1422
box 0 0 6 6
use CELL  971
transform -1 0 2999 0 1 1431
box 0 0 6 6
use CELL  972
transform -1 0 2996 0 -1 1500
box 0 0 6 6
use CELL  973
transform 1 0 3538 0 1 1647
box 0 0 6 6
use CELL  974
transform -1 0 2952 0 1 1692
box 0 0 6 6
use CELL  975
transform -1 0 3821 0 1 1512
box 0 0 6 6
use CELL  976
transform 1 0 2946 0 -1 1590
box 0 0 6 6
use CELL  977
transform -1 0 2946 0 1 1548
box 0 0 6 6
use CELL  978
transform -1 0 2996 0 1 1503
box 0 0 6 6
use CELL  979
transform -1 0 2937 0 1 1449
box 0 0 6 6
use CELL  980
transform -1 0 2820 0 1 1557
box 0 0 6 6
use CELL  981
transform -1 0 2911 0 1 1575
box 0 0 6 6
use CELL  982
transform -1 0 3818 0 1 1494
box 0 0 6 6
use CELL  983
transform -1 0 3700 0 1 1449
box 0 0 6 6
use CELL  984
transform -1 0 3891 0 1 1494
box 0 0 6 6
use CELL  985
transform 1 0 2821 0 -1 1527
box 0 0 6 6
use CELL  986
transform -1 0 3219 0 1 1530
box 0 0 6 6
use CELL  987
transform -1 0 3828 0 1 1458
box 0 0 6 6
use CELL  988
transform 1 0 3722 0 1 1449
box 0 0 6 6
use CELL  989
transform -1 0 3791 0 1 1593
box 0 0 6 6
use CELL  990
transform 1 0 2821 0 -1 1518
box 0 0 6 6
use CELL  991
transform 1 0 2931 0 1 1530
box 0 0 6 6
use CELL  992
transform -1 0 3856 0 1 1494
box 0 0 6 6
use CELL  993
transform -1 0 2965 0 1 1449
box 0 0 6 6
use CELL  994
transform -1 0 3015 0 1 1575
box 0 0 6 6
use CELL  995
transform -1 0 2905 0 1 1557
box 0 0 6 6
use CELL  996
transform -1 0 3006 0 1 1638
box 0 0 6 6
use CELL  997
transform 1 0 2906 0 -1 1545
box 0 0 6 6
use CELL  998
transform 1 0 2898 0 -1 1482
box 0 0 6 6
use CELL  999
transform 1 0 3520 0 1 1431
box 0 0 6 6
use CELL  1000
transform 1 0 2815 0 -1 1455
box 0 0 6 6
<< metal1 >>
rect 3221 1420 3222 1423
rect 3221 1420 3489 1421
rect 3489 1420 3490 1431
rect 3815 1474 3816 1477
rect 3815 1474 3818 1475
rect 3818 1465 3819 1475
rect 3806 1465 3819 1466
rect 3806 1456 3807 1466
rect 3806 1456 3837 1457
rect 3837 1456 3838 1458
rect 3635 1573 3636 1621
rect 3435 1573 3636 1574
rect 3435 1537 3436 1574
rect 3429 1537 3436 1538
rect 3429 1537 3430 1539
rect 3708 1627 3709 1630
rect 3007 1627 3709 1628
rect 3007 1627 3008 1654
rect 2993 1654 3008 1655
rect 2993 1654 2994 1665
rect 2822 1519 2823 1522
rect 2815 1519 2823 1520
rect 2815 1519 2816 1521
rect 3920 1483 3921 1486
rect 3803 1483 3921 1484
rect 3803 1483 3804 1537
rect 3795 1537 3804 1538
rect 3795 1537 3796 1539
rect 2995 1600 2996 1621
rect 2995 1600 3106 1601
rect 3106 1582 3107 1601
rect 3106 1582 3112 1583
rect 3112 1582 3113 1584
rect 2914 1555 2915 1558
rect 2914 1555 2958 1556
rect 2958 1555 2959 1564
rect 2958 1564 2961 1565
rect 2961 1564 2962 1573
rect 2949 1573 2962 1574
rect 2949 1573 2950 1575
rect 2957 1465 2958 1468
rect 2957 1465 2974 1466
rect 2974 1465 2975 1474
rect 2964 1474 2975 1475
rect 2964 1474 2965 1483
rect 2964 1483 2971 1484
rect 2971 1483 2972 1492
rect 2958 1492 2972 1493
rect 2958 1492 2959 1494
rect 3664 1553 3665 1555
rect 3437 1555 3665 1556
rect 3437 1535 3438 1556
rect 3220 1535 3438 1536
rect 3220 1535 3221 1546
rect 3196 1546 3221 1547
rect 3196 1546 3197 1548
rect 2906 1429 2907 1432
rect 2906 1429 2929 1430
rect 2929 1429 2930 1456
rect 2929 1456 2998 1457
rect 2998 1456 2999 1510
rect 2998 1510 3000 1511
rect 3000 1510 3001 1519
rect 2987 1519 3001 1520
rect 2987 1519 2988 1521
rect 3123 1501 3124 1504
rect 3002 1501 3124 1502
rect 3002 1501 3003 1528
rect 2914 1528 3003 1529
rect 2914 1483 2915 1529
rect 2890 1483 2915 1484
rect 2890 1465 2891 1484
rect 2890 1465 2907 1466
rect 2907 1465 2908 1467
rect 3594 1510 3595 1513
rect 3576 1510 3595 1511
rect 3576 1510 3577 1539
rect 2928 1636 2929 1639
rect 2928 1636 2949 1637
rect 2949 1636 2950 1638
rect 3885 1472 3886 1481
rect 3885 1481 3936 1482
rect 3936 1481 3937 1501
rect 3878 1501 3937 1502
rect 3878 1501 3879 1519
rect 3878 1519 3891 1520
rect 3891 1519 3892 1521
rect 3011 1645 3012 1666
rect 3011 1645 3071 1646
rect 3071 1645 3072 1647
rect 2978 1537 2979 1540
rect 2890 1537 2979 1538
rect 2890 1528 2891 1538
rect 2890 1528 2907 1529
rect 2907 1528 2908 1530
rect 2867 1609 2868 1612
rect 2867 1609 2877 1610
rect 2877 1609 2878 1618
rect 2866 1618 2878 1619
rect 2866 1618 2867 1620
rect 3611 1474 3612 1513
rect 3142 1474 3612 1475
rect 3142 1474 3143 1476
rect 3592 1575 3593 1585
rect 3425 1575 3593 1576
rect 3425 1555 3426 1576
rect 3190 1555 3426 1556
rect 3190 1528 3191 1556
rect 3190 1528 3570 1529
rect 3570 1528 3571 1546
rect 3570 1546 3724 1547
rect 3724 1546 3725 1618
rect 3724 1618 3735 1619
rect 3735 1618 3736 1620
rect 3608 1618 3609 1621
rect 3138 1618 3609 1619
rect 3138 1483 3139 1619
rect 3136 1483 3139 1484
rect 3136 1465 3137 1484
rect 3136 1465 3745 1466
rect 3745 1465 3746 1501
rect 3745 1501 3752 1502
rect 3752 1501 3753 1537
rect 3752 1537 3760 1538
rect 3760 1537 3761 1573
rect 3760 1573 3770 1574
rect 3770 1573 3771 1611
rect 3033 1537 3034 1540
rect 3028 1537 3034 1538
rect 3028 1537 3029 1555
rect 3025 1555 3029 1556
rect 3025 1553 3026 1556
rect 2966 1429 2967 1432
rect 2966 1429 3090 1430
rect 3090 1429 3091 1467
rect 2896 1501 2897 1504
rect 2884 1501 2897 1502
rect 2884 1492 2885 1502
rect 2884 1492 2894 1493
rect 2894 1492 2895 1494
rect 3792 1537 3793 1540
rect 3762 1537 3793 1538
rect 3762 1492 3763 1538
rect 3754 1492 3763 1493
rect 3754 1465 3755 1493
rect 3747 1465 3755 1466
rect 3747 1456 3748 1466
rect 3134 1456 3748 1457
rect 3134 1456 3135 1501
rect 3134 1501 3136 1502
rect 3136 1501 3137 1573
rect 3092 1573 3137 1574
rect 3092 1573 3093 1575
rect 3883 1582 3884 1585
rect 3876 1582 3884 1583
rect 3876 1582 3877 1584
rect 3540 1636 3541 1639
rect 3009 1636 3541 1637
rect 3009 1636 3010 1663
rect 2996 1663 3010 1664
rect 2996 1663 2997 1672
rect 2984 1672 2997 1673
rect 2984 1654 2985 1673
rect 2976 1654 2985 1655
rect 2976 1627 2977 1655
rect 2976 1627 3005 1628
rect 3005 1609 3006 1628
rect 3005 1609 3129 1610
rect 3129 1600 3130 1610
rect 3129 1600 3132 1601
rect 3132 1600 3133 1602
rect 3022 1447 3023 1459
rect 2935 1447 3023 1448
rect 2935 1429 2936 1448
rect 2935 1429 2964 1430
rect 2964 1420 2965 1430
rect 2896 1420 2965 1421
rect 2896 1420 2897 1456
rect 2896 1456 2928 1457
rect 2928 1456 2929 1474
rect 2928 1474 2961 1475
rect 2961 1474 2962 1483
rect 2941 1483 2962 1484
rect 2941 1483 2942 1492
rect 2941 1492 2948 1493
rect 2948 1492 2949 1501
rect 2948 1501 2987 1502
rect 2987 1501 2988 1503
rect 2925 1600 2926 1603
rect 2925 1600 2958 1601
rect 2958 1600 2959 1620
rect 3763 1465 3764 1477
rect 3763 1465 3776 1466
rect 3776 1454 3777 1466
rect 3776 1454 3963 1455
rect 3963 1454 3964 1528
rect 3867 1528 3964 1529
rect 3867 1519 3868 1529
rect 3867 1519 3876 1520
rect 3876 1501 3877 1520
rect 3841 1501 3877 1502
rect 3841 1492 3842 1502
rect 3841 1492 3844 1493
rect 3844 1492 3845 1494
rect 3815 1546 3816 1549
rect 3815 1546 3866 1547
rect 3866 1546 3867 1555
rect 3843 1555 3867 1556
rect 3843 1555 3844 1557
rect 2860 1573 2861 1576
rect 2860 1573 2870 1574
rect 2870 1564 2871 1574
rect 2867 1564 2871 1565
rect 2867 1564 2868 1566
rect 3251 1663 3252 1675
rect 3251 1663 3283 1664
rect 3283 1663 3284 1665
rect 2941 1438 2942 1441
rect 2941 1438 2948 1439
rect 2948 1436 2949 1439
rect 3117 1580 3118 1603
rect 3095 1580 3118 1581
rect 3095 1580 3096 1591
rect 2965 1591 3096 1592
rect 2965 1591 2966 1620
rect 3502 1654 3503 1657
rect 3099 1654 3503 1655
rect 3099 1654 3100 1663
rect 3091 1663 3100 1664
rect 3091 1663 3092 1665
rect 3325 1663 3326 1666
rect 3325 1663 3575 1664
rect 3575 1645 3576 1664
rect 3575 1645 3648 1646
rect 3648 1645 3649 1647
rect 2860 1519 2861 1567
rect 2860 1519 2893 1520
rect 2893 1519 2894 1521
rect 3867 1564 3868 1567
rect 3867 1564 3874 1565
rect 3874 1564 3875 1566
rect 3479 1429 3480 1432
rect 3469 1429 3480 1430
rect 3469 1429 3470 1438
rect 3469 1438 3559 1439
rect 3559 1438 3560 1440
rect 2907 1555 2908 1558
rect 2890 1555 2908 1556
rect 2890 1555 2891 1564
rect 2890 1564 2897 1565
rect 2897 1564 2898 1566
rect 2984 1600 2985 1603
rect 2968 1600 2985 1601
rect 2968 1600 2969 1627
rect 2896 1627 2969 1628
rect 2896 1618 2897 1628
rect 2896 1618 2954 1619
rect 2954 1616 2955 1619
rect 3764 1627 3765 1630
rect 3764 1627 3824 1628
rect 3824 1609 3825 1628
rect 3811 1609 3825 1610
rect 3811 1609 3812 1611
rect 3599 1654 3600 1657
rect 3599 1654 3669 1655
rect 3669 1645 3670 1655
rect 3669 1645 3679 1646
rect 3679 1645 3680 1647
rect 2924 1465 2925 1468
rect 2914 1465 2925 1466
rect 2914 1465 2915 1467
rect 3808 1600 3809 1603
rect 3808 1600 3850 1601
rect 3850 1600 3851 1602
rect 3652 1447 3653 1450
rect 3198 1447 3653 1448
rect 3198 1429 3199 1448
rect 3195 1429 3199 1430
rect 3195 1429 3196 1431
rect 3577 1438 3578 1441
rect 3577 1438 3659 1439
rect 3659 1438 3660 1449
rect 2955 1591 2956 1594
rect 2884 1591 2956 1592
rect 2884 1591 2885 1681
rect 2884 1681 3073 1682
rect 3073 1672 3074 1682
rect 3073 1672 3076 1673
rect 3076 1672 3077 1674
rect 2930 1546 2931 1549
rect 2916 1546 2931 1547
rect 2916 1546 2917 1548
rect 3859 1591 3860 1594
rect 3859 1591 3910 1592
rect 3910 1582 3911 1592
rect 3904 1582 3911 1583
rect 3904 1582 3905 1584
rect 2986 1546 2987 1549
rect 2980 1546 2987 1547
rect 2980 1546 2981 1582
rect 2882 1582 2981 1583
rect 2882 1582 2883 1690
rect 2882 1690 3076 1691
rect 3076 1681 3077 1691
rect 3076 1681 3089 1682
rect 3089 1681 3090 1683
rect 2803 1627 2804 1630
rect 2803 1627 2810 1628
rect 2810 1627 2811 1629
rect 3769 1546 3770 1549
rect 3763 1546 3770 1547
rect 3763 1546 3764 1564
rect 3763 1564 3773 1565
rect 3773 1564 3774 1566
rect 3847 1456 3848 1459
rect 3847 1456 3857 1457
rect 3857 1456 3858 1465
rect 3825 1465 3858 1466
rect 3825 1465 3826 1476
rect 3953 1501 3954 1504
rect 3946 1501 3954 1502
rect 3946 1501 3947 1503
rect 3656 1636 3657 1639
rect 3613 1636 3657 1637
rect 3613 1636 3614 1638
rect 2825 1654 2826 1657
rect 2815 1654 2826 1655
rect 2815 1654 2816 1656
rect 3566 1654 3567 1657
rect 3503 1654 3567 1655
rect 3503 1652 3504 1655
rect 3085 1652 3504 1653
rect 3085 1652 3086 1679
rect 3085 1679 3094 1680
rect 3094 1679 3095 1681
rect 3094 1681 3298 1682
rect 3298 1672 3299 1682
rect 3298 1672 3308 1673
rect 3308 1672 3309 1674
rect 3836 1474 3837 1477
rect 3829 1474 3837 1475
rect 3829 1474 3830 1476
rect 3005 1456 3006 1459
rect 3002 1456 3006 1457
rect 3002 1456 3003 1465
rect 3002 1465 3084 1466
rect 3084 1465 3085 1474
rect 3084 1474 3093 1475
rect 3093 1411 3094 1475
rect 2972 1411 3094 1412
rect 2972 1411 2973 1413
rect 3058 1474 3059 1477
rect 3058 1474 3083 1475
rect 3083 1474 3084 1476
rect 3083 1476 3132 1477
rect 3132 1420 3133 1477
rect 3132 1420 3142 1421
rect 3142 1420 3143 1422
rect 2940 1510 2941 1513
rect 2940 1510 2950 1511
rect 2950 1510 2951 1521
rect 2875 1463 2876 1468
rect 3871 1537 3872 1540
rect 3871 1537 3891 1538
rect 3891 1537 3892 1562
rect 3863 1562 3892 1563
rect 3863 1562 3864 1564
rect 3818 1564 3864 1565
rect 3818 1564 3819 1566
rect 3787 1609 3788 1612
rect 3783 1609 3788 1610
rect 3783 1591 3784 1610
rect 3783 1591 3842 1592
rect 3842 1591 3843 1593
rect 2815 1636 2816 1639
rect 2815 1636 2822 1637
rect 2822 1636 2823 1638
rect 3457 1670 3458 1681
rect 3331 1681 3458 1682
rect 3331 1679 3332 1682
rect 3514 1429 3515 1432
rect 3510 1429 3515 1430
rect 3510 1429 3511 1431
rect 2816 1447 2817 1450
rect 2809 1447 2817 1448
rect 2809 1447 2810 1449
rect 3802 1573 3803 1576
rect 3790 1573 3803 1574
rect 3790 1573 3791 1582
rect 3777 1582 3791 1583
rect 3777 1582 3778 1593
rect 2941 1654 2942 1657
rect 2941 1654 2952 1655
rect 2952 1645 2953 1655
rect 2949 1645 2953 1646
rect 2949 1645 2950 1647
rect 3804 1474 3805 1477
rect 3801 1474 3805 1475
rect 3801 1474 3802 1476
rect 3524 1429 3525 1432
rect 3524 1429 3965 1430
rect 3965 1429 3966 1636
rect 3680 1636 3966 1637
rect 3680 1636 3681 1638
rect 3714 1618 3715 1621
rect 3644 1618 3715 1619
rect 3644 1618 3645 1620
<< metal2 >>
rect 3895 1465 3896 1468
rect 3895 1465 3925 1466
rect 3925 1465 3926 1483
rect 3896 1483 3926 1484
rect 3896 1483 3897 1485
rect 3857 1483 3858 1486
rect 3778 1483 3858 1484
rect 3778 1483 3779 1485
rect 2992 1618 2993 1621
rect 2992 1618 3034 1619
rect 3034 1618 3035 1645
rect 3034 1645 3049 1646
rect 3049 1645 3050 1647
rect 2920 1474 2921 1477
rect 2920 1474 2929 1475
rect 2929 1456 2930 1475
rect 2929 1456 2935 1457
rect 2935 1456 2936 1458
rect 2994 1429 2995 1432
rect 2994 1429 3000 1430
rect 3000 1429 3001 1438
rect 2973 1438 3001 1439
rect 2973 1438 2974 1440
rect 3731 1573 3732 1576
rect 3684 1573 3732 1574
rect 3684 1555 3685 1574
rect 3681 1555 3685 1556
rect 3681 1555 3682 1557
rect 3566 1618 3567 1621
rect 3325 1618 3567 1619
rect 3325 1618 3326 1663
rect 3318 1663 3326 1664
rect 3318 1663 3319 1674
rect 2935 1483 2936 1486
rect 2910 1483 2936 1484
rect 2910 1483 2911 1485
rect 2945 1555 2946 1558
rect 2945 1555 2957 1556
rect 2957 1546 2958 1556
rect 2957 1546 2960 1547
rect 2960 1537 2961 1547
rect 2957 1537 2961 1538
rect 2957 1537 2958 1539
rect 3072 1429 3073 1432
rect 3002 1429 3073 1430
rect 3002 1429 3003 1447
rect 2981 1447 3003 1448
rect 2981 1447 2982 1449
rect 3794 1553 3795 1555
rect 3794 1555 3850 1556
rect 3850 1553 3851 1556
rect 3735 1591 3736 1594
rect 3708 1591 3736 1592
rect 3708 1591 3709 1593
rect 2938 1438 2939 1441
rect 2935 1438 2939 1439
rect 2935 1438 2936 1447
rect 2935 1447 2939 1448
rect 2939 1447 2940 1449
rect 3790 1528 3791 1531
rect 3741 1528 3791 1529
rect 3741 1528 3742 1600
rect 3693 1600 3742 1601
rect 3693 1600 3694 1602
rect 2910 1519 2911 1522
rect 2910 1519 2929 1520
rect 2929 1519 2930 1521
rect 3656 1609 3657 1612
rect 3656 1609 3783 1610
rect 3783 1591 3784 1610
rect 3783 1591 3793 1592
rect 3793 1573 3794 1592
rect 3793 1573 3820 1574
rect 3820 1573 3821 1575
rect 3705 1575 3706 1594
rect 3425 1575 3706 1576
rect 3425 1492 3426 1576
rect 3084 1492 3426 1493
rect 3084 1492 3085 1494
rect 2910 1465 2911 1468
rect 2890 1465 2911 1466
rect 2890 1465 2891 1492
rect 2890 1492 2917 1493
rect 2917 1492 2918 1510
rect 2917 1510 2933 1511
rect 2933 1510 2934 1512
rect 2934 1474 2935 1477
rect 2934 1474 2964 1475
rect 2964 1474 2965 1483
rect 2964 1483 2971 1484
rect 2971 1483 2972 1510
rect 2960 1510 2972 1511
rect 2960 1510 2961 1528
rect 2884 1528 2961 1529
rect 2884 1420 2885 1529
rect 2884 1420 2918 1421
rect 2918 1420 2919 1422
rect 3821 1519 3822 1522
rect 3821 1519 3825 1520
rect 3825 1501 3826 1520
rect 3825 1501 3872 1502
rect 3872 1501 3873 1503
rect 3905 1501 3906 1504
rect 3875 1501 3906 1502
rect 3875 1501 3876 1510
rect 3866 1510 3876 1511
rect 3866 1510 3867 1512
rect 3021 1528 3022 1540
rect 2981 1528 3022 1529
rect 2981 1528 2982 1530
rect 2909 1429 2910 1432
rect 2909 1429 2988 1430
rect 2988 1420 2989 1430
rect 2988 1420 3078 1421
rect 3078 1420 3079 1456
rect 2956 1456 3079 1457
rect 2956 1456 2957 1458
rect 2997 1636 2998 1639
rect 2997 1636 3032 1637
rect 3032 1636 3033 1654
rect 3032 1654 3316 1655
rect 3316 1616 3317 1655
rect 3316 1616 3578 1617
rect 3578 1616 3579 1629
rect 3623 1636 3624 1657
rect 3623 1636 3910 1637
rect 3910 1537 3911 1637
rect 3793 1537 3911 1538
rect 3793 1492 3794 1538
rect 3541 1492 3794 1493
rect 3541 1429 3542 1493
rect 3475 1429 3542 1430
rect 3475 1429 3476 1431
rect 3114 1600 3115 1603
rect 3027 1600 3115 1601
rect 3027 1600 3028 1602
rect 3124 1429 3125 1486
rect 3124 1429 3473 1430
rect 3473 1427 3474 1430
rect 3473 1427 3748 1428
rect 3748 1427 3749 1485
rect 3429 1663 3430 1666
rect 3355 1663 3430 1664
rect 3355 1663 3356 1681
rect 2944 1681 3356 1682
rect 2944 1672 2945 1682
rect 2934 1672 2945 1673
rect 2934 1672 2935 1674
rect 2983 1510 2984 1513
rect 2983 1510 3019 1511
rect 3019 1510 3020 1521
rect 3101 1627 3102 1630
rect 3043 1627 3102 1628
rect 3043 1618 3044 1628
rect 3037 1618 3044 1619
rect 3037 1618 3038 1620
rect 2970 1474 2971 1477
rect 2970 1474 2987 1475
rect 2987 1474 2988 1483
rect 2974 1483 2988 1484
rect 2974 1483 2975 1501
rect 2974 1501 2980 1502
rect 2980 1501 2981 1503
rect 3861 1519 3862 1522
rect 3861 1519 3963 1520
rect 3963 1463 3964 1520
rect 3871 1463 3964 1464
rect 3871 1463 3872 1467
rect 3854 1492 3855 1495
rect 3854 1492 3863 1493
rect 3863 1474 3864 1493
rect 3797 1474 3864 1475
rect 3797 1474 3798 1476
rect 2958 1564 2959 1567
rect 2958 1564 2962 1565
rect 2962 1564 2963 1618
rect 2962 1618 2968 1619
rect 2968 1618 2969 1636
rect 2952 1636 2969 1637
rect 2952 1636 2953 1654
rect 2951 1654 2953 1655
rect 2951 1654 2952 1663
rect 2946 1663 2952 1664
rect 2946 1663 2947 1665
rect 3104 1609 3105 1639
rect 2984 1609 3105 1610
rect 2984 1609 2985 1645
rect 2984 1645 3027 1646
rect 3027 1645 3028 1672
rect 3027 1672 3067 1673
rect 3067 1672 3068 1674
rect 3569 1618 3570 1621
rect 3569 1618 3575 1619
rect 3575 1618 3576 1636
rect 3575 1636 3598 1637
rect 3598 1618 3599 1637
rect 3594 1618 3599 1619
rect 3594 1609 3595 1619
rect 3594 1609 3597 1610
rect 3597 1609 3598 1611
rect 3259 1420 3260 1423
rect 3184 1420 3260 1421
rect 3184 1420 3185 1422
rect 3837 1582 3838 1585
rect 3824 1582 3838 1583
rect 3824 1582 3825 1591
rect 3824 1591 3863 1592
rect 3863 1591 3864 1627
rect 3701 1627 3864 1628
rect 3701 1627 3702 1629
rect 3860 1461 3861 1468
rect 3860 1461 3965 1462
rect 3965 1461 3966 1528
rect 3844 1528 3966 1529
rect 3844 1528 3845 1530
rect 2943 1537 2944 1540
rect 2882 1537 2944 1538
rect 2882 1411 2883 1538
rect 2882 1411 3087 1412
rect 3087 1411 3088 1465
rect 3034 1465 3088 1466
rect 3034 1465 3035 1537
rect 3027 1537 3035 1538
rect 3027 1537 3028 1546
rect 2975 1546 3028 1547
rect 2975 1519 2976 1547
rect 2975 1519 2991 1520
rect 2991 1519 2992 1521
rect 3496 1519 3497 1522
rect 3496 1519 3695 1520
rect 3695 1519 3696 1521
rect 3387 1501 3388 1513
rect 3057 1501 3388 1502
rect 3057 1492 3058 1502
rect 3051 1492 3058 1493
rect 3051 1492 3052 1494
rect 2964 1555 2965 1558
rect 2964 1555 3042 1556
rect 3042 1510 3043 1556
rect 3042 1510 3048 1511
rect 3048 1483 3049 1511
rect 3048 1483 3093 1484
rect 3093 1409 3094 1484
rect 2872 1409 3094 1410
rect 2872 1409 2873 1573
rect 2872 1573 2878 1574
rect 2878 1573 2879 1575
rect 3721 1618 3722 1621
rect 3600 1618 3722 1619
rect 3600 1618 3601 1654
rect 3575 1654 3601 1655
rect 3575 1654 3576 1663
rect 3575 1663 3654 1664
rect 3654 1645 3655 1664
rect 3651 1645 3655 1646
rect 3651 1645 3652 1647
rect 3698 1519 3699 1522
rect 3698 1519 3779 1520
rect 3779 1519 3780 1521
rect 2954 1420 2955 1423
rect 2954 1420 2961 1421
rect 2961 1420 2962 1422
rect 2948 1591 2949 1594
rect 2948 1591 2960 1592
rect 2960 1573 2961 1592
rect 2946 1573 2961 1574
rect 2946 1573 2947 1575
rect 2941 1600 2942 1603
rect 2909 1600 2942 1601
rect 2909 1600 2910 1602
rect 2910 1609 2911 1612
rect 2896 1609 2911 1610
rect 2896 1591 2897 1610
rect 2896 1591 2924 1592
rect 2924 1591 2925 1593
rect 2899 1627 2900 1657
rect 2899 1627 2922 1628
rect 2922 1627 2923 1629
rect 3352 1654 3353 1666
rect 3352 1654 3562 1655
rect 3562 1654 3563 1656
rect 2971 1465 2972 1468
rect 2964 1465 2972 1466
rect 2964 1465 2965 1467
rect 3055 1528 3056 1594
rect 3055 1528 3121 1529
rect 3121 1528 3122 1530
rect 2937 1609 2938 1612
rect 2937 1609 2957 1610
rect 2957 1609 2958 1618
rect 2937 1618 2958 1619
rect 2937 1618 2938 1620
rect 3889 1483 3890 1486
rect 3872 1483 3890 1484
rect 3872 1483 3873 1494
rect 3857 1420 3858 1468
rect 3276 1420 3858 1421
rect 3276 1420 3277 1422
rect 3780 1573 3781 1576
rect 3765 1573 3781 1574
rect 3765 1573 3766 1582
rect 3757 1582 3766 1583
rect 3757 1582 3758 1584
rect 2928 1555 2929 1558
rect 2924 1555 2929 1556
rect 2924 1555 2925 1557
rect 2984 1492 2985 1495
rect 2984 1492 2998 1493
rect 2998 1465 2999 1493
rect 2998 1465 3011 1466
rect 3011 1465 3012 1467
rect 2928 1645 2929 1648
rect 2908 1645 2929 1646
rect 2908 1636 2909 1646
rect 2908 1636 2932 1637
rect 2932 1636 2933 1638
rect 3856 1546 3857 1549
rect 3856 1546 3889 1547
rect 3889 1546 3890 1582
rect 3848 1582 3890 1583
rect 3848 1582 3849 1584
rect 3529 1447 3530 1450
rect 3529 1447 3539 1448
rect 3539 1447 3540 1510
rect 3539 1510 3779 1511
rect 3779 1510 3780 1512
rect 3132 1609 3133 1612
rect 3120 1609 3133 1610
rect 3120 1582 3121 1610
rect 3076 1582 3121 1583
rect 3076 1582 3077 1584
rect 3542 1645 3543 1648
rect 3542 1645 3572 1646
rect 3572 1645 3573 1690
rect 2992 1690 3573 1691
rect 2992 1690 2993 1692
<< end >>
