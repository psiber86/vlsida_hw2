magic
tech scmos
timestamp 1395743126
<< m1p >>
use CELL  1
transform -1 0 2477 0 1 2481
box 0 0 6 6
use CELL  2
transform 1 0 2587 0 1 2076
box 0 0 6 6
use CELL  3
transform 1 0 2369 0 1 2076
box 0 0 6 6
use CELL  4
transform -1 0 2572 0 -1 3503
box 0 0 6 6
use CELL  5
transform -1 0 2796 0 -1 2487
box 0 0 6 6
use CELL  6
transform 1 0 2362 0 1 2076
box 0 0 6 6
use CELL  7
transform -1 0 2467 0 1 3458
box 0 0 6 6
use CELL  8
transform 1 0 2819 0 1 2600
box 0 0 6 6
use CELL  9
transform -1 0 2350 0 1 3458
box 0 0 6 6
use CELL  10
transform -1 0 2807 0 1 1826
box 0 0 6 6
use CELL  11
transform -1 0 2306 0 1 2600
box 0 0 6 6
use CELL  12
transform -1 0 2386 0 1 1432
box 0 0 6 6
use CELL  13
transform -1 0 2464 0 1 1513
box 0 0 6 6
use CELL  14
transform -1 0 2521 0 1 1717
box 0 0 6 6
use CELL  15
transform 1 0 2468 0 1 2870
box 0 0 6 6
use CELL  16
transform 1 0 2477 0 1 3306
box 0 0 6 6
use CELL  17
transform 1 0 2742 0 1 2971
box 0 0 6 6
use CELL  18
transform -1 0 2400 0 1 1235
box 0 0 6 6
use CELL  19
transform -1 0 2359 0 1 2199
box 0 0 6 6
use CELL  20
transform 1 0 2512 0 -1 1519
box 0 0 6 6
use CELL  21
transform 1 0 2356 0 -1 2348
box 0 0 6 6
use CELL  22
transform 1 0 2552 0 1 3100
box 0 0 6 6
use CELL  23
transform 1 0 2862 0 -1 2205
box 0 0 6 6
use CELL  24
transform -1 0 2590 0 1 1513
box 0 0 6 6
use CELL  25
transform 1 0 2401 0 1 3541
box 0 0 6 6
use CELL  26
transform -1 0 2322 0 1 3100
box 0 0 6 6
use CELL  27
transform -1 0 2607 0 -1 1438
box 0 0 6 6
use CELL  28
transform -1 0 2328 0 -1 2082
box 0 0 6 6
use CELL  29
transform -1 0 2707 0 1 1717
box 0 0 6 6
use CELL  30
transform 1 0 2847 0 1 2600
box 0 0 6 6
use CELL  31
transform 1 0 2668 0 1 3100
box 0 0 6 6
use CELL  32
transform 1 0 2580 0 1 3458
box 0 0 6 6
use CELL  33
transform 1 0 2389 0 1 2870
box 0 0 6 6
use CELL  34
transform -1 0 2325 0 1 2600
box 0 0 6 6
use CELL  35
transform 1 0 2473 0 -1 1157
box 0 0 6 6
use CELL  36
transform -1 0 2626 0 1 3306
box 0 0 6 6
use CELL  37
transform -1 0 2466 0 1 1365
box 0 0 6 6
use CELL  38
transform -1 0 2613 0 -1 3195
box 0 0 6 6
use CELL  39
transform -1 0 2482 0 1 1290
box 0 0 6 6
use CELL  40
transform 1 0 2761 0 -1 2348
box 0 0 6 6
use CELL  41
transform -1 0 2659 0 -1 1723
box 0 0 6 6
use CELL  42
transform 1 0 2708 0 1 3100
box 0 0 6 6
use CELL  43
transform 1 0 2706 0 1 2342
box 0 0 6 6
use CELL  44
transform 1 0 2642 0 1 3100
box 0 0 6 6
use CELL  45
transform -1 0 2413 0 1 1432
box 0 0 6 6
use CELL  46
transform 1 0 2642 0 -1 2876
box 0 0 6 6
use CELL  47
transform 1 0 2652 0 1 1290
box 0 0 6 6
use CELL  48
transform -1 0 2325 0 -1 1832
box 0 0 6 6
use CELL  49
transform 1 0 2719 0 1 3189
box 0 0 6 6
use CELL  50
transform -1 0 2311 0 1 3189
box 0 0 6 6
use CELL  51
transform 1 0 2364 0 1 2745
box 0 0 6 6
use CELL  52
transform 1 0 2342 0 -1 1519
box 0 0 6 6
use CELL  53
transform -1 0 2372 0 1 1365
box 0 0 6 6
use CELL  54
transform 1 0 2327 0 1 3306
box 0 0 6 6
use CELL  55
transform 1 0 2665 0 1 3306
box 0 0 6 6
use CELL  56
transform -1 0 2362 0 -1 1519
box 0 0 6 6
use CELL  57
transform 1 0 2825 0 1 2481
box 0 0 6 6
use CELL  58
transform -1 0 2678 0 1 3306
box 0 0 6 6
use CELL  59
transform -1 0 2336 0 1 3458
box 0 0 6 6
use CELL  60
transform 1 0 2855 0 1 2199
box 0 0 6 6
use CELL  61
transform -1 0 2623 0 -1 3395
box 0 0 6 6
use CELL  62
transform 1 0 2680 0 -1 1519
box 0 0 6 6
use CELL  63
transform -1 0 2809 0 1 2342
box 0 0 6 6
use CELL  64
transform 1 0 2796 0 -1 2348
box 0 0 6 6
use CELL  65
transform -1 0 2453 0 1 3541
box 0 0 6 6
use CELL  66
transform 1 0 2350 0 -1 1438
box 0 0 6 6
use CELL  67
transform -1 0 2344 0 1 1290
box 0 0 6 6
use CELL  68
transform 1 0 2396 0 1 2870
box 0 0 6 6
use CELL  69
transform 1 0 2624 0 1 3389
box 0 0 6 6
use CELL  70
transform 1 0 2624 0 -1 2977
box 0 0 6 6
use CELL  71
transform 1 0 2286 0 -1 2606
box 0 0 6 6
use CELL  72
transform 1 0 2450 0 1 1151
box 0 0 6 6
use CELL  73
transform 1 0 2329 0 1 3497
box 0 0 6 6
use CELL  74
transform -1 0 2304 0 1 3306
box 0 0 6 6
use CELL  75
transform 1 0 2328 0 1 3518
box 0 0 6 6
use CELL  76
transform 1 0 2349 0 -1 1519
box 0 0 6 6
use CELL  77
transform 1 0 2335 0 1 3518
box 0 0 6 6
use CELL  78
transform 1 0 2342 0 1 3518
box 0 0 6 6
use CELL  79
transform -1 0 2403 0 1 3306
box 0 0 6 6
use CELL  80
transform -1 0 2745 0 1 1717
box 0 0 6 6
use CELL  81
transform 1 0 2349 0 1 3518
box 0 0 6 6
use CELL  82
transform 1 0 2725 0 -1 1723
box 0 0 6 6
use CELL  83
transform 1 0 2329 0 1 2076
box 0 0 6 6
use CELL  84
transform -1 0 2528 0 1 3497
box 0 0 6 6
use CELL  85
transform -1 0 2832 0 1 2600
box 0 0 6 6
use CELL  86
transform -1 0 2339 0 -1 1832
box 0 0 6 6
use CELL  87
transform -1 0 2715 0 -1 2977
box 0 0 6 6
use CELL  88
transform 1 0 2555 0 1 2870
box 0 0 6 6
use CELL  89
transform -1 0 2474 0 1 1941
box 0 0 6 6
use CELL  90
transform 1 0 2323 0 1 1941
box 0 0 6 6
use CELL  91
transform 1 0 2364 0 -1 2606
box 0 0 6 6
use CELL  92
transform 1 0 2395 0 1 2600
box 0 0 6 6
use CELL  93
transform 1 0 2711 0 1 1622
box 0 0 6 6
use CELL  94
transform -1 0 2324 0 1 2481
box 0 0 6 6
use CELL  95
transform 1 0 2716 0 -1 2751
box 0 0 6 6
use CELL  96
transform 1 0 2570 0 1 1365
box 0 0 6 6
use CELL  97
transform 1 0 2545 0 1 3306
box 0 0 6 6
use CELL  98
transform -1 0 2744 0 -1 2205
box 0 0 6 6
use CELL  99
transform 1 0 2308 0 -1 2348
box 0 0 6 6
use CELL  100
transform -1 0 2411 0 1 3189
box 0 0 6 6
use CELL  101
transform -1 0 2382 0 -1 3547
box 0 0 6 6
use CELL  102
transform 1 0 2646 0 1 3189
box 0 0 6 6
use CELL  103
transform 1 0 2732 0 1 1717
box 0 0 6 6
use CELL  104
transform 1 0 2457 0 -1 1157
box 0 0 6 6
use CELL  105
transform -1 0 2640 0 1 1365
box 0 0 6 6
use CELL  106
transform -1 0 2356 0 1 2076
box 0 0 6 6
use CELL  107
transform -1 0 2677 0 1 1290
box 0 0 6 6
use CELL  108
transform 1 0 2385 0 1 2745
box 0 0 6 6
use CELL  109
transform 1 0 2738 0 -1 2487
box 0 0 6 6
use CELL  110
transform -1 0 2298 0 1 2870
box 0 0 6 6
use CELL  111
transform -1 0 2377 0 1 2745
box 0 0 6 6
use CELL  112
transform -1 0 2376 0 1 2971
box 0 0 6 6
use CELL  113
transform -1 0 2881 0 1 2199
box 0 0 6 6
use CELL  114
transform -1 0 2729 0 1 2745
box 0 0 6 6
use CELL  115
transform -1 0 2388 0 -1 2876
box 0 0 6 6
use CELL  116
transform 1 0 2632 0 1 3306
box 0 0 6 6
use CELL  117
transform -1 0 2330 0 -1 3195
box 0 0 6 6
use CELL  118
transform 1 0 2639 0 1 3306
box 0 0 6 6
use CELL  119
transform 1 0 2286 0 1 3458
box 0 0 6 6
use CELL  120
transform -1 0 2796 0 -1 2205
box 0 0 6 6
use CELL  121
transform 1 0 2280 0 1 2342
box 0 0 6 6
use CELL  122
transform -1 0 2518 0 1 1365
box 0 0 6 6
use CELL  123
transform -1 0 2379 0 1 1622
box 0 0 6 6
use CELL  124
transform -1 0 2753 0 1 1622
box 0 0 6 6
use CELL  125
transform 1 0 2385 0 1 3306
box 0 0 6 6
use CELL  126
transform 1 0 2364 0 -1 1157
box 0 0 6 6
use CELL  127
transform -1 0 2399 0 1 2481
box 0 0 6 6
use CELL  128
transform 1 0 2552 0 1 2971
box 0 0 6 6
use CELL  129
transform 1 0 2811 0 1 2481
box 0 0 6 6
use CELL  130
transform 1 0 2350 0 1 1365
box 0 0 6 6
use CELL  131
transform 1 0 2378 0 1 1365
box 0 0 6 6
use CELL  132
transform 1 0 2390 0 1 1365
box 0 0 6 6
use CELL  133
transform 1 0 2527 0 1 1432
box 0 0 6 6
use CELL  134
transform 1 0 2394 0 1 3541
box 0 0 6 6
use CELL  135
transform 1 0 2453 0 1 1365
box 0 0 6 6
use CELL  136
transform 1 0 2716 0 -1 2977
box 0 0 6 6
use CELL  137
transform -1 0 2355 0 1 2342
box 0 0 6 6
use CELL  138
transform 1 0 2345 0 1 1622
box 0 0 6 6
use CELL  139
transform -1 0 2311 0 1 3306
box 0 0 6 6
use CELL  140
transform 1 0 2573 0 1 3458
box 0 0 6 6
use CELL  141
transform -1 0 2737 0 1 2199
box 0 0 6 6
use CELL  142
transform -1 0 2311 0 -1 1832
box 0 0 6 6
use CELL  143
transform -1 0 2705 0 1 3306
box 0 0 6 6
use CELL  144
transform 1 0 2692 0 -1 3312
box 0 0 6 6
use CELL  145
transform -1 0 2814 0 1 1826
box 0 0 6 6
use CELL  146
transform 1 0 2621 0 -1 1947
box 0 0 6 6
use CELL  147
transform -1 0 2318 0 1 2870
box 0 0 6 6
use CELL  148
transform 1 0 2510 0 1 2870
box 0 0 6 6
use CELL  149
transform -1 0 2377 0 1 1432
box 0 0 6 6
use CELL  150
transform 1 0 2423 0 1 2342
box 0 0 6 6
use CELL  151
transform 1 0 2313 0 -1 2977
box 0 0 6 6
use CELL  152
transform -1 0 2549 0 -1 3464
box 0 0 6 6
use CELL  153
transform 1 0 2566 0 1 1432
box 0 0 6 6
use CELL  154
transform 1 0 2843 0 1 1826
box 0 0 6 6
use CELL  155
transform 1 0 2768 0 -1 2348
box 0 0 6 6
use CELL  156
transform -1 0 2584 0 -1 1723
box 0 0 6 6
use CELL  157
transform 1 0 2472 0 -1 2751
box 0 0 6 6
use CELL  158
transform -1 0 2328 0 -1 1204
box 0 0 6 6
use CELL  159
transform 1 0 2573 0 1 1432
box 0 0 6 6
use CELL  160
transform -1 0 2576 0 -1 2348
box 0 0 6 6
use CELL  161
transform 1 0 2833 0 -1 2205
box 0 0 6 6
use CELL  162
transform 1 0 2374 0 1 2199
box 0 0 6 6
use CELL  163
transform -1 0 2732 0 1 3189
box 0 0 6 6
use CELL  164
transform 1 0 2339 0 -1 1723
box 0 0 6 6
use CELL  165
transform 1 0 2539 0 1 1365
box 0 0 6 6
use CELL  166
transform -1 0 2651 0 1 1290
box 0 0 6 6
use CELL  167
transform 1 0 2540 0 1 3389
box 0 0 6 6
use CELL  168
transform 1 0 2778 0 1 2600
box 0 0 6 6
use CELL  169
transform 1 0 2768 0 1 2745
box 0 0 6 6
use CELL  170
transform 1 0 2673 0 1 1513
box 0 0 6 6
use CELL  171
transform -1 0 2311 0 1 2870
box 0 0 6 6
use CELL  172
transform 1 0 2543 0 1 3497
box 0 0 6 6
use CELL  173
transform 1 0 2375 0 1 2342
box 0 0 6 6
use CELL  174
transform 1 0 2360 0 1 1717
box 0 0 6 6
use CELL  175
transform 1 0 2336 0 1 1198
box 0 0 6 6
use CELL  176
transform 1 0 2329 0 1 1151
box 0 0 6 6
use CELL  177
transform 1 0 2726 0 -1 1628
box 0 0 6 6
use CELL  178
transform 1 0 2336 0 1 1151
box 0 0 6 6
use CELL  179
transform 1 0 2317 0 -1 3395
box 0 0 6 6
use CELL  180
transform 1 0 2443 0 1 1151
box 0 0 6 6
use CELL  181
transform 1 0 2528 0 1 3518
box 0 0 6 6
use CELL  182
transform 1 0 2521 0 1 3518
box 0 0 6 6
use CELL  183
transform 1 0 2761 0 1 2745
box 0 0 6 6
use CELL  184
transform 1 0 2500 0 1 3518
box 0 0 6 6
use CELL  185
transform -1 0 2423 0 -1 3395
box 0 0 6 6
use CELL  186
transform -1 0 2497 0 1 2745
box 0 0 6 6
use CELL  187
transform 1 0 2448 0 1 3518
box 0 0 6 6
use CELL  188
transform -1 0 2347 0 1 2481
box 0 0 6 6
use CELL  189
transform 1 0 2363 0 1 3518
box 0 0 6 6
use CELL  190
transform 1 0 2368 0 -1 1832
box 0 0 6 6
use CELL  191
transform 1 0 2518 0 1 1198
box 0 0 6 6
use CELL  192
transform 1 0 2377 0 1 3518
box 0 0 6 6
use CELL  193
transform -1 0 2657 0 -1 3312
box 0 0 6 6
use CELL  194
transform -1 0 2334 0 1 1513
box 0 0 6 6
use CELL  195
transform 1 0 2589 0 1 3189
box 0 0 6 6
use CELL  196
transform -1 0 2671 0 -1 2606
box 0 0 6 6
use CELL  197
transform 1 0 2630 0 1 2870
box 0 0 6 6
use CELL  198
transform -1 0 2367 0 -1 1832
box 0 0 6 6
use CELL  199
transform 1 0 2827 0 1 2076
box 0 0 6 6
use CELL  200
transform 1 0 2854 0 1 2600
box 0 0 6 6
use CELL  201
transform 1 0 2420 0 1 3518
box 0 0 6 6
use CELL  202
transform 1 0 2836 0 1 1826
box 0 0 6 6
use CELL  203
transform -1 0 2835 0 1 1826
box 0 0 6 6
use CELL  204
transform 1 0 2441 0 1 3518
box 0 0 6 6
use CELL  205
transform 1 0 2322 0 1 1432
box 0 0 6 6
use CELL  206
transform -1 0 2528 0 1 2481
box 0 0 6 6
use CELL  207
transform 1 0 2356 0 1 3518
box 0 0 6 6
use CELL  208
transform 1 0 2761 0 1 1622
box 0 0 6 6
use CELL  209
transform 1 0 2455 0 1 3518
box 0 0 6 6
use CELL  210
transform -1 0 2394 0 1 2076
box 0 0 6 6
use CELL  211
transform 1 0 2515 0 1 3458
box 0 0 6 6
use CELL  212
transform -1 0 2558 0 -1 3503
box 0 0 6 6
use CELL  213
transform -1 0 2358 0 1 1622
box 0 0 6 6
use CELL  214
transform -1 0 2298 0 1 2971
box 0 0 6 6
use CELL  215
transform -1 0 2521 0 1 1432
box 0 0 6 6
use CELL  216
transform -1 0 2395 0 1 3497
box 0 0 6 6
use CELL  217
transform 1 0 2754 0 -1 1628
box 0 0 6 6
use CELL  218
transform 1 0 2434 0 1 3518
box 0 0 6 6
use CELL  219
transform 1 0 2591 0 1 3100
box 0 0 6 6
use CELL  220
transform 1 0 2370 0 1 3518
box 0 0 6 6
use CELL  221
transform 1 0 2564 0 1 3458
box 0 0 6 6
use CELL  222
transform 1 0 2635 0 1 1432
box 0 0 6 6
use CELL  223
transform 1 0 2330 0 1 1941
box 0 0 6 6
use CELL  224
transform 1 0 2473 0 1 3518
box 0 0 6 6
use CELL  225
transform 1 0 2690 0 -1 2606
box 0 0 6 6
use CELL  226
transform -1 0 2719 0 1 2342
box 0 0 6 6
use CELL  227
transform -1 0 2743 0 -1 2348
box 0 0 6 6
use CELL  228
transform -1 0 2399 0 1 3518
box 0 0 6 6
use CELL  229
transform 1 0 2401 0 -1 3464
box 0 0 6 6
use CELL  230
transform 1 0 2441 0 1 1198
box 0 0 6 6
use CELL  231
transform 1 0 2800 0 -1 2606
box 0 0 6 6
use CELL  232
transform 1 0 2323 0 1 3458
box 0 0 6 6
use CELL  233
transform 1 0 2411 0 1 3518
box 0 0 6 6
use CELL  234
transform -1 0 2328 0 -1 3503
box 0 0 6 6
use CELL  235
transform 1 0 2842 0 1 2199
box 0 0 6 6
use CELL  236
transform 1 0 2705 0 -1 2487
box 0 0 6 6
use CELL  237
transform 1 0 2625 0 1 1365
box 0 0 6 6
use CELL  238
transform -1 0 2358 0 1 2600
box 0 0 6 6
use CELL  239
transform -1 0 2794 0 1 1622
box 0 0 6 6
use CELL  240
transform 1 0 2657 0 1 1432
box 0 0 6 6
use CELL  241
transform 1 0 2392 0 1 2971
box 0 0 6 6
use CELL  242
transform 1 0 2331 0 1 1622
box 0 0 6 6
use CELL  243
transform -1 0 2316 0 -1 3395
box 0 0 6 6
use CELL  244
transform -1 0 2490 0 -1 2751
box 0 0 6 6
use CELL  245
transform -1 0 2597 0 1 2971
box 0 0 6 6
use CELL  246
transform -1 0 2360 0 1 2870
box 0 0 6 6
use CELL  247
transform 1 0 2411 0 -1 3106
box 0 0 6 6
use CELL  248
transform -1 0 2446 0 1 3541
box 0 0 6 6
use CELL  249
transform -1 0 2477 0 -1 2977
box 0 0 6 6
use CELL  250
transform 1 0 2577 0 1 1365
box 0 0 6 6
use CELL  251
transform -1 0 2855 0 -1 2205
box 0 0 6 6
use CELL  252
transform 1 0 2332 0 1 1717
box 0 0 6 6
use CELL  253
transform 1 0 2760 0 1 1717
box 0 0 6 6
use CELL  254
transform 1 0 2495 0 1 2971
box 0 0 6 6
use CELL  255
transform -1 0 2332 0 1 1826
box 0 0 6 6
use CELL  256
transform 1 0 2611 0 1 1235
box 0 0 6 6
use CELL  257
transform 1 0 2834 0 1 2076
box 0 0 6 6
use CELL  258
transform -1 0 2564 0 -1 1296
box 0 0 6 6
use CELL  259
transform 1 0 2671 0 1 1432
box 0 0 6 6
use CELL  260
transform 1 0 2361 0 1 3497
box 0 0 6 6
use CELL  261
transform 1 0 2753 0 1 1717
box 0 0 6 6
use CELL  262
transform -1 0 2773 0 1 1717
box 0 0 6 6
use CELL  263
transform -1 0 2335 0 1 1432
box 0 0 6 6
use CELL  264
transform -1 0 2329 0 -1 1241
box 0 0 6 6
use CELL  265
transform 1 0 2293 0 -1 1519
box 0 0 6 6
use CELL  266
transform -1 0 2473 0 -1 1723
box 0 0 6 6
use CELL  267
transform 1 0 2314 0 1 2199
box 0 0 6 6
use CELL  268
transform 1 0 2539 0 1 1826
box 0 0 6 6
use CELL  269
transform -1 0 2821 0 -1 1947
box 0 0 6 6
use CELL  270
transform -1 0 2305 0 1 2870
box 0 0 6 6
use CELL  271
transform 1 0 2322 0 1 1151
box 0 0 6 6
use CELL  272
transform 1 0 2611 0 1 1365
box 0 0 6 6
use CELL  273
transform -1 0 2377 0 1 1151
box 0 0 6 6
use CELL  274
transform -1 0 2473 0 -1 1832
box 0 0 6 6
use CELL  275
transform 1 0 2350 0 1 1198
box 0 0 6 6
use CELL  276
transform 1 0 2364 0 1 1198
box 0 0 6 6
use CELL  277
transform -1 0 2821 0 1 1826
box 0 0 6 6
use CELL  278
transform 1 0 2358 0 1 1124
box 0 0 6 6
use CELL  279
transform 1 0 2378 0 1 1198
box 0 0 6 6
use CELL  280
transform 1 0 2399 0 1 1198
box 0 0 6 6
use CELL  281
transform -1 0 2364 0 -1 1947
box 0 0 6 6
use CELL  282
transform -1 0 2506 0 1 3458
box 0 0 6 6
use CELL  283
transform -1 0 2574 0 1 3189
box 0 0 6 6
use CELL  284
transform -1 0 2338 0 1 2199
box 0 0 6 6
use CELL  285
transform 1 0 2453 0 1 1198
box 0 0 6 6
use CELL  286
transform -1 0 2595 0 1 1432
box 0 0 6 6
use CELL  287
transform -1 0 2419 0 1 1717
box 0 0 6 6
use CELL  288
transform 1 0 2490 0 1 1198
box 0 0 6 6
use CELL  289
transform -1 0 2304 0 1 2076
box 0 0 6 6
use CELL  290
transform 1 0 2703 0 1 1941
box 0 0 6 6
use CELL  291
transform 1 0 2534 0 1 1198
box 0 0 6 6
use CELL  292
transform 1 0 2550 0 1 1198
box 0 0 6 6
use CELL  293
transform -1 0 2423 0 -1 3503
box 0 0 6 6
use CELL  294
transform 1 0 2454 0 1 3497
box 0 0 6 6
use CELL  295
transform -1 0 2788 0 -1 1628
box 0 0 6 6
use CELL  296
transform -1 0 2333 0 1 2745
box 0 0 6 6
use CELL  297
transform -1 0 2799 0 1 2600
box 0 0 6 6
use CELL  298
transform 1 0 2410 0 -1 2205
box 0 0 6 6
use CELL  299
transform -1 0 2356 0 -1 1157
box 0 0 6 6
use CELL  300
transform -1 0 2774 0 1 1622
box 0 0 6 6
use CELL  301
transform 1 0 2578 0 1 1198
box 0 0 6 6
use CELL  302
transform 1 0 2587 0 -1 3312
box 0 0 6 6
use CELL  303
transform 1 0 2507 0 1 3518
box 0 0 6 6
use CELL  304
transform -1 0 2522 0 1 2342
box 0 0 6 6
use CELL  305
transform -1 0 2374 0 1 2342
box 0 0 6 6
use CELL  306
transform 1 0 2535 0 1 3518
box 0 0 6 6
use CELL  307
transform 1 0 2426 0 1 1365
box 0 0 6 6
use CELL  308
transform 1 0 2563 0 1 1365
box 0 0 6 6
use CELL  309
transform -1 0 2317 0 1 1717
box 0 0 6 6
use CELL  310
transform 1 0 2749 0 1 2971
box 0 0 6 6
use CELL  311
transform 1 0 2623 0 1 2199
box 0 0 6 6
use CELL  312
transform 1 0 2682 0 1 3100
box 0 0 6 6
use CELL  313
transform 1 0 2359 0 1 3189
box 0 0 6 6
use CELL  314
transform 1 0 2286 0 1 2199
box 0 0 6 6
use CELL  315
transform 1 0 2346 0 -1 2205
box 0 0 6 6
use CELL  316
transform 1 0 2348 0 1 3306
box 0 0 6 6
use CELL  317
transform 1 0 2746 0 1 1941
box 0 0 6 6
use CELL  318
transform 1 0 2364 0 1 3389
box 0 0 6 6
use CELL  319
transform -1 0 2875 0 -1 2205
box 0 0 6 6
use CELL  320
transform 1 0 2394 0 1 3389
box 0 0 6 6
use CELL  321
transform -1 0 2812 0 -1 2082
box 0 0 6 6
use CELL  322
transform 1 0 2480 0 1 1151
box 0 0 6 6
use CELL  323
transform -1 0 2380 0 1 1717
box 0 0 6 6
use CELL  324
transform 1 0 2709 0 1 2745
box 0 0 6 6
use CELL  325
transform 1 0 2410 0 1 1622
box 0 0 6 6
use CELL  326
transform 1 0 2307 0 1 2199
box 0 0 6 6
use CELL  327
transform -1 0 2323 0 -1 3195
box 0 0 6 6
use CELL  328
transform 1 0 2531 0 1 3389
box 0 0 6 6
use CELL  329
transform -1 0 2533 0 -1 1204
box 0 0 6 6
use CELL  330
transform 1 0 2601 0 1 1622
box 0 0 6 6
use CELL  331
transform -1 0 2853 0 -1 2082
box 0 0 6 6
use CELL  332
transform 1 0 2524 0 1 2600
box 0 0 6 6
use CELL  333
transform -1 0 2381 0 -1 3503
box 0 0 6 6
use CELL  334
transform 1 0 2705 0 1 3189
box 0 0 6 6
use CELL  335
transform 1 0 2631 0 1 1622
box 0 0 6 6
use CELL  336
transform 1 0 2376 0 1 2600
box 0 0 6 6
use CELL  337
transform -1 0 2317 0 1 3306
box 0 0 6 6
use CELL  338
transform -1 0 2330 0 1 1622
box 0 0 6 6
use CELL  339
transform 1 0 2350 0 1 3389
box 0 0 6 6
use CELL  340
transform 1 0 2744 0 -1 2876
box 0 0 6 6
use CELL  341
transform 1 0 2610 0 1 3389
box 0 0 6 6
use CELL  342
transform 1 0 2358 0 1 3458
box 0 0 6 6
use CELL  343
transform 1 0 2550 0 1 1622
box 0 0 6 6
use CELL  344
transform 1 0 2675 0 1 3100
box 0 0 6 6
use CELL  345
transform -1 0 2503 0 1 1198
box 0 0 6 6
use CELL  346
transform 1 0 2644 0 -1 1723
box 0 0 6 6
use CELL  347
transform 1 0 2345 0 1 3189
box 0 0 6 6
use CELL  348
transform 1 0 2423 0 1 3458
box 0 0 6 6
use CELL  349
transform 1 0 2468 0 1 3458
box 0 0 6 6
use CELL  350
transform 1 0 2475 0 1 3458
box 0 0 6 6
use CELL  351
transform 1 0 2482 0 1 3458
box 0 0 6 6
use CELL  352
transform -1 0 2414 0 1 1151
box 0 0 6 6
use CELL  353
transform 1 0 2775 0 1 2971
box 0 0 6 6
use CELL  354
transform 1 0 2789 0 -1 2348
box 0 0 6 6
use CELL  355
transform 1 0 2797 0 1 2481
box 0 0 6 6
use CELL  356
transform -1 0 2784 0 1 2481
box 0 0 6 6
use CELL  357
transform 1 0 2341 0 1 3306
box 0 0 6 6
use CELL  358
transform 1 0 2398 0 1 3189
box 0 0 6 6
use CELL  359
transform 1 0 2667 0 -1 3195
box 0 0 6 6
use CELL  360
transform 1 0 2468 0 1 3389
box 0 0 6 6
use CELL  361
transform 1 0 2415 0 -1 1157
box 0 0 6 6
use CELL  362
transform 1 0 2524 0 1 3389
box 0 0 6 6
use CELL  363
transform -1 0 2464 0 -1 1628
box 0 0 6 6
use CELL  364
transform 1 0 2636 0 1 1513
box 0 0 6 6
use CELL  365
transform -1 0 2367 0 1 2870
box 0 0 6 6
use CELL  366
transform 1 0 2589 0 1 3389
box 0 0 6 6
use CELL  367
transform -1 0 2361 0 1 3306
box 0 0 6 6
use CELL  368
transform 1 0 2841 0 1 2076
box 0 0 6 6
use CELL  369
transform 1 0 2596 0 1 3389
box 0 0 6 6
use CELL  370
transform -1 0 2678 0 1 2481
box 0 0 6 6
use CELL  371
transform 1 0 2410 0 1 3389
box 0 0 6 6
use CELL  372
transform -1 0 2703 0 1 2870
box 0 0 6 6
use CELL  373
transform -1 0 2310 0 1 2481
box 0 0 6 6
use CELL  374
transform 1 0 2709 0 1 1513
box 0 0 6 6
use CELL  375
transform 1 0 2500 0 1 1290
box 0 0 6 6
use CELL  376
transform -1 0 2507 0 -1 1157
box 0 0 6 6
use CELL  377
transform 1 0 2340 0 -1 1832
box 0 0 6 6
use CELL  378
transform -1 0 2780 0 -1 1723
box 0 0 6 6
use CELL  379
transform 1 0 2454 0 1 3458
box 0 0 6 6
use CELL  380
transform -1 0 2351 0 1 2600
box 0 0 6 6
use CELL  381
transform 1 0 2784 0 1 2076
box 0 0 6 6
use CELL  382
transform 1 0 2352 0 1 1290
box 0 0 6 6
use CELL  383
transform -1 0 2702 0 -1 1947
box 0 0 6 6
use CELL  384
transform -1 0 2299 0 1 2600
box 0 0 6 6
use CELL  385
transform 1 0 2359 0 1 1290
box 0 0 6 6
use CELL  386
transform -1 0 2725 0 1 2870
box 0 0 6 6
use CELL  387
transform -1 0 2767 0 1 2971
box 0 0 6 6
use CELL  388
transform -1 0 2443 0 -1 2606
box 0 0 6 6
use CELL  389
transform 1 0 2366 0 1 1290
box 0 0 6 6
use CELL  390
transform -1 0 2348 0 1 3100
box 0 0 6 6
use CELL  391
transform 1 0 2588 0 -1 2876
box 0 0 6 6
use CELL  392
transform 1 0 2770 0 1 2870
box 0 0 6 6
use CELL  393
transform -1 0 2587 0 -1 1832
box 0 0 6 6
use CELL  394
transform -1 0 2426 0 1 3306
box 0 0 6 6
use CELL  395
transform 1 0 2494 0 1 1365
box 0 0 6 6
use CELL  396
transform 1 0 2392 0 1 1290
box 0 0 6 6
use CELL  397
transform 1 0 2452 0 1 1290
box 0 0 6 6
use CELL  398
transform -1 0 2431 0 -1 1832
box 0 0 6 6
use CELL  399
transform 1 0 2531 0 1 3306
box 0 0 6 6
use CELL  400
transform 1 0 2395 0 -1 3106
box 0 0 6 6
use CELL  401
transform 1 0 2763 0 1 2870
box 0 0 6 6
use CELL  402
transform 1 0 2651 0 1 2481
box 0 0 6 6
use CELL  403
transform -1 0 2491 0 1 2600
box 0 0 6 6
use CELL  404
transform -1 0 2322 0 1 1941
box 0 0 6 6
use CELL  405
transform 1 0 2595 0 1 1365
box 0 0 6 6
use CELL  406
transform -1 0 2670 0 1 1290
box 0 0 6 6
use CELL  407
transform 1 0 2537 0 1 1290
box 0 0 6 6
use CELL  408
transform 1 0 2394 0 -1 3464
box 0 0 6 6
use CELL  409
transform 1 0 2569 0 1 3306
box 0 0 6 6
use CELL  410
transform -1 0 2342 0 1 2076
box 0 0 6 6
use CELL  411
transform -1 0 2317 0 1 2481
box 0 0 6 6
use CELL  412
transform 1 0 2617 0 1 1432
box 0 0 6 6
use CELL  413
transform 1 0 2672 0 1 2600
box 0 0 6 6
use CELL  414
transform 1 0 2638 0 1 1622
box 0 0 6 6
use CELL  415
transform 1 0 2351 0 1 1941
box 0 0 6 6
use CELL  416
transform 1 0 2787 0 1 1941
box 0 0 6 6
use CELL  417
transform -1 0 2300 0 -1 2348
box 0 0 6 6
use CELL  418
transform 1 0 2826 0 1 2199
box 0 0 6 6
use CELL  419
transform 1 0 2782 0 1 2342
box 0 0 6 6
use CELL  420
transform -1 0 2661 0 1 1513
box 0 0 6 6
use CELL  421
transform -1 0 2449 0 -1 1296
box 0 0 6 6
use CELL  422
transform -1 0 2432 0 -1 3503
box 0 0 6 6
use CELL  423
transform 1 0 2357 0 1 3389
box 0 0 6 6
use CELL  424
transform 1 0 2647 0 1 2199
box 0 0 6 6
use CELL  425
transform -1 0 2386 0 1 1622
box 0 0 6 6
use CELL  426
transform -1 0 2331 0 1 2481
box 0 0 6 6
use CELL  427
transform -1 0 2655 0 1 3100
box 0 0 6 6
use CELL  428
transform 1 0 2357 0 1 1432
box 0 0 6 6
use CELL  429
transform 1 0 2376 0 1 3458
box 0 0 6 6
use CELL  430
transform -1 0 2509 0 1 1622
box 0 0 6 6
use CELL  431
transform -1 0 2334 0 1 3100
box 0 0 6 6
use CELL  432
transform -1 0 2371 0 -1 1130
box 0 0 6 6
use CELL  433
transform 1 0 2615 0 1 2342
box 0 0 6 6
use CELL  434
transform -1 0 2392 0 1 1124
box 0 0 6 6
use CELL  435
transform 1 0 2818 0 1 2481
box 0 0 6 6
use CELL  436
transform -1 0 2752 0 1 1717
box 0 0 6 6
use CELL  437
transform -1 0 2331 0 -1 1723
box 0 0 6 6
use CELL  438
transform 1 0 2401 0 1 1151
box 0 0 6 6
use CELL  439
transform -1 0 2306 0 1 2199
box 0 0 6 6
use CELL  440
transform 1 0 2691 0 1 2342
box 0 0 6 6
use CELL  441
transform 1 0 2374 0 1 2481
box 0 0 6 6
use CELL  442
transform 1 0 2351 0 1 3458
box 0 0 6 6
use CELL  443
transform -1 0 2386 0 -1 1832
box 0 0 6 6
use CELL  444
transform 1 0 2334 0 1 3306
box 0 0 6 6
use CELL  445
transform 1 0 2440 0 1 1432
box 0 0 6 6
use CELL  446
transform 1 0 2458 0 1 1432
box 0 0 6 6
use CELL  447
transform 1 0 2691 0 1 2745
box 0 0 6 6
use CELL  448
transform 1 0 2368 0 -1 2876
box 0 0 6 6
use CELL  449
transform -1 0 2539 0 1 2745
box 0 0 6 6
use CELL  450
transform -1 0 2327 0 -1 1519
box 0 0 6 6
use CELL  451
transform 1 0 2508 0 1 1151
box 0 0 6 6
use CELL  452
transform 1 0 2425 0 1 1513
box 0 0 6 6
use CELL  453
transform -1 0 2293 0 1 2342
box 0 0 6 6
use CELL  454
transform -1 0 2838 0 1 2481
box 0 0 6 6
use CELL  455
transform -1 0 2632 0 1 1826
box 0 0 6 6
use CELL  456
transform -1 0 2363 0 -1 1157
box 0 0 6 6
use CELL  457
transform -1 0 2728 0 1 2199
box 0 0 6 6
use CELL  458
transform 1 0 2404 0 1 1513
box 0 0 6 6
use CELL  459
transform 1 0 2377 0 1 1513
box 0 0 6 6
use CELL  460
transform -1 0 2528 0 -1 1157
box 0 0 6 6
use CELL  461
transform -1 0 2616 0 1 1432
box 0 0 6 6
use CELL  462
transform 1 0 2656 0 1 3100
box 0 0 6 6
use CELL  463
transform 1 0 2745 0 1 2481
box 0 0 6 6
use CELL  464
transform 1 0 2797 0 1 2199
box 0 0 6 6
use CELL  465
transform -1 0 2476 0 1 1432
box 0 0 6 6
use CELL  466
transform -1 0 2307 0 1 2342
box 0 0 6 6
use CELL  467
transform -1 0 2774 0 1 2971
box 0 0 6 6
use CELL  468
transform -1 0 2358 0 1 3189
box 0 0 6 6
use CELL  469
transform -1 0 2527 0 1 1826
box 0 0 6 6
use CELL  470
transform -1 0 2514 0 1 3389
box 0 0 6 6
use CELL  471
transform 1 0 2627 0 1 2481
box 0 0 6 6
use CELL  472
transform 1 0 2293 0 1 2199
box 0 0 6 6
use CELL  473
transform 1 0 2510 0 1 1622
box 0 0 6 6
use CELL  474
transform -1 0 2637 0 -1 3195
box 0 0 6 6
use CELL  475
transform -1 0 2389 0 1 2600
box 0 0 6 6
use CELL  476
transform 1 0 2747 0 1 2745
box 0 0 6 6
use CELL  477
transform 1 0 2519 0 1 3100
box 0 0 6 6
use CELL  478
transform -1 0 2825 0 1 2199
box 0 0 6 6
use CELL  479
transform -1 0 2645 0 -1 2977
box 0 0 6 6
use CELL  480
transform 1 0 2507 0 1 1290
box 0 0 6 6
use CELL  481
transform 1 0 2617 0 1 1513
box 0 0 6 6
use CELL  482
transform -1 0 2772 0 1 2481
box 0 0 6 6
use CELL  483
transform 1 0 2643 0 1 1513
box 0 0 6 6
use CELL  484
transform -1 0 2670 0 1 2745
box 0 0 6 6
use CELL  485
transform -1 0 2387 0 -1 2487
box 0 0 6 6
use CELL  486
transform -1 0 2661 0 -1 2348
box 0 0 6 6
use CELL  487
transform 1 0 2784 0 1 2870
box 0 0 6 6
use CELL  488
transform -1 0 2716 0 -1 1947
box 0 0 6 6
use CELL  489
transform 1 0 2397 0 1 2745
box 0 0 6 6
use CELL  490
transform -1 0 2332 0 1 2600
box 0 0 6 6
use CELL  491
transform -1 0 2372 0 1 1622
box 0 0 6 6
use CELL  492
transform 1 0 2697 0 1 2971
box 0 0 6 6
use CELL  493
transform 1 0 2451 0 1 2745
box 0 0 6 6
use CELL  494
transform -1 0 2326 0 1 2971
box 0 0 6 6
use CELL  495
transform 1 0 2353 0 1 1717
box 0 0 6 6
use CELL  496
transform 1 0 2754 0 -1 2751
box 0 0 6 6
use CELL  497
transform 1 0 2812 0 1 2600
box 0 0 6 6
use CELL  498
transform -1 0 2670 0 1 1432
box 0 0 6 6
use CELL  499
transform -1 0 2751 0 1 2199
box 0 0 6 6
use CELL  500
transform -1 0 2659 0 1 3189
box 0 0 6 6
use CELL  501
transform 1 0 2473 0 1 2600
box 0 0 6 6
use CELL  502
transform 1 0 2608 0 1 1513
box 0 0 6 6
use CELL  503
transform -1 0 2306 0 1 1513
box 0 0 6 6
use CELL  504
transform -1 0 2391 0 1 3541
box 0 0 6 6
use CELL  505
transform 1 0 2370 0 1 1513
box 0 0 6 6
use CELL  506
transform -1 0 2417 0 1 1941
box 0 0 6 6
use CELL  507
transform -1 0 2334 0 1 2342
box 0 0 6 6
use CELL  508
transform 1 0 2579 0 1 3100
box 0 0 6 6
use CELL  509
transform 1 0 2567 0 1 1290
box 0 0 6 6
use CELL  510
transform 1 0 2576 0 1 1290
box 0 0 6 6
use CELL  511
transform 1 0 2573 0 -1 3395
box 0 0 6 6
use CELL  512
transform -1 0 2402 0 1 1941
box 0 0 6 6
use CELL  513
transform -1 0 2369 0 1 2971
box 0 0 6 6
use CELL  514
transform -1 0 2507 0 1 3389
box 0 0 6 6
use CELL  515
transform -1 0 2320 0 1 2342
box 0 0 6 6
use CELL  516
transform 1 0 2583 0 1 1290
box 0 0 6 6
use CELL  517
transform 1 0 2590 0 1 1290
box 0 0 6 6
use CELL  518
transform 1 0 2602 0 1 1290
box 0 0 6 6
use CELL  519
transform 1 0 2343 0 1 1365
box 0 0 6 6
use CELL  520
transform 1 0 2343 0 1 1432
box 0 0 6 6
use CELL  521
transform -1 0 2370 0 -1 1438
box 0 0 6 6
use CELL  522
transform 1 0 2799 0 1 2076
box 0 0 6 6
use CELL  523
transform 1 0 2440 0 1 2199
box 0 0 6 6
use CELL  524
transform 1 0 2404 0 1 1717
box 0 0 6 6
use CELL  525
transform -1 0 2741 0 1 2745
box 0 0 6 6
use CELL  526
transform 1 0 2318 0 1 3306
box 0 0 6 6
use CELL  527
transform 1 0 2347 0 1 1826
box 0 0 6 6
use CELL  528
transform 1 0 2822 0 1 1826
box 0 0 6 6
use CELL  529
transform 1 0 2771 0 1 1826
box 0 0 6 6
use CELL  530
transform 1 0 2605 0 1 1717
box 0 0 6 6
use CELL  531
transform 1 0 2794 0 1 1941
box 0 0 6 6
use CELL  532
transform -1 0 2414 0 1 2971
box 0 0 6 6
use CELL  533
transform -1 0 2447 0 1 2342
box 0 0 6 6
use CELL  534
transform 1 0 2560 0 1 2199
box 0 0 6 6
use CELL  535
transform 1 0 2377 0 -1 1130
box 0 0 6 6
use CELL  536
transform 1 0 2422 0 1 1151
box 0 0 6 6
use CELL  537
transform -1 0 2586 0 1 3389
box 0 0 6 6
use CELL  538
transform 1 0 2482 0 1 3518
box 0 0 6 6
use CELL  539
transform 1 0 2723 0 1 2971
box 0 0 6 6
use CELL  540
transform 1 0 2385 0 1 3458
box 0 0 6 6
use CELL  541
transform -1 0 2373 0 -1 1723
box 0 0 6 6
use CELL  542
transform -1 0 2459 0 1 2481
box 0 0 6 6
use CELL  543
transform 1 0 2812 0 1 2342
box 0 0 6 6
use CELL  544
transform -1 0 2725 0 1 2076
box 0 0 6 6
use CELL  545
transform 1 0 2360 0 1 2199
box 0 0 6 6
use CELL  546
transform 1 0 2412 0 1 3189
box 0 0 6 6
use CELL  547
transform -1 0 2869 0 1 2600
box 0 0 6 6
use CELL  548
transform 1 0 2427 0 1 3189
box 0 0 6 6
use CELL  549
transform -1 0 2609 0 1 3389
box 0 0 6 6
use CELL  550
transform -1 0 2339 0 1 2600
box 0 0 6 6
use CELL  551
transform -1 0 2391 0 1 1290
box 0 0 6 6
use CELL  552
transform -1 0 2692 0 1 3306
box 0 0 6 6
use CELL  553
transform 1 0 2586 0 1 1365
box 0 0 6 6
use CELL  554
transform 1 0 2445 0 1 3189
box 0 0 6 6
use CELL  555
transform 1 0 2534 0 1 3458
box 0 0 6 6
use CELL  556
transform 1 0 2532 0 1 3189
box 0 0 6 6
use CELL  557
transform -1 0 2330 0 -1 3395
box 0 0 6 6
use CELL  558
transform -1 0 2453 0 1 3458
box 0 0 6 6
use CELL  559
transform -1 0 2807 0 -1 1947
box 0 0 6 6
use CELL  560
transform -1 0 2699 0 1 3189
box 0 0 6 6
use CELL  561
transform 1 0 2729 0 1 2600
box 0 0 6 6
use CELL  562
transform 1 0 2820 0 -1 2082
box 0 0 6 6
use CELL  563
transform 1 0 2714 0 -1 1832
box 0 0 6 6
use CELL  564
transform -1 0 2351 0 1 1290
box 0 0 6 6
use CELL  565
transform 1 0 2350 0 1 2481
box 0 0 6 6
use CELL  566
transform 1 0 2433 0 -1 3547
box 0 0 6 6
use CELL  567
transform -1 0 2786 0 1 1941
box 0 0 6 6
use CELL  568
transform -1 0 2349 0 1 2076
box 0 0 6 6
use CELL  569
transform 1 0 2515 0 1 1151
box 0 0 6 6
use CELL  570
transform -1 0 2636 0 1 3389
box 0 0 6 6
use CELL  571
transform -1 0 2398 0 1 1151
box 0 0 6 6
use CELL  572
transform 1 0 2638 0 -1 2751
box 0 0 6 6
use CELL  573
transform -1 0 2384 0 1 2745
box 0 0 6 6
use CELL  574
transform 1 0 2670 0 1 2870
box 0 0 6 6
use CELL  575
transform 1 0 2373 0 1 1290
box 0 0 6 6
use CELL  576
transform -1 0 2674 0 -1 1723
box 0 0 6 6
use CELL  577
transform -1 0 2647 0 1 1365
box 0 0 6 6
use CELL  578
transform -1 0 2839 0 -1 2606
box 0 0 6 6
use CELL  579
transform -1 0 2854 0 -1 2487
box 0 0 6 6
use CELL  580
transform -1 0 2810 0 -1 2487
box 0 0 6 6
use CELL  581
transform -1 0 2292 0 1 1513
box 0 0 6 6
use CELL  582
transform 1 0 2401 0 -1 3395
box 0 0 6 6
use CELL  583
transform -1 0 2390 0 1 3518
box 0 0 6 6
use CELL  584
transform -1 0 2367 0 1 3100
box 0 0 6 6
use CELL  585
transform 1 0 2569 0 1 1235
box 0 0 6 6
use CELL  586
transform 1 0 2735 0 -1 2977
box 0 0 6 6
use CELL  587
transform 1 0 2316 0 -1 3464
box 0 0 6 6
use CELL  588
transform 1 0 2408 0 -1 3547
box 0 0 6 6
use CELL  589
transform -1 0 2316 0 1 1622
box 0 0 6 6
use CELL  590
transform 1 0 2286 0 -1 3395
box 0 0 6 6
use CELL  591
transform 1 0 2298 0 1 3189
box 0 0 6 6
use CELL  592
transform -1 0 2663 0 1 2971
box 0 0 6 6
use CELL  593
transform 1 0 2658 0 1 3306
box 0 0 6 6
use CELL  594
transform 1 0 2555 0 1 1235
box 0 0 6 6
use CELL  595
transform 1 0 2306 0 1 2971
box 0 0 6 6
use CELL  596
transform -1 0 2521 0 1 2076
box 0 0 6 6
use CELL  597
transform -1 0 2371 0 1 1941
box 0 0 6 6
use CELL  598
transform -1 0 2781 0 1 1622
box 0 0 6 6
use CELL  599
transform -1 0 2744 0 1 2076
box 0 0 6 6
use CELL  600
transform -1 0 2330 0 1 1290
box 0 0 6 6
use CELL  601
transform -1 0 2628 0 1 2342
box 0 0 6 6
use CELL  602
transform -1 0 2672 0 1 1622
box 0 0 6 6
use CELL  603
transform 1 0 2597 0 1 1235
box 0 0 6 6
use CELL  604
transform 1 0 2465 0 1 3100
box 0 0 6 6
use CELL  605
transform -1 0 2626 0 -1 1296
box 0 0 6 6
use CELL  606
transform 1 0 2509 0 1 1235
box 0 0 6 6
use CELL  607
transform 1 0 2564 0 -1 1204
box 0 0 6 6
use CELL  608
transform 1 0 2527 0 1 3458
box 0 0 6 6
use CELL  609
transform 1 0 2335 0 1 1513
box 0 0 6 6
use CELL  610
transform 1 0 2638 0 1 1290
box 0 0 6 6
use CELL  611
transform -1 0 2819 0 1 2076
box 0 0 6 6
use CELL  612
transform 1 0 2372 0 1 1235
box 0 0 6 6
use CELL  613
transform -1 0 2520 0 1 3518
box 0 0 6 6
use CELL  614
transform -1 0 2305 0 1 2971
box 0 0 6 6
use CELL  615
transform -1 0 2341 0 1 3100
box 0 0 6 6
use CELL  616
transform 1 0 2733 0 -1 1628
box 0 0 6 6
use CELL  617
transform 1 0 2382 0 1 3497
box 0 0 6 6
use CELL  618
transform -1 0 2610 0 1 1365
box 0 0 6 6
use CELL  619
transform -1 0 2419 0 1 1826
box 0 0 6 6
use CELL  620
transform 1 0 2316 0 -1 1241
box 0 0 6 6
use CELL  621
transform 1 0 2368 0 1 3497
box 0 0 6 6
use CELL  622
transform -1 0 2765 0 1 1826
box 0 0 6 6
use CELL  623
transform -1 0 2764 0 1 1941
box 0 0 6 6
use CELL  624
transform 1 0 2372 0 1 1941
box 0 0 6 6
use CELL  625
transform -1 0 2551 0 -1 1519
box 0 0 6 6
use CELL  626
transform 1 0 2664 0 1 2971
box 0 0 6 6
use CELL  627
transform 1 0 2712 0 1 3189
box 0 0 6 6
use CELL  628
transform -1 0 2419 0 1 3306
box 0 0 6 6
use CELL  629
transform 1 0 2339 0 1 2199
box 0 0 6 6
use CELL  630
transform -1 0 2472 0 -1 1157
box 0 0 6 6
use CELL  631
transform 1 0 2529 0 1 3497
box 0 0 6 6
use CELL  632
transform -1 0 2737 0 1 2076
box 0 0 6 6
use CELL  633
transform -1 0 2362 0 1 2971
box 0 0 6 6
use CELL  634
transform 1 0 2494 0 1 1235
box 0 0 6 6
use CELL  635
transform 1 0 2457 0 1 1235
box 0 0 6 6
use CELL  636
transform -1 0 2407 0 1 2971
box 0 0 6 6
use CELL  637
transform -1 0 2326 0 1 2199
box 0 0 6 6
use CELL  638
transform 1 0 2312 0 -1 1832
box 0 0 6 6
use CELL  639
transform -1 0 2636 0 1 3100
box 0 0 6 6
use CELL  640
transform -1 0 2713 0 1 1826
box 0 0 6 6
use CELL  641
transform 1 0 2494 0 1 1151
box 0 0 6 6
use CELL  642
transform -1 0 2350 0 1 1941
box 0 0 6 6
use CELL  643
transform 1 0 2379 0 1 1235
box 0 0 6 6
use CELL  644
transform -1 0 2700 0 1 3100
box 0 0 6 6
use CELL  645
transform 1 0 2402 0 1 3100
box 0 0 6 6
use CELL  646
transform 1 0 2312 0 -1 2606
box 0 0 6 6
use CELL  647
transform 1 0 2337 0 1 1235
box 0 0 6 6
use CELL  648
transform 1 0 2536 0 1 3497
box 0 0 6 6
use CELL  649
transform 1 0 2585 0 1 1198
box 0 0 6 6
use CELL  650
transform -1 0 2412 0 1 3306
box 0 0 6 6
use CELL  651
transform -1 0 2324 0 1 1717
box 0 0 6 6
use CELL  652
transform -1 0 2681 0 1 1941
box 0 0 6 6
use CELL  653
transform 1 0 2771 0 1 2600
box 0 0 6 6
use CELL  654
transform -1 0 2365 0 -1 1628
box 0 0 6 6
use CELL  655
transform 1 0 2536 0 1 1235
box 0 0 6 6
use CELL  656
transform -1 0 2316 0 1 1290
box 0 0 6 6
use CELL  657
transform 1 0 2543 0 -1 1241
box 0 0 6 6
use CELL  658
transform 1 0 2701 0 -1 3106
box 0 0 6 6
use CELL  659
transform 1 0 2357 0 1 1198
box 0 0 6 6
use CELL  660
transform 1 0 2343 0 1 1198
box 0 0 6 6
use CELL  661
transform 1 0 2318 0 1 2745
box 0 0 6 6
use CELL  662
transform -1 0 2783 0 -1 2082
box 0 0 6 6
use CELL  663
transform -1 0 2341 0 -1 2348
box 0 0 6 6
use CELL  664
transform -1 0 2337 0 1 3389
box 0 0 6 6
use CELL  665
transform 1 0 2395 0 1 2076
box 0 0 6 6
use CELL  666
transform -1 0 2683 0 1 1717
box 0 0 6 6
use CELL  667
transform 1 0 2483 0 1 1198
box 0 0 6 6
use CELL  668
transform -1 0 2677 0 1 2076
box 0 0 6 6
use CELL  669
transform 1 0 2343 0 1 3389
box 0 0 6 6
use CELL  670
transform -1 0 2323 0 1 1622
box 0 0 6 6
use CELL  671
transform -1 0 2847 0 1 2481
box 0 0 6 6
use CELL  672
transform -1 0 2310 0 1 1717
box 0 0 6 6
use CELL  673
transform 1 0 2433 0 1 3497
box 0 0 6 6
use CELL  674
transform -1 0 2337 0 1 3189
box 0 0 6 6
use CELL  675
transform -1 0 2422 0 -1 3464
box 0 0 6 6
use CELL  676
transform 1 0 2674 0 1 3189
box 0 0 6 6
use CELL  677
transform -1 0 2651 0 -1 2751
box 0 0 6 6
use CELL  678
transform -1 0 2467 0 -1 2082
box 0 0 6 6
use CELL  679
transform 1 0 2642 0 1 1432
box 0 0 6 6
use CELL  680
transform 1 0 2429 0 1 3389
box 0 0 6 6
use CELL  681
transform 1 0 2702 0 1 1513
box 0 0 6 6
use CELL  682
transform -1 0 2655 0 -1 2876
box 0 0 6 6
use CELL  683
transform 1 0 2746 0 -1 2348
box 0 0 6 6
use CELL  684
transform 1 0 2338 0 1 1622
box 0 0 6 6
use CELL  685
transform -1 0 2363 0 1 2745
box 0 0 6 6
use CELL  686
transform 1 0 2338 0 1 3189
box 0 0 6 6
use CELL  687
transform 1 0 2695 0 -1 1519
box 0 0 6 6
use CELL  688
transform -1 0 2328 0 1 1365
box 0 0 6 6
use CELL  689
transform -1 0 2560 0 -1 1519
box 0 0 6 6
use CELL  690
transform -1 0 2544 0 1 3306
box 0 0 6 6
use CELL  691
transform 1 0 2337 0 1 1941
box 0 0 6 6
use CELL  692
transform 1 0 2336 0 1 1432
box 0 0 6 6
use CELL  693
transform 1 0 2427 0 1 3518
box 0 0 6 6
use CELL  694
transform -1 0 2335 0 1 1365
box 0 0 6 6
use CELL  695
transform 1 0 2329 0 1 1198
box 0 0 6 6
use CELL  696
transform -1 0 2746 0 -1 1628
box 0 0 6 6
use CELL  697
transform 1 0 2311 0 -1 2751
box 0 0 6 6
use CELL  698
transform 1 0 2371 0 1 1198
box 0 0 6 6
use CELL  699
transform -1 0 2365 0 -1 1371
box 0 0 6 6
use CELL  700
transform 1 0 2390 0 1 1198
box 0 0 6 6
use CELL  701
transform -1 0 2382 0 1 2076
box 0 0 6 6
use CELL  702
transform 1 0 2314 0 -1 1519
box 0 0 6 6
use CELL  703
transform 1 0 2592 0 1 1198
box 0 0 6 6
use CELL  704
transform 1 0 2317 0 -1 1296
box 0 0 6 6
use CELL  705
transform 1 0 2732 0 1 3189
box 0 0 6 6
use CELL  706
transform 1 0 2367 0 1 2199
box 0 0 6 6
use CELL  707
transform -1 0 2533 0 1 1717
box 0 0 6 6
use CELL  708
transform 1 0 2541 0 1 1198
box 0 0 6 6
use CELL  709
transform -1 0 2588 0 -1 1438
box 0 0 6 6
use CELL  710
transform 1 0 2557 0 1 1198
box 0 0 6 6
use CELL  711
transform 1 0 2571 0 1 1198
box 0 0 6 6
use CELL  712
transform 1 0 2351 0 1 1235
box 0 0 6 6
use CELL  713
transform 1 0 2365 0 1 1235
box 0 0 6 6
use CELL  714
transform -1 0 2360 0 1 3100
box 0 0 6 6
use CELL  715
transform -1 0 2506 0 1 1432
box 0 0 6 6
use CELL  716
transform -1 0 2327 0 -1 2348
box 0 0 6 6
use CELL  717
transform 1 0 2487 0 1 1151
box 0 0 6 6
use CELL  718
transform 1 0 2432 0 -1 3106
box 0 0 6 6
use CELL  719
transform -1 0 2360 0 1 1826
box 0 0 6 6
use CELL  720
transform -1 0 2560 0 1 1365
box 0 0 6 6
use CELL  721
transform -1 0 2666 0 -1 3195
box 0 0 6 6
use CELL  722
transform 1 0 2629 0 1 2076
box 0 0 6 6
use CELL  723
transform -1 0 2718 0 1 2870
box 0 0 6 6
use CELL  724
transform 1 0 2403 0 1 1235
box 0 0 6 6
use CELL  725
transform 1 0 2332 0 -1 2487
box 0 0 6 6
use CELL  726
transform 1 0 2645 0 -1 1628
box 0 0 6 6
use CELL  727
transform -1 0 2473 0 -1 1371
box 0 0 6 6
use CELL  728
transform -1 0 2311 0 1 2076
box 0 0 6 6
use CELL  729
transform -1 0 2522 0 1 3306
box 0 0 6 6
use CELL  730
transform 1 0 2444 0 1 1941
box 0 0 6 6
use CELL  731
transform -1 0 2567 0 1 1941
box 0 0 6 6
use CELL  732
transform -1 0 2292 0 1 2481
box 0 0 6 6
use CELL  733
transform 1 0 2517 0 1 1622
box 0 0 6 6
use CELL  734
transform -1 0 2381 0 1 2870
box 0 0 6 6
use CELL  735
transform 1 0 2343 0 1 1151
box 0 0 6 6
use CELL  736
transform 1 0 2840 0 1 2600
box 0 0 6 6
use CELL  737
transform -1 0 2444 0 1 2870
box 0 0 6 6
use CELL  738
transform 1 0 2558 0 1 2481
box 0 0 6 6
use CELL  739
transform -1 0 2576 0 1 3100
box 0 0 6 6
use CELL  740
transform 1 0 2775 0 -1 2348
box 0 0 6 6
use CELL  741
transform 1 0 2456 0 1 2971
box 0 0 6 6
use CELL  742
transform 1 0 2274 0 1 2199
box 0 0 6 6
use CELL  743
transform -1 0 2500 0 -1 2205
box 0 0 6 6
use CELL  744
transform 1 0 2368 0 1 3100
box 0 0 6 6
use CELL  745
transform 1 0 2469 0 -1 1130
box 0 0 6 6
use CELL  746
transform -1 0 2783 0 -1 2876
box 0 0 6 6
use CELL  747
transform 1 0 2337 0 1 3458
box 0 0 6 6
use CELL  748
transform 1 0 2557 0 1 3458
box 0 0 6 6
use CELL  749
transform 1 0 2383 0 -1 3195
box 0 0 6 6
use CELL  750
transform -1 0 2383 0 1 2971
box 0 0 6 6
use CELL  751
transform 1 0 2336 0 1 3497
box 0 0 6 6
use CELL  752
transform 1 0 2343 0 1 3497
box 0 0 6 6
use CELL  753
transform -1 0 2446 0 -1 3503
box 0 0 6 6
use CELL  754
transform 1 0 2618 0 1 1365
box 0 0 6 6
use CELL  755
transform -1 0 2663 0 -1 2751
box 0 0 6 6
use CELL  756
transform -1 0 2624 0 -1 1241
box 0 0 6 6
use CELL  757
transform 1 0 2517 0 1 3389
box 0 0 6 6
use CELL  758
transform 1 0 2396 0 1 3497
box 0 0 6 6
use CELL  759
transform 1 0 2576 0 1 1235
box 0 0 6 6
use CELL  760
transform 1 0 2487 0 1 1235
box 0 0 6 6
use CELL  761
transform -1 0 2304 0 1 1826
box 0 0 6 6
use CELL  762
transform 1 0 2344 0 1 1235
box 0 0 6 6
use CELL  763
transform 1 0 2358 0 1 1235
box 0 0 6 6
use CELL  764
transform -1 0 2732 0 -1 2876
box 0 0 6 6
use CELL  765
transform 1 0 2756 0 1 2870
box 0 0 6 6
use CELL  766
transform -1 0 2779 0 1 1941
box 0 0 6 6
use CELL  767
transform -1 0 2695 0 1 1826
box 0 0 6 6
use CELL  768
transform 1 0 2445 0 1 1235
box 0 0 6 6
use CELL  769
transform 1 0 2346 0 1 1717
box 0 0 6 6
use CELL  770
transform -1 0 2337 0 1 1290
box 0 0 6 6
use CELL  771
transform 1 0 2562 0 1 1235
box 0 0 6 6
use CELL  772
transform 1 0 2550 0 1 3458
box 0 0 6 6
use CELL  773
transform 1 0 2686 0 1 3189
box 0 0 6 6
use CELL  774
transform 1 0 2336 0 1 1365
box 0 0 6 6
use CELL  775
transform 1 0 2362 0 1 2481
box 0 0 6 6
use CELL  776
transform -1 0 2348 0 1 2342
box 0 0 6 6
use CELL  777
transform 1 0 2447 0 1 3497
box 0 0 6 6
use CELL  778
transform 1 0 2304 0 -1 2751
box 0 0 6 6
use CELL  779
transform 1 0 2408 0 1 3497
box 0 0 6 6
use CELL  780
transform -1 0 2801 0 1 1622
box 0 0 6 6
use CELL  781
transform -1 0 2630 0 1 1513
box 0 0 6 6
use CELL  782
transform 1 0 2588 0 1 1235
box 0 0 6 6
use CELL  783
transform -1 0 2313 0 1 1513
box 0 0 6 6
use CELL  784
transform 1 0 2418 0 1 1124
box 0 0 6 6
use CELL  785
transform -1 0 2712 0 -1 3312
box 0 0 6 6
use CELL  786
transform 1 0 2479 0 1 3497
box 0 0 6 6
use CELL  787
transform -1 0 2818 0 1 2199
box 0 0 6 6
use CELL  788
transform 1 0 2559 0 1 3497
box 0 0 6 6
use CELL  789
transform 1 0 2506 0 1 3497
box 0 0 6 6
use CELL  790
transform 1 0 2712 0 -1 3312
box 0 0 6 6
use CELL  791
transform 1 0 2604 0 1 1235
box 0 0 6 6
use CELL  792
transform 1 0 2330 0 1 1235
box 0 0 6 6
use CELL  793
transform 1 0 2513 0 1 3497
box 0 0 6 6
use CELL  794
transform 1 0 2461 0 1 3497
box 0 0 6 6
use CELL  795
transform -1 0 2781 0 1 2745
box 0 0 6 6
use CELL  796
transform -1 0 2814 0 1 1941
box 0 0 6 6
use CELL  797
transform -1 0 2685 0 1 3306
box 0 0 6 6
use CELL  798
transform 1 0 2870 0 -1 2606
box 0 0 6 6
use CELL  799
transform 1 0 2363 0 -1 1519
box 0 0 6 6
use CELL  800
transform 1 0 2494 0 1 3497
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 2603 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 2567 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 2572 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 2572 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 2540 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 2536 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 2524 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 2526 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 2629 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 2504 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 2476 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 2452 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 2432 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 2461 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 2449 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 2437 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 2485 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 2758 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 2806 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 2793 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 2764 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 2795 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 2719 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 2705 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 2798 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 2783 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 2722 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 2708 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 2503 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 2398 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 2476 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 2536 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 2548 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 2552 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 2536 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 2400 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 2396 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 2467 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 2476 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 2479 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 2452 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 2464 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 2473 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 2476 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 2453 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 2449 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 2509 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 2531 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 2567 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 2575 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 2548 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 2577 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 2590 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 2605 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 2627 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 2653 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 2665 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 2637 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 2666 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 2678 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 2351 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 2389 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 2501 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 2332 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 2327 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 2512 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 2494 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 2674 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 2720 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 2716 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 2744 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 2772 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 2725 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 2751 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 2784 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 2345 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 2342 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 2344 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 2545 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 2351 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 2348 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 2350 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 2567 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 2494 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 2473 0 1 3497
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 2467 0 1 3518
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 2430 0 1 3541
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 2614 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 2617 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 2570 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 2497 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 2476 0 1 3497
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 2470 0 1 3518
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 2491 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 2506 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 2491 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 2478 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 2474 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 2497 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 2484 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 2480 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 2469 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 2465 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 2809 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 2796 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 2754 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 2790 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 2729 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-109
transform 1 0 2738 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-110
transform 1 0 2629 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-111
transform 1 0 2622 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-112
transform 1 0 2596 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-113
transform 1 0 2548 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-114
transform 1 0 2545 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-115
transform 1 0 2546 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-116
transform 1 0 2521 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-117
transform 1 0 2509 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-118
transform 1 0 2463 0 1 1151
box 0 0 3 6
use FEEDTHRU  F-119
transform 1 0 2728 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-120
transform 1 0 2716 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-121
transform 1 0 2687 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-122
transform 1 0 2683 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-123
transform 1 0 2636 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-124
transform 1 0 2703 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-125
transform 1 0 2703 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-126
transform 1 0 2630 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-127
transform 1 0 2567 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-128
transform 1 0 2580 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-129
transform 1 0 2525 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-130
transform 1 0 2314 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-131
transform 1 0 2533 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-132
transform 1 0 2537 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-133
transform 1 0 2495 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-134
transform 1 0 2450 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-135
transform 1 0 2455 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-136
transform 1 0 2431 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-137
transform 1 0 2500 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-138
transform 1 0 2482 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-139
transform 1 0 2476 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-140
transform 1 0 2477 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-141
transform 1 0 2512 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-142
transform 1 0 2512 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-143
transform 1 0 2546 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-144
transform 1 0 2555 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-145
transform 1 0 2599 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-146
transform 1 0 2560 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-147
transform 1 0 2552 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-148
transform 1 0 2546 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-149
transform 1 0 2416 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-150
transform 1 0 2411 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-151
transform 1 0 2425 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-152
transform 1 0 2424 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-153
transform 1 0 2420 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-154
transform 1 0 2645 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-155
transform 1 0 2699 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-156
transform 1 0 2438 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-157
transform 1 0 2540 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-158
transform 1 0 2519 0 1 3497
box 0 0 3 6
use FEEDTHRU  F-159
transform 1 0 2649 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-160
transform 1 0 2693 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-161
transform 1 0 2695 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-162
transform 1 0 2765 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-163
transform 1 0 2752 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-164
transform 1 0 2771 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-165
transform 1 0 2784 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-166
transform 1 0 2752 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-167
transform 1 0 2772 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-168
transform 1 0 2803 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-169
transform 1 0 2790 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-170
transform 1 0 2767 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-171
transform 1 0 2392 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-172
transform 1 0 2437 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-173
transform 1 0 2455 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-174
transform 1 0 2464 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-175
transform 1 0 2624 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-176
transform 1 0 2632 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-177
transform 1 0 2656 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-178
transform 1 0 2621 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-179
transform 1 0 2597 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-180
transform 1 0 2587 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-181
transform 1 0 2324 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-182
transform 1 0 2318 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-183
transform 1 0 2311 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-184
transform 1 0 2298 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-185
transform 1 0 2465 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-186
transform 1 0 2465 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-187
transform 1 0 2481 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-188
transform 1 0 2410 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-189
transform 1 0 2696 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-190
transform 1 0 2494 0 1 3518
box 0 0 3 6
use FEEDTHRU  F-191
transform 1 0 2732 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-192
transform 1 0 2732 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-193
transform 1 0 2729 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-194
transform 1 0 2662 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-195
transform 1 0 2680 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-196
transform 1 0 2626 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-197
transform 1 0 2586 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-198
transform 1 0 2521 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-199
transform 1 0 2500 0 1 3497
box 0 0 3 6
use FEEDTHRU  F-200
transform 1 0 2497 0 1 3518
box 0 0 3 6
use FEEDTHRU  F-201
transform 1 0 2453 0 1 3541
box 0 0 3 6
use FEEDTHRU  F-202
transform 1 0 2422 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-203
transform 1 0 2422 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-204
transform 1 0 2419 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-205
transform 1 0 2416 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-206
transform 1 0 2377 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-207
transform 1 0 2356 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-208
transform 1 0 2522 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-209
transform 1 0 2566 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-210
transform 1 0 2358 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-211
transform 1 0 2531 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-212
transform 1 0 2700 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-213
transform 1 0 2765 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-214
transform 1 0 2431 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-215
transform 1 0 2347 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-216
transform 1 0 2403 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-217
transform 1 0 2407 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-218
transform 1 0 2391 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-219
transform 1 0 2408 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-220
transform 1 0 2468 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-221
transform 1 0 2459 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-222
transform 1 0 2566 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-223
transform 1 0 2470 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-224
transform 1 0 2468 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-225
transform 1 0 2447 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-226
transform 1 0 2446 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-227
transform 1 0 2458 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-228
transform 1 0 2438 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-229
transform 1 0 2443 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-230
transform 1 0 2382 0 1 3541
box 0 0 3 6
use FEEDTHRU  F-231
transform 1 0 2390 0 1 3518
box 0 0 3 6
use FEEDTHRU  F-232
transform 1 0 2405 0 1 3497
box 0 0 3 6
use FEEDTHRU  F-233
transform 1 0 2407 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-234
transform 1 0 2648 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-235
transform 1 0 2686 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-236
transform 1 0 2717 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-237
transform 1 0 2473 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-238
transform 1 0 2431 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-239
transform 1 0 2440 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-240
transform 1 0 2658 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-241
transform 1 0 2631 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-242
transform 1 0 2654 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-243
transform 1 0 2692 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-244
transform 1 0 2415 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-245
transform 1 0 2413 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-246
transform 1 0 2405 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-247
transform 1 0 2339 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-248
transform 1 0 2554 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-249
transform 1 0 2593 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-250
transform 1 0 2839 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-251
transform 1 0 2809 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-252
transform 1 0 2838 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-253
transform 1 0 2860 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-254
transform 1 0 2781 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-255
transform 1 0 2790 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-256
transform 1 0 2706 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-257
transform 1 0 2709 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-258
transform 1 0 2700 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-259
transform 1 0 2717 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-260
transform 1 0 2768 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-261
transform 1 0 2338 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-262
transform 1 0 2500 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-263
transform 1 0 2446 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-264
transform 1 0 2428 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-265
transform 1 0 2423 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-266
transform 1 0 2434 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-267
transform 1 0 2439 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-268
transform 1 0 2435 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-269
transform 1 0 2699 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-270
transform 1 0 2667 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-271
transform 1 0 2629 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-272
transform 1 0 2707 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-273
transform 1 0 2777 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-274
transform 1 0 2465 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-275
transform 1 0 2467 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-276
transform 1 0 2466 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-277
transform 1 0 2456 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-278
transform 1 0 2743 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-279
transform 1 0 2781 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-280
transform 1 0 2480 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-281
transform 1 0 2509 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-282
transform 1 0 2500 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-283
transform 1 0 2483 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-284
transform 1 0 2480 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-285
transform 1 0 2480 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-286
transform 1 0 2472 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-287
transform 1 0 2468 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-288
transform 1 0 2453 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-289
transform 1 0 2447 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-290
transform 1 0 2431 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-291
transform 1 0 2433 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-292
transform 1 0 2414 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-293
transform 1 0 2438 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-294
transform 1 0 2383 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-295
transform 1 0 2371 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-296
transform 1 0 2367 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-297
transform 1 0 2376 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-298
transform 1 0 2382 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-299
transform 1 0 2324 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-300
transform 1 0 2753 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-301
transform 1 0 2740 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-302
transform 1 0 2753 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-303
transform 1 0 2766 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-304
transform 1 0 2756 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-305
transform 1 0 2603 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-306
transform 1 0 2386 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-307
transform 1 0 2348 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-308
transform 1 0 2425 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-309
transform 1 0 2402 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-310
transform 1 0 2410 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-311
transform 1 0 2415 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-312
transform 1 0 2411 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-313
transform 1 0 2414 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-314
transform 1 0 2416 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-315
transform 1 0 2427 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-316
transform 1 0 2423 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-317
transform 1 0 2389 0 1 1151
box 0 0 3 6
use FEEDTHRU  F-318
transform 1 0 2420 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-319
transform 1 0 2431 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-320
transform 1 0 2436 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-321
transform 1 0 2432 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-322
transform 1 0 2386 0 1 1151
box 0 0 3 6
use FEEDTHRU  F-323
transform 1 0 2374 0 1 1124
box 0 0 3 6
use FEEDTHRU  F-324
transform 1 0 2719 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-325
transform 1 0 2769 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-326
transform 1 0 2563 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-327
transform 1 0 2575 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-328
transform 1 0 2606 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-329
transform 1 0 2611 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-330
transform 1 0 2605 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-331
transform 1 0 2564 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-332
transform 1 0 2597 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-333
transform 1 0 2635 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-334
transform 1 0 2614 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-335
transform 1 0 2603 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-336
transform 1 0 2612 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-337
transform 1 0 2540 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-338
transform 1 0 2544 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-339
transform 1 0 2513 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-340
transform 1 0 2495 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-341
transform 1 0 2444 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-342
transform 1 0 2762 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-343
transform 1 0 2725 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-344
transform 1 0 2738 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-345
transform 1 0 2683 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-346
transform 1 0 2684 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-347
transform 1 0 2688 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-348
transform 1 0 2755 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-349
transform 1 0 2750 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-350
transform 1 0 2741 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-351
transform 1 0 2806 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-352
transform 1 0 2784 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-353
transform 1 0 2410 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-354
transform 1 0 2410 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-355
transform 1 0 2402 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-356
transform 1 0 2500 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-357
transform 1 0 2506 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-358
transform 1 0 2381 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-359
transform 1 0 2417 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-360
transform 1 0 2425 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-361
transform 1 0 2524 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-362
transform 1 0 2507 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-363
transform 1 0 2492 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-364
transform 1 0 2632 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-365
transform 1 0 2594 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-366
transform 1 0 2635 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-367
transform 1 0 2601 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-368
transform 1 0 2632 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-369
transform 1 0 2670 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-370
transform 1 0 2702 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-371
transform 1 0 2710 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-372
transform 1 0 2780 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-373
transform 1 0 2557 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-374
transform 1 0 2637 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-375
transform 1 0 2639 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-376
transform 1 0 2706 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-377
transform 1 0 2706 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-378
transform 1 0 2679 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-379
transform 1 0 2702 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-380
transform 1 0 2699 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-381
transform 1 0 2679 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-382
transform 1 0 2716 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-383
transform 1 0 2701 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-384
transform 1 0 2398 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-385
transform 1 0 2465 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-386
transform 1 0 2507 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-387
transform 1 0 2523 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-388
transform 1 0 2602 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-389
transform 1 0 2435 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-390
transform 1 0 2387 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-391
transform 1 0 2392 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-392
transform 1 0 2399 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-393
transform 1 0 2608 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-394
transform 1 0 2401 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-395
transform 1 0 2401 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-396
transform 1 0 2455 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-397
transform 1 0 2459 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-398
transform 1 0 2401 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-399
transform 1 0 2485 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-400
transform 1 0 2401 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-401
transform 1 0 2392 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-402
transform 1 0 2392 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-403
transform 1 0 2392 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-404
transform 1 0 2653 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-405
transform 1 0 2635 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-406
transform 1 0 2627 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-407
transform 1 0 2728 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-408
transform 1 0 2759 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-409
transform 1 0 2763 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-410
transform 1 0 2734 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-411
transform 1 0 2757 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-412
transform 1 0 2398 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-413
transform 1 0 2398 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-414
transform 1 0 2398 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-415
transform 1 0 2398 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-416
transform 1 0 2390 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-417
transform 1 0 2561 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-418
transform 1 0 2557 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-419
transform 1 0 2527 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-420
transform 1 0 2486 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-421
transform 1 0 2500 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-422
transform 1 0 2509 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-423
transform 1 0 2549 0 1 3497
box 0 0 3 6
use FEEDTHRU  F-424
transform 1 0 2570 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-425
transform 1 0 2636 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-426
transform 1 0 2383 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-427
transform 1 0 2551 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-428
transform 1 0 2580 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-429
transform 1 0 2402 0 1 3497
box 0 0 3 6
use FEEDTHRU  F-430
transform 1 0 2413 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-431
transform 1 0 2477 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-432
transform 1 0 2492 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-433
transform 1 0 2508 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-434
transform 1 0 2516 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-435
transform 1 0 2567 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-436
transform 1 0 2522 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-437
transform 1 0 2584 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-438
transform 1 0 2611 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-439
transform 1 0 2692 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-440
transform 1 0 2750 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-441
transform 1 0 2770 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-442
transform 1 0 2682 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-443
transform 1 0 2719 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-444
transform 1 0 2704 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-445
transform 1 0 2657 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-446
transform 1 0 2656 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-447
transform 1 0 2707 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-448
transform 1 0 2695 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-449
transform 1 0 2669 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-450
transform 1 0 2668 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-451
transform 1 0 2638 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-452
transform 1 0 2408 0 1 3518
box 0 0 3 6
use FEEDTHRU  F-453
transform 1 0 2414 0 1 3497
box 0 0 3 6
use FEEDTHRU  F-454
transform 1 0 2405 0 1 3518
box 0 0 3 6
use FEEDTHRU  F-455
transform 1 0 2462 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-456
transform 1 0 2447 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-457
transform 1 0 2511 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-458
transform 1 0 2531 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-459
transform 1 0 2582 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-460
transform 1 0 2579 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-461
transform 1 0 2590 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-462
transform 1 0 2548 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-463
transform 1 0 2540 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-464
transform 1 0 2537 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-465
transform 1 0 2521 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-466
transform 1 0 2521 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-467
transform 1 0 2480 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-468
transform 1 0 2485 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-469
transform 1 0 2494 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-470
transform 1 0 2479 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-471
transform 1 0 2464 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-472
transform 1 0 2446 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-473
transform 1 0 2441 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-474
transform 1 0 2464 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-475
transform 1 0 2787 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-476
transform 1 0 2358 0 1 3497
box 0 0 3 6
use FEEDTHRU  F-477
transform 1 0 2373 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-478
transform 1 0 2391 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-479
transform 1 0 2382 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-480
transform 1 0 2657 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-481
transform 1 0 2628 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-482
transform 1 0 2635 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-483
transform 1 0 2641 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-484
transform 1 0 2609 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-485
transform 1 0 2723 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-486
transform 1 0 2554 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-487
transform 1 0 2435 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-488
transform 1 0 2448 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-489
transform 1 0 2515 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-490
transform 1 0 2501 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-491
transform 1 0 2516 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-492
transform 1 0 2405 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-493
transform 1 0 2419 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-494
transform 1 0 2398 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-495
transform 1 0 2468 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-496
transform 1 0 2429 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-497
transform 1 0 2449 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-498
transform 1 0 2445 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-499
transform 1 0 2432 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-500
transform 1 0 2432 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-501
transform 1 0 2380 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-502
transform 1 0 2442 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-503
transform 1 0 2379 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-504
transform 1 0 2388 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-505
transform 1 0 2370 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-506
transform 1 0 2355 0 1 3497
box 0 0 3 6
use FEEDTHRU  F-507
transform 1 0 2548 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-508
transform 1 0 2551 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-509
transform 1 0 2599 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-510
transform 1 0 2625 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-511
transform 1 0 2632 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-512
transform 1 0 2686 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-513
transform 1 0 2732 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-514
transform 1 0 2719 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-515
transform 1 0 2747 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-516
transform 1 0 2751 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-517
transform 1 0 2728 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-518
transform 1 0 2787 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-519
transform 1 0 2413 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-520
transform 1 0 2416 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-521
transform 1 0 2419 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-522
transform 1 0 2419 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-523
transform 1 0 2417 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-524
transform 1 0 2437 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-525
transform 1 0 2518 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-526
transform 1 0 2513 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-527
transform 1 0 2549 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-528
transform 1 0 2569 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-529
transform 1 0 2457 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-530
transform 1 0 2531 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-531
transform 1 0 2534 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-532
transform 1 0 2486 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-533
transform 1 0 2478 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-534
transform 1 0 2462 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-535
transform 1 0 2391 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-536
transform 1 0 2383 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-537
transform 1 0 2515 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-538
transform 1 0 2492 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-539
transform 1 0 2533 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-540
transform 1 0 2554 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-541
transform 1 0 2558 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-542
transform 1 0 2582 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-543
transform 1 0 2617 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-544
transform 1 0 2593 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-545
transform 1 0 2428 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-546
transform 1 0 2583 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-547
transform 1 0 2516 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-548
transform 1 0 2768 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-549
transform 1 0 2698 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-550
transform 1 0 2657 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-551
transform 1 0 2652 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-552
transform 1 0 2695 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-553
transform 1 0 2371 0 1 1124
box 0 0 3 6
use FEEDTHRU  F-554
transform 1 0 2383 0 1 1151
box 0 0 3 6
use FEEDTHRU  F-555
transform 1 0 2429 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-556
transform 1 0 2433 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-557
transform 1 0 2461 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-558
transform 1 0 2545 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-559
transform 1 0 2536 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-560
transform 1 0 2474 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-561
transform 1 0 2483 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-562
transform 1 0 2518 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-563
transform 1 0 2515 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-564
transform 1 0 2537 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-565
transform 1 0 2561 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-566
transform 1 0 2510 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-567
transform 1 0 2552 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-568
transform 1 0 2546 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-569
transform 1 0 2563 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-570
transform 1 0 2643 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-571
transform 1 0 2612 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-572
transform 1 0 2694 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-573
transform 1 0 2688 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-574
transform 1 0 2703 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-575
transform 1 0 2723 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-576
transform 1 0 2720 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-577
transform 1 0 2703 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-578
transform 1 0 2710 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-579
transform 1 0 2698 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-580
transform 1 0 2672 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-581
transform 1 0 2671 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-582
transform 1 0 2641 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-583
transform 1 0 2607 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-584
transform 1 0 2590 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-585
transform 1 0 2562 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-586
transform 1 0 2561 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-587
transform 1 0 2618 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-588
transform 1 0 2612 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-589
transform 1 0 2617 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-590
transform 1 0 2638 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-591
transform 1 0 2615 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-592
transform 1 0 2600 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-593
transform 1 0 2590 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-594
transform 1 0 2584 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-595
transform 1 0 2558 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-596
transform 1 0 2500 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-597
transform 1 0 2491 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-598
transform 1 0 2425 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-599
transform 1 0 2435 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-600
transform 1 0 2486 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-601
transform 1 0 2696 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-602
transform 1 0 2551 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-603
transform 1 0 2417 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-604
transform 1 0 2421 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-605
transform 1 0 2422 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-606
transform 1 0 2408 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-607
transform 1 0 2413 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-608
transform 1 0 2434 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-609
transform 1 0 2452 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-610
transform 1 0 2461 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-611
transform 1 0 2446 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-612
transform 1 0 2450 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-613
transform 1 0 2473 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-614
transform 1 0 2470 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-615
transform 1 0 2471 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-616
transform 1 0 2477 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-617
transform 1 0 2506 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-618
transform 1 0 2497 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-619
transform 1 0 2480 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-620
transform 1 0 2477 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-621
transform 1 0 2423 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-622
transform 1 0 2418 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-623
transform 1 0 2579 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-624
transform 1 0 2614 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-625
transform 1 0 2599 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-626
transform 1 0 2573 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-627
transform 1 0 2576 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-628
transform 1 0 2525 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-629
transform 1 0 2517 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-630
transform 1 0 2495 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-631
transform 1 0 2509 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-632
transform 1 0 2509 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-633
transform 1 0 2474 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-634
transform 1 0 2473 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-635
transform 1 0 2479 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-636
transform 1 0 2470 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-637
transform 1 0 2458 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-638
transform 1 0 2422 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-639
transform 1 0 2575 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-640
transform 1 0 2543 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-641
transform 1 0 2560 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-642
transform 1 0 2542 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-643
transform 1 0 2541 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-644
transform 1 0 2530 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-645
transform 1 0 2494 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-646
transform 1 0 2491 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-647
transform 1 0 2494 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-648
transform 1 0 2481 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-649
transform 1 0 2477 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-650
transform 1 0 2440 0 1 1151
box 0 0 3 6
use FEEDTHRU  F-651
transform 1 0 2458 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-652
transform 1 0 2438 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-653
transform 1 0 2695 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-654
transform 1 0 2488 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-655
transform 1 0 2470 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-656
transform 1 0 2428 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-657
transform 1 0 2530 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-658
transform 1 0 2552 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-659
transform 1 0 2533 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-660
transform 1 0 2542 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-661
transform 1 0 2560 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-662
transform 1 0 2595 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-663
transform 1 0 2599 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-664
transform 1 0 2659 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-665
transform 1 0 2660 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-666
transform 1 0 2647 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-667
transform 1 0 2641 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-668
transform 1 0 2631 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-669
transform 1 0 2702 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-670
transform 1 0 2705 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-671
transform 1 0 2682 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-672
transform 1 0 2636 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-673
transform 1 0 2645 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-674
transform 1 0 2585 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-675
transform 1 0 2640 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-676
transform 1 0 2560 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-677
transform 1 0 2537 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-678
transform 1 0 2632 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-679
transform 1 0 2594 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-680
transform 1 0 2576 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-681
transform 1 0 2566 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-682
transform 1 0 2563 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-683
transform 1 0 2410 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-684
transform 1 0 2447 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-685
transform 1 0 2438 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-686
transform 1 0 2484 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-687
transform 1 0 2492 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-688
transform 1 0 2507 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-689
transform 1 0 2516 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-690
transform 1 0 2539 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-691
transform 1 0 2560 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-692
transform 1 0 2552 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-693
transform 1 0 2522 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-694
transform 1 0 2395 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-695
transform 1 0 2741 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-696
transform 1 0 2500 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-697
transform 1 0 2525 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-698
transform 1 0 2599 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-699
transform 1 0 2383 0 1 1124
box 0 0 3 6
use FEEDTHRU  F-700
transform 1 0 2613 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-701
transform 1 0 2437 0 1 1151
box 0 0 3 6
use FEEDTHRU  F-702
transform 1 0 2750 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-703
transform 1 0 2669 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-704
transform 1 0 2471 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-705
transform 1 0 2505 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-706
transform 1 0 2513 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-707
transform 1 0 2564 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-708
transform 1 0 2561 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-709
transform 1 0 2581 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-710
transform 1 0 2608 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-711
transform 1 0 2585 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-712
transform 1 0 2555 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-713
transform 1 0 2548 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-714
transform 1 0 2548 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-715
transform 1 0 2507 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-716
transform 1 0 2512 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-717
transform 1 0 2506 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-718
transform 1 0 2636 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-719
transform 1 0 2576 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-720
transform 1 0 2583 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-721
transform 1 0 2547 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-722
transform 1 0 2552 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-723
transform 1 0 2573 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-724
transform 1 0 2560 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-725
transform 1 0 2579 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-726
transform 1 0 2593 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-727
transform 1 0 2628 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-728
transform 1 0 2635 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-729
transform 1 0 2650 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-730
transform 1 0 2743 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-731
transform 1 0 2756 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-732
transform 1 0 2683 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-733
transform 1 0 2722 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-734
transform 1 0 2696 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-735
transform 1 0 2720 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-736
transform 1 0 2676 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-737
transform 1 0 2667 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-738
transform 1 0 2670 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-739
transform 1 0 2609 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-740
transform 1 0 2616 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-741
transform 1 0 2611 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-742
transform 1 0 2558 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-743
transform 1 0 2506 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-744
transform 1 0 2485 0 1 3497
box 0 0 3 6
use FEEDTHRU  F-745
transform 1 0 2479 0 1 3518
box 0 0 3 6
use FEEDTHRU  F-746
transform 1 0 2691 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-747
transform 1 0 2627 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-748
transform 1 0 2682 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-749
transform 1 0 2606 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-750
transform 1 0 2615 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-751
transform 1 0 2543 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-752
transform 1 0 2547 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-753
transform 1 0 2510 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-754
transform 1 0 2492 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-755
transform 1 0 2441 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-756
transform 1 0 2423 0 1 3497
box 0 0 3 6
use FEEDTHRU  F-757
transform 1 0 2417 0 1 3518
box 0 0 3 6
use FEEDTHRU  F-758
transform 1 0 2391 0 1 3541
box 0 0 3 6
use FEEDTHRU  F-759
transform 1 0 2566 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-760
transform 1 0 2556 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-761
transform 1 0 2518 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-762
transform 1 0 2497 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-763
transform 1 0 2537 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-764
transform 1 0 2540 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-765
transform 1 0 2441 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-766
transform 1 0 2506 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-767
transform 1 0 2614 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-768
transform 1 0 2585 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-769
transform 1 0 2617 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-770
transform 1 0 2474 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-771
transform 1 0 2489 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-772
transform 1 0 2586 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-773
transform 1 0 2497 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-774
transform 1 0 2488 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-775
transform 1 0 2491 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-776
transform 1 0 2492 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-777
transform 1 0 2459 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-778
transform 1 0 2498 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-779
transform 1 0 2512 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-780
transform 1 0 2488 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-781
transform 1 0 2482 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-782
transform 1 0 2488 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-783
transform 1 0 2488 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-784
transform 1 0 2475 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-785
transform 1 0 2471 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-786
transform 1 0 2434 0 1 1151
box 0 0 3 6
use FEEDTHRU  F-787
transform 1 0 2581 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-788
transform 1 0 2581 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-789
transform 1 0 2555 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-790
transform 1 0 2557 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-791
transform 1 0 2741 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-792
transform 1 0 2452 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-793
transform 1 0 2456 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-794
transform 1 0 2491 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-795
transform 1 0 2482 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-796
transform 1 0 2465 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-797
transform 1 0 2461 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-798
transform 1 0 2638 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-799
transform 1 0 2644 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-800
transform 1 0 2612 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-801
transform 1 0 2602 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-802
transform 1 0 2569 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-803
transform 1 0 2574 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-804
transform 1 0 2527 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-805
transform 1 0 2506 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-806
transform 1 0 2503 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-807
transform 1 0 2528 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-808
transform 1 0 2424 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-809
transform 1 0 2429 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-810
transform 1 0 2489 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-811
transform 1 0 2504 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-812
transform 1 0 2521 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-813
transform 1 0 2530 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-814
transform 1 0 2534 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-815
transform 1 0 2492 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-816
transform 1 0 2503 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-817
transform 1 0 2449 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-818
transform 1 0 2435 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-819
transform 1 0 2455 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-820
transform 1 0 2630 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-821
transform 1 0 2656 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-822
transform 1 0 2398 0 1 1151
box 0 0 3 6
use FEEDTHRU  F-823
transform 1 0 2438 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-824
transform 1 0 2442 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-825
transform 1 0 2449 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-826
transform 1 0 2432 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-827
transform 1 0 2437 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-828
transform 1 0 2449 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-829
transform 1 0 2485 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-830
transform 1 0 2491 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-831
transform 1 0 2491 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-832
transform 1 0 2498 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-833
transform 1 0 2542 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-834
transform 1 0 2533 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-835
transform 1 0 2528 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-836
transform 1 0 2564 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-837
transform 1 0 2572 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-838
transform 1 0 2545 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-839
transform 1 0 2534 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-840
transform 1 0 2525 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-841
transform 1 0 2459 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-842
transform 1 0 2502 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-843
transform 1 0 2486 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-844
transform 1 0 2668 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-845
transform 1 0 2640 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-846
transform 1 0 2639 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-847
transform 1 0 2466 0 1 1124
box 0 0 3 6
use FEEDTHRU  F-848
transform 1 0 2456 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-849
transform 1 0 2489 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-850
transform 1 0 2500 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-851
transform 1 0 2478 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-852
transform 1 0 2462 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-853
transform 1 0 2462 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-854
transform 1 0 2688 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-855
transform 1 0 2621 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-856
transform 1 0 2702 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-857
transform 1 0 2648 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-858
transform 1 0 2450 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-859
transform 1 0 2539 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-860
transform 1 0 2535 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-861
transform 1 0 2494 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-862
transform 1 0 2488 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-863
transform 1 0 2485 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-864
transform 1 0 2584 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-865
transform 1 0 2596 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-866
transform 1 0 2557 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-867
transform 1 0 2549 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-868
transform 1 0 2543 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-869
transform 1 0 2489 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-870
transform 1 0 2481 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-871
transform 1 0 2671 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-872
transform 1 0 2633 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-873
transform 1 0 2543 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-874
transform 1 0 2603 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-875
transform 1 0 2633 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-876
transform 1 0 2681 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-877
transform 1 0 2623 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-878
transform 1 0 2609 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-879
transform 1 0 2609 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-880
transform 1 0 2558 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-881
transform 1 0 2559 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-882
transform 1 0 2528 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-883
transform 1 0 2514 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-884
transform 1 0 2497 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-885
transform 1 0 2563 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-886
transform 1 0 2492 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-887
transform 1 0 2503 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-888
transform 1 0 2536 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-889
transform 1 0 2510 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-890
transform 1 0 2501 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-891
transform 1 0 2498 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-892
transform 1 0 2509 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-893
transform 1 0 2542 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-894
transform 1 0 2516 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-895
transform 1 0 2486 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-896
transform 1 0 2500 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-897
transform 1 0 2503 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-898
transform 1 0 2735 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-899
transform 1 0 2732 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-900
transform 1 0 2665 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-901
transform 1 0 2683 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-902
transform 1 0 2629 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-903
transform 1 0 2651 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-904
transform 1 0 2689 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-905
transform 1 0 2720 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-906
transform 1 0 2650 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-907
transform 1 0 2735 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-908
transform 1 0 2722 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-909
transform 1 0 2707 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-910
transform 1 0 2754 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-911
transform 1 0 2731 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-912
transform 1 0 2711 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-913
transform 1 0 2809 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-914
transform 1 0 2744 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-915
transform 1 0 2753 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-916
transform 1 0 2758 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-917
transform 1 0 2691 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-918
transform 1 0 2619 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-919
transform 1 0 2599 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-920
transform 1 0 2635 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-921
transform 1 0 2531 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-922
transform 1 0 2527 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-923
transform 1 0 2510 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-924
transform 1 0 2515 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-925
transform 1 0 2501 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-926
transform 1 0 2444 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-927
transform 1 0 2433 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-928
transform 1 0 2432 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-929
transform 1 0 2423 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-930
transform 1 0 2498 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-931
transform 1 0 2522 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-932
transform 1 0 2565 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-933
transform 1 0 2564 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-934
transform 1 0 2621 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-935
transform 1 0 2594 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-936
transform 1 0 2605 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-937
transform 1 0 2644 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-938
transform 1 0 2618 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-939
transform 1 0 2498 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-940
transform 1 0 2528 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-941
transform 1 0 2452 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-942
transform 1 0 2447 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-943
transform 1 0 2458 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-944
transform 1 0 2439 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-945
transform 1 0 2723 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-946
transform 1 0 2729 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-947
transform 1 0 2759 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-948
transform 1 0 2697 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-949
transform 1 0 2685 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-950
transform 1 0 2685 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-951
transform 1 0 2624 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-952
transform 1 0 2628 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-953
transform 1 0 2762 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-954
transform 1 0 2732 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-955
transform 1 0 2697 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-956
transform 1 0 2713 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-957
transform 1 0 2713 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-958
transform 1 0 2693 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-959
transform 1 0 2680 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-960
transform 1 0 2659 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-961
transform 1 0 2663 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-962
transform 1 0 2614 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-963
transform 1 0 2607 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-964
transform 1 0 2592 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-965
transform 1 0 2524 0 1 3458
box 0 0 3 6
use FEEDTHRU  F-966
transform 1 0 2503 0 1 3497
box 0 0 3 6
use FEEDTHRU  F-967
transform 1 0 2566 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-968
transform 1 0 2546 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-969
transform 1 0 2731 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-970
transform 1 0 2602 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-971
transform 1 0 2598 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-972
transform 1 0 2563 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-973
transform 1 0 2545 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-974
transform 1 0 2536 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-975
transform 1 0 2555 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-976
transform 1 0 2533 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-977
transform 1 0 2515 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-978
transform 1 0 2661 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-979
transform 1 0 2582 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-980
transform 1 0 2735 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-981
transform 1 0 2471 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-982
transform 1 0 2477 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-983
transform 1 0 2469 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-984
transform 1 0 2465 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-985
transform 1 0 2450 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-986
transform 1 0 2455 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-987
transform 1 0 2458 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-988
transform 1 0 2629 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-989
transform 1 0 2428 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-990
transform 1 0 2591 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-991
transform 1 0 2608 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-992
transform 1 0 2614 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-993
transform 1 0 2549 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-994
transform 1 0 2564 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-995
transform 1 0 2551 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-996
transform 1 0 2560 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-997
transform 1 0 2572 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-998
transform 1 0 2616 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-999
transform 1 0 2617 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-1000
transform 1 0 2638 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-1001
transform 1 0 2755 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-1002
transform 1 0 2774 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1003
transform 1 0 2787 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-1004
transform 1 0 2755 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-1005
transform 1 0 2775 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-1006
transform 1 0 2714 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-1007
transform 1 0 2563 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-1008
transform 1 0 2566 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-1009
transform 1 0 2610 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-1010
transform 1 0 2611 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-1011
transform 1 0 2632 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-1012
transform 1 0 2639 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-1013
transform 1 0 2659 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1014
transform 1 0 2653 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-1015
transform 1 0 2643 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-1016
transform 1 0 2678 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-1017
transform 1 0 2717 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-1018
transform 1 0 2533 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-1019
transform 1 0 2538 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-1020
transform 1 0 2504 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-1021
transform 1 0 2520 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-1022
transform 1 0 2528 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-1023
transform 1 0 2579 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-1024
transform 1 0 2576 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-1025
transform 1 0 2587 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-1026
transform 1 0 2626 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-1027
transform 1 0 2600 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-1028
transform 1 0 2564 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-1029
transform 1 0 2569 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-1030
transform 1 0 2569 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1031
transform 1 0 2537 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-1032
transform 1 0 2533 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-1033
transform 1 0 2521 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-1034
transform 1 0 2523 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-1035
transform 1 0 2482 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-1036
transform 1 0 2476 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-1037
transform 1 0 2473 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-1038
transform 1 0 2512 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-1039
transform 1 0 2524 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-1040
transform 1 0 2549 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-1041
transform 1 0 2506 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-1042
transform 1 0 2509 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-1043
transform 1 0 2521 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-1044
transform 1 0 2568 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-1045
transform 1 0 2572 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-1046
transform 1 0 2593 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-1047
transform 1 0 2690 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-1048
transform 1 0 2513 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-1049
transform 1 0 2501 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-1050
transform 1 0 2493 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-1051
transform 1 0 2558 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-1052
transform 1 0 2507 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-1053
transform 1 0 2499 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-1054
transform 1 0 2483 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-1055
transform 1 0 2524 0 1 1198
box 0 0 3 6
use FEEDTHRU  F-1056
transform 1 0 2527 0 1 1235
box 0 0 3 6
use FEEDTHRU  F-1057
transform 1 0 2543 0 1 1290
box 0 0 3 6
use FEEDTHRU  F-1058
transform 1 0 2530 0 1 1365
box 0 0 3 6
use FEEDTHRU  F-1059
transform 1 0 2533 0 1 1432
box 0 0 3 6
use FEEDTHRU  F-1060
transform 1 0 2542 0 1 1513
box 0 0 3 6
use FEEDTHRU  F-1061
transform 1 0 2513 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-1062
transform 1 0 2509 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-1063
transform 1 0 2435 0 1 3389
box 0 0 3 6
use FEEDTHRU  F-1064
transform 1 0 2459 0 1 3306
box 0 0 3 6
use FEEDTHRU  F-1065
transform 1 0 2475 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-1066
transform 1 0 2483 0 1 3100
box 0 0 3 6
use FEEDTHRU  F-1067
transform 1 0 2531 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-1068
transform 1 0 2528 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-1069
transform 1 0 2549 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-1070
transform 1 0 2545 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-1071
transform 1 0 2533 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-1072
transform 1 0 2556 0 1 3189
box 0 0 3 6
use FEEDTHRU  F-1073
transform 1 0 2549 0 1 2971
box 0 0 3 6
use FEEDTHRU  F-1074
transform 1 0 2546 0 1 2870
box 0 0 3 6
use FEEDTHRU  F-1075
transform 1 0 2551 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-1076
transform 1 0 2590 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-1077
transform 1 0 2570 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-1078
transform 1 0 2534 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-1079
transform 1 0 2539 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-1080
transform 1 0 2539 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1081
transform 1 0 2510 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-1082
transform 1 0 2506 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-1083
transform 1 0 2605 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1084
transform 1 0 2579 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-1085
transform 1 0 2578 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-1086
transform 1 0 2551 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-1087
transform 1 0 2559 0 1 1622
box 0 0 3 6
use FEEDTHRU  F-1088
transform 1 0 2545 0 1 1717
box 0 0 3 6
use FEEDTHRU  F-1089
transform 1 0 2563 0 1 1826
box 0 0 3 6
use FEEDTHRU  F-1090
transform 1 0 2573 0 1 1941
box 0 0 3 6
use FEEDTHRU  F-1091
transform 1 0 2599 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1092
transform 1 0 2593 0 1 2199
box 0 0 3 6
use FEEDTHRU  F-1093
transform 1 0 2594 0 1 2342
box 0 0 3 6
use FEEDTHRU  F-1094
transform 1 0 2624 0 1 2481
box 0 0 3 6
use FEEDTHRU  F-1095
transform 1 0 2650 0 1 2600
box 0 0 3 6
use FEEDTHRU  F-1096
transform 1 0 2611 0 1 2745
box 0 0 3 6
use FEEDTHRU  F-1097
transform 1 0 2600 0 1 2870
box 0 0 3 6
<< metal1 >>
rect 2359 1121 2373 1122
rect 2375 1121 2379 1122
rect 2384 1121 2388 1122
rect 2467 1121 2474 1122
rect 2361 1131 2400 1132
rect 2375 1133 2388 1134
rect 2384 1135 2410 1136
rect 2372 1137 2385 1138
rect 2372 1139 2397 1140
rect 2390 1141 2436 1142
rect 2369 1143 2391 1144
rect 2419 1143 2439 1144
rect 2422 1145 2465 1146
rect 2441 1147 2492 1148
rect 2467 1149 2527 1150
rect 2354 1158 2419 1159
rect 2368 1160 2478 1161
rect 2375 1162 2394 1163
rect 2384 1164 2431 1165
rect 2387 1166 2434 1167
rect 2390 1168 2425 1169
rect 2397 1170 2413 1171
rect 2402 1172 2413 1173
rect 2421 1172 2566 1173
rect 2426 1174 2439 1175
rect 2399 1176 2440 1177
rect 2435 1178 2473 1179
rect 2323 1180 2437 1181
rect 2441 1180 2479 1181
rect 2458 1182 2476 1183
rect 2461 1184 2467 1185
rect 2464 1186 2511 1187
rect 2470 1188 2514 1189
rect 2481 1190 2499 1191
rect 2495 1192 2526 1193
rect 2505 1194 2549 1195
rect 2516 1196 2597 1197
rect 2327 1205 2393 1206
rect 2397 1205 2402 1206
rect 2412 1205 2417 1206
rect 2424 1205 2429 1206
rect 2421 1207 2426 1208
rect 2418 1209 2423 1210
rect 2439 1209 2444 1210
rect 2436 1211 2441 1212
rect 2433 1213 2438 1214
rect 2430 1215 2435 1216
rect 2466 1215 2471 1216
rect 2481 1215 2486 1216
rect 2478 1217 2483 1218
rect 2475 1219 2480 1220
rect 2472 1221 2477 1222
rect 2510 1221 2523 1222
rect 2516 1223 2535 1224
rect 2525 1225 2529 1226
rect 2513 1227 2526 1228
rect 2548 1227 2554 1228
rect 2547 1229 2584 1230
rect 2550 1231 2569 1232
rect 2586 1231 2623 1232
rect 2595 1233 2620 1234
rect 2317 1242 2393 1243
rect 2325 1244 2340 1245
rect 2332 1246 2466 1247
rect 2335 1248 2460 1249
rect 2395 1250 2469 1251
rect 2398 1252 2402 1253
rect 2411 1252 2417 1253
rect 2417 1254 2429 1255
rect 2314 1256 2430 1257
rect 2432 1258 2438 1259
rect 2434 1260 2463 1261
rect 2435 1262 2441 1263
rect 2443 1262 2451 1263
rect 2476 1262 2490 1263
rect 2470 1264 2478 1265
rect 2479 1264 2493 1265
rect 2482 1266 2496 1267
rect 2485 1268 2499 1269
rect 2522 1268 2548 1269
rect 2528 1270 2545 1271
rect 2386 1272 2530 1273
rect 2534 1272 2557 1273
rect 2550 1274 2566 1275
rect 2525 1276 2551 1277
rect 2501 1278 2527 1279
rect 2553 1278 2575 1279
rect 2531 1280 2554 1281
rect 2583 1280 2663 1281
rect 2586 1282 2616 1283
rect 2595 1284 2634 1285
rect 2618 1286 2666 1287
rect 2636 1288 2650 1289
rect 2659 1288 2676 1289
rect 2314 1297 2319 1298
rect 2323 1297 2331 1298
rect 2325 1299 2430 1300
rect 2349 1301 2594 1302
rect 2357 1303 2643 1304
rect 2360 1305 2487 1306
rect 2403 1307 2412 1308
rect 2409 1309 2424 1310
rect 2412 1311 2427 1312
rect 2415 1313 2418 1314
rect 2421 1313 2433 1314
rect 2424 1315 2436 1316
rect 2433 1317 2451 1318
rect 2367 1319 2452 1320
rect 2442 1321 2466 1322
rect 2444 1323 2463 1324
rect 2448 1325 2460 1326
rect 2464 1325 2493 1326
rect 2468 1327 2478 1328
rect 2471 1329 2527 1330
rect 2480 1331 2499 1332
rect 2492 1333 2496 1334
rect 2501 1333 2517 1334
rect 2504 1335 2530 1336
rect 2507 1337 2551 1338
rect 2531 1339 2545 1340
rect 2534 1341 2554 1342
rect 2537 1343 2557 1344
rect 2549 1345 2560 1346
rect 2474 1347 2559 1348
rect 2552 1349 2566 1350
rect 2561 1351 2575 1352
rect 2602 1351 2637 1352
rect 2605 1353 2622 1354
rect 2615 1355 2666 1356
rect 2584 1357 2616 1358
rect 2618 1357 2643 1358
rect 2633 1359 2650 1360
rect 2632 1361 2660 1362
rect 2645 1363 2663 1364
rect 2323 1372 2382 1373
rect 2351 1374 2394 1375
rect 2357 1376 2379 1377
rect 2372 1378 2422 1379
rect 2375 1380 2416 1381
rect 2403 1382 2427 1383
rect 2409 1384 2415 1385
rect 2399 1386 2409 1387
rect 2412 1386 2418 1387
rect 2424 1386 2430 1387
rect 2433 1386 2439 1387
rect 2448 1386 2454 1387
rect 2442 1388 2448 1389
rect 2451 1388 2457 1389
rect 2471 1388 2499 1389
rect 2477 1390 2481 1391
rect 2474 1392 2478 1393
rect 2483 1392 2490 1393
rect 2486 1394 2490 1395
rect 2492 1394 2496 1395
rect 2464 1396 2493 1397
rect 2507 1396 2511 1397
rect 2504 1398 2508 1399
rect 2504 1400 2517 1401
rect 2513 1402 2588 1403
rect 2534 1404 2544 1405
rect 2531 1406 2535 1407
rect 2564 1406 2609 1407
rect 2581 1408 2631 1409
rect 2561 1410 2581 1411
rect 2552 1412 2562 1413
rect 2549 1414 2553 1415
rect 2546 1416 2550 1417
rect 2537 1418 2547 1419
rect 2584 1418 2616 1419
rect 2501 1420 2584 1421
rect 2593 1420 2609 1421
rect 2632 1420 2656 1421
rect 2602 1422 2634 1423
rect 2602 1424 2666 1425
rect 2635 1426 2650 1427
rect 2638 1428 2676 1429
rect 2652 1430 2669 1431
rect 2290 1439 2385 1440
rect 2304 1441 2309 1442
rect 2329 1441 2403 1442
rect 2343 1443 2487 1444
rect 2350 1445 2412 1446
rect 2357 1447 2418 1448
rect 2365 1449 2454 1450
rect 2372 1451 2427 1452
rect 2378 1453 2418 1454
rect 2381 1455 2400 1456
rect 2323 1457 2400 1458
rect 2414 1457 2436 1458
rect 2333 1459 2415 1460
rect 2432 1459 2457 1460
rect 2438 1461 2451 1462
rect 2393 1463 2439 1464
rect 2447 1463 2466 1464
rect 2429 1465 2448 1466
rect 2453 1465 2481 1466
rect 2471 1467 2556 1468
rect 2495 1469 2532 1470
rect 2489 1471 2496 1472
rect 2483 1473 2490 1474
rect 2477 1475 2484 1476
rect 2498 1475 2520 1476
rect 2507 1477 2529 1478
rect 2492 1479 2508 1480
rect 2510 1479 2523 1480
rect 2504 1481 2511 1482
rect 2549 1481 2598 1482
rect 2552 1483 2601 1484
rect 2516 1485 2553 1486
rect 2561 1485 2574 1486
rect 2543 1487 2562 1488
rect 2534 1489 2544 1490
rect 2534 1491 2550 1492
rect 2564 1491 2568 1492
rect 2546 1493 2565 1494
rect 2580 1493 2595 1494
rect 2583 1495 2591 1496
rect 2591 1497 2612 1498
rect 2608 1499 2616 1500
rect 2630 1499 2669 1500
rect 2633 1501 2672 1502
rect 2649 1503 2688 1504
rect 2650 1505 2685 1506
rect 2652 1507 2691 1508
rect 2653 1509 2660 1510
rect 2655 1511 2694 1512
rect 2287 1520 2302 1521
rect 2297 1522 2385 1523
rect 2308 1524 2424 1525
rect 2311 1526 2316 1527
rect 2353 1526 2412 1527
rect 2370 1528 2499 1529
rect 2374 1530 2448 1531
rect 2393 1532 2403 1533
rect 2332 1534 2403 1535
rect 2411 1534 2472 1535
rect 2417 1536 2421 1537
rect 2414 1538 2418 1539
rect 2432 1538 2502 1539
rect 2438 1540 2457 1541
rect 2438 1542 2487 1543
rect 2450 1544 2487 1545
rect 2322 1546 2451 1547
rect 2321 1548 2472 1549
rect 2459 1550 2478 1551
rect 2465 1552 2481 1553
rect 2453 1554 2466 1555
rect 2435 1556 2454 1557
rect 2483 1556 2525 1557
rect 2489 1558 2505 1559
rect 2367 1560 2490 1561
rect 2367 1562 2493 1563
rect 2495 1562 2537 1563
rect 2510 1564 2514 1565
rect 2507 1566 2515 1567
rect 2507 1568 2707 1569
rect 2519 1570 2558 1571
rect 2522 1572 2570 1573
rect 2528 1574 2576 1575
rect 2360 1576 2528 1577
rect 2534 1576 2540 1577
rect 2543 1576 2697 1577
rect 2531 1578 2543 1579
rect 2552 1578 2582 1579
rect 2567 1580 2612 1581
rect 2573 1582 2618 1583
rect 2578 1584 2586 1585
rect 2591 1584 2609 1585
rect 2594 1586 2630 1587
rect 2597 1588 2624 1589
rect 2561 1590 2597 1591
rect 2560 1592 2626 1593
rect 2600 1594 2627 1595
rect 2564 1596 2600 1597
rect 2615 1596 2665 1597
rect 2653 1598 2659 1599
rect 2656 1600 2710 1601
rect 2668 1602 2701 1603
rect 2671 1604 2704 1605
rect 2670 1606 2698 1607
rect 2685 1608 2780 1609
rect 2687 1610 2719 1611
rect 2690 1612 2722 1613
rect 2693 1614 2745 1615
rect 2650 1616 2695 1617
rect 2649 1618 2668 1619
rect 2724 1618 2793 1619
rect 2765 1620 2773 1621
rect 2311 1629 2451 1630
rect 2312 1631 2424 1632
rect 2325 1633 2511 1634
rect 2326 1635 2647 1636
rect 2340 1637 2412 1638
rect 2353 1639 2368 1640
rect 2368 1641 2499 1642
rect 2375 1643 2490 1644
rect 2414 1645 2517 1646
rect 2420 1647 2424 1648
rect 2417 1649 2421 1650
rect 2417 1651 2493 1652
rect 2438 1653 2451 1654
rect 2453 1653 2463 1654
rect 2459 1655 2582 1656
rect 2319 1657 2460 1658
rect 2465 1657 2475 1658
rect 2456 1659 2466 1660
rect 2314 1661 2457 1662
rect 2480 1661 2496 1662
rect 2471 1663 2481 1664
rect 2483 1663 2502 1664
rect 2384 1665 2502 1666
rect 2486 1667 2493 1668
rect 2507 1667 2779 1668
rect 2518 1669 2547 1670
rect 2522 1671 2525 1672
rect 2525 1673 2528 1674
rect 2531 1673 2535 1674
rect 2539 1673 2682 1674
rect 2536 1675 2541 1676
rect 2477 1677 2538 1678
rect 2552 1677 2561 1678
rect 2557 1679 2568 1680
rect 2569 1679 2574 1680
rect 2570 1681 2576 1682
rect 2578 1681 2592 1682
rect 2564 1683 2580 1684
rect 2599 1683 2604 1684
rect 2596 1685 2601 1686
rect 2608 1685 2643 1686
rect 2626 1687 2634 1688
rect 2629 1689 2637 1690
rect 2623 1691 2631 1692
rect 2639 1691 2772 1692
rect 2651 1693 2722 1694
rect 2660 1695 2665 1696
rect 2675 1695 2731 1696
rect 2697 1697 2741 1698
rect 2694 1699 2697 1700
rect 2693 1701 2756 1702
rect 2700 1703 2752 1704
rect 2658 1705 2700 1706
rect 2703 1705 2712 1706
rect 2706 1707 2721 1708
rect 2718 1709 2735 1710
rect 2724 1711 2787 1712
rect 2709 1713 2724 1714
rect 2708 1715 2749 1716
rect 2792 1715 2800 1716
rect 2312 1724 2460 1725
rect 2323 1726 2331 1727
rect 2326 1728 2454 1729
rect 2341 1730 2445 1731
rect 2369 1732 2475 1733
rect 2375 1734 2427 1735
rect 2417 1736 2502 1737
rect 2447 1738 2463 1739
rect 2450 1740 2463 1741
rect 2417 1742 2451 1743
rect 2456 1742 2460 1743
rect 2402 1744 2457 1745
rect 2465 1744 2469 1745
rect 2471 1744 2517 1745
rect 2474 1746 2481 1747
rect 2477 1748 2484 1749
rect 2486 1748 2496 1749
rect 2501 1748 2511 1749
rect 2355 1750 2511 1751
rect 2507 1752 2514 1753
rect 2299 1754 2508 1755
rect 2537 1754 2550 1755
rect 2525 1756 2538 1757
rect 2543 1756 2562 1757
rect 2552 1758 2580 1759
rect 2558 1760 2761 1761
rect 2564 1762 2577 1763
rect 2546 1764 2565 1765
rect 2534 1766 2547 1767
rect 2522 1768 2535 1769
rect 2522 1770 2541 1771
rect 2567 1770 2583 1771
rect 2573 1772 2595 1773
rect 2591 1774 2607 1775
rect 2603 1776 2716 1777
rect 2570 1778 2604 1779
rect 2630 1778 2655 1779
rect 2630 1780 2658 1781
rect 2633 1782 2688 1783
rect 2612 1784 2634 1785
rect 2639 1784 2670 1785
rect 2618 1786 2640 1787
rect 2651 1786 2737 1787
rect 2636 1788 2652 1789
rect 2672 1788 2682 1789
rect 2642 1790 2673 1791
rect 2660 1792 2682 1793
rect 2600 1794 2661 1795
rect 2600 1796 2646 1797
rect 2675 1796 2706 1797
rect 2684 1798 2740 1799
rect 2627 1800 2685 1801
rect 2693 1800 2752 1801
rect 2696 1802 2767 1803
rect 2696 1804 2820 1805
rect 2699 1806 2770 1807
rect 2708 1808 2779 1809
rect 2528 1810 2709 1811
rect 2711 1810 2782 1811
rect 2720 1812 2797 1813
rect 2702 1814 2722 1815
rect 2723 1814 2785 1815
rect 2729 1816 2800 1817
rect 2733 1818 2772 1819
rect 2724 1820 2773 1821
rect 2742 1822 2748 1823
rect 2754 1822 2813 1823
rect 2757 1824 2810 1825
rect 2302 1833 2307 1834
rect 2316 1833 2460 1834
rect 2320 1835 2443 1836
rect 2330 1837 2407 1838
rect 2337 1839 2424 1840
rect 2358 1841 2688 1842
rect 2362 1843 2782 1844
rect 2381 1845 2394 1846
rect 2391 1847 2400 1848
rect 2403 1847 2412 1848
rect 2412 1849 2529 1850
rect 2415 1851 2533 1852
rect 2418 1853 2421 1854
rect 2433 1853 2463 1854
rect 2439 1855 2445 1856
rect 2456 1855 2461 1856
rect 2453 1857 2458 1858
rect 2450 1859 2455 1860
rect 2447 1861 2452 1862
rect 2469 1861 2524 1862
rect 2481 1863 2487 1864
rect 2487 1865 2502 1866
rect 2492 1867 2500 1868
rect 2493 1869 2517 1870
rect 2471 1871 2518 1872
rect 2537 1871 2542 1872
rect 2534 1873 2539 1874
rect 2544 1873 2562 1874
rect 2549 1875 2554 1876
rect 2546 1877 2551 1878
rect 2556 1877 2559 1878
rect 2313 1879 2560 1880
rect 2564 1879 2575 1880
rect 2600 1879 2694 1880
rect 2603 1881 2614 1882
rect 2604 1883 2677 1884
rect 2610 1885 2691 1886
rect 2594 1887 2692 1888
rect 2627 1889 2632 1890
rect 2606 1891 2629 1892
rect 2576 1893 2608 1894
rect 2651 1893 2745 1894
rect 2681 1895 2695 1896
rect 2684 1897 2689 1898
rect 2696 1897 2782 1898
rect 2711 1899 2743 1900
rect 2714 1901 2764 1902
rect 2717 1903 2722 1904
rect 2720 1905 2734 1906
rect 2724 1907 2760 1908
rect 2723 1909 2737 1910
rect 2726 1911 2740 1912
rect 2729 1913 2834 1914
rect 2741 1915 2755 1916
rect 2751 1917 2772 1918
rect 2753 1919 2767 1920
rect 2757 1921 2763 1922
rect 2639 1923 2757 1924
rect 2633 1925 2641 1926
rect 2765 1925 2797 1926
rect 2769 1927 2817 1928
rect 2768 1929 2820 1930
rect 2778 1931 2848 1932
rect 2777 1933 2813 1934
rect 2732 1935 2813 1936
rect 2784 1937 2803 1938
rect 2799 1939 2806 1940
rect 2302 1948 2427 1949
rect 2309 1950 2430 1951
rect 2317 1952 2390 1953
rect 2320 1954 2446 1955
rect 2324 1956 2401 1957
rect 2323 1958 2496 1959
rect 2345 1960 2515 1961
rect 2348 1962 2692 1963
rect 2359 1964 2547 1965
rect 2366 1966 2392 1967
rect 2397 1966 2533 1967
rect 2403 1968 2502 1969
rect 2402 1970 2461 1971
rect 2406 1972 2421 1973
rect 2439 1972 2460 1973
rect 2418 1974 2439 1975
rect 2465 1974 2551 1975
rect 2469 1976 2623 1977
rect 2478 1978 2514 1979
rect 2454 1980 2478 1981
rect 2433 1982 2454 1983
rect 2380 1984 2433 1985
rect 2487 1984 2529 1985
rect 2493 1986 2535 1987
rect 2457 1988 2493 1989
rect 2508 1988 2550 1989
rect 2442 1990 2508 1991
rect 2351 1992 2442 1993
rect 2517 1992 2566 1993
rect 2504 1994 2517 1995
rect 2523 1994 2568 1995
rect 2481 1996 2523 1997
rect 2538 1996 2571 1997
rect 2537 1998 2554 1999
rect 2544 2000 2577 2001
rect 2499 2002 2544 2003
rect 2337 2004 2499 2005
rect 2556 2004 2583 2005
rect 2559 2006 2586 2007
rect 2564 2008 2698 2009
rect 2574 2010 2601 2011
rect 2541 2012 2574 2013
rect 2511 2014 2541 2015
rect 2475 2016 2511 2017
rect 2451 2018 2475 2019
rect 2604 2018 2626 2019
rect 2610 2020 2643 2021
rect 2613 2022 2646 2023
rect 2607 2024 2613 2025
rect 2580 2026 2607 2027
rect 2615 2026 2779 2027
rect 2628 2028 2655 2029
rect 2648 2030 2662 2031
rect 2640 2032 2661 2033
rect 2658 2034 2706 2035
rect 2631 2036 2658 2037
rect 2670 2036 2697 2037
rect 2673 2038 2700 2039
rect 2672 2040 2798 2041
rect 2694 2042 2715 2043
rect 2702 2044 2852 2045
rect 2708 2046 2724 2047
rect 2720 2048 2749 2049
rect 2676 2050 2721 2051
rect 2726 2050 2764 2051
rect 2729 2052 2761 2053
rect 2732 2054 2806 2055
rect 2636 2056 2733 2057
rect 2751 2056 2846 2057
rect 2765 2058 2795 2059
rect 2768 2060 2792 2061
rect 2771 2062 2775 2063
rect 2753 2064 2773 2065
rect 2741 2066 2755 2067
rect 2756 2066 2776 2067
rect 2744 2068 2758 2069
rect 2717 2070 2746 2071
rect 2688 2072 2718 2073
rect 2812 2072 2817 2073
rect 2817 2074 2825 2075
rect 2294 2083 2457 2084
rect 2301 2085 2427 2086
rect 2306 2087 2463 2088
rect 2315 2089 2430 2090
rect 2308 2091 2430 2092
rect 2324 2093 2517 2094
rect 2344 2095 2442 2096
rect 2351 2097 2433 2098
rect 2299 2099 2433 2100
rect 2347 2101 2351 2102
rect 2357 2101 2478 2102
rect 2375 2103 2496 2104
rect 2377 2105 2508 2106
rect 2392 2107 2568 2108
rect 2336 2109 2394 2110
rect 2396 2109 2538 2110
rect 2399 2111 2421 2112
rect 2402 2113 2487 2114
rect 2414 2115 2553 2116
rect 2438 2117 2520 2118
rect 2447 2119 2460 2120
rect 2287 2121 2460 2122
rect 2453 2123 2478 2124
rect 2471 2125 2475 2126
rect 2354 2127 2475 2128
rect 2483 2127 2493 2128
rect 2489 2129 2499 2130
rect 2501 2129 2508 2130
rect 2501 2131 2505 2132
rect 2275 2133 2505 2134
rect 2528 2133 2559 2134
rect 2534 2135 2556 2136
rect 2534 2137 2544 2138
rect 2537 2139 2547 2140
rect 2564 2139 2568 2140
rect 2576 2139 2628 2140
rect 2585 2141 2592 2142
rect 2588 2143 2880 2144
rect 2594 2145 2601 2146
rect 2606 2145 2631 2146
rect 2606 2147 2613 2148
rect 2609 2149 2616 2150
rect 2630 2149 2740 2150
rect 2639 2151 2646 2152
rect 2654 2151 2667 2152
rect 2654 2153 2661 2154
rect 2657 2155 2733 2156
rect 2669 2157 2724 2158
rect 2672 2159 2771 2160
rect 2672 2161 2818 2162
rect 2684 2163 2758 2164
rect 2699 2165 2712 2166
rect 2705 2167 2721 2168
rect 2717 2169 2730 2170
rect 2702 2171 2718 2172
rect 2735 2171 2783 2172
rect 2751 2173 2825 2174
rect 2748 2175 2753 2176
rect 2754 2175 2768 2176
rect 2708 2177 2756 2178
rect 2696 2179 2709 2180
rect 2696 2181 2808 2182
rect 2763 2183 2838 2184
rect 2760 2185 2765 2186
rect 2772 2185 2786 2186
rect 2745 2187 2774 2188
rect 2636 2189 2747 2190
rect 2636 2191 2643 2192
rect 2642 2193 2649 2194
rect 2775 2193 2789 2194
rect 2791 2193 2805 2194
rect 2794 2195 2808 2196
rect 2797 2197 2811 2198
rect 2816 2197 2821 2198
rect 2840 2197 2877 2198
rect 2288 2206 2457 2207
rect 2291 2208 2437 2209
rect 2301 2210 2430 2211
rect 2304 2212 2463 2213
rect 2305 2214 2458 2215
rect 2309 2216 2433 2217
rect 2318 2218 2500 2219
rect 2333 2220 2487 2221
rect 2343 2222 2490 2223
rect 2357 2224 2533 2225
rect 2369 2226 2511 2227
rect 2372 2228 2553 2229
rect 2378 2230 2475 2231
rect 2382 2232 2508 2233
rect 2388 2234 2394 2235
rect 2399 2234 2470 2235
rect 2329 2236 2401 2237
rect 2439 2236 2460 2237
rect 2322 2238 2461 2239
rect 2445 2240 2545 2241
rect 2466 2242 2484 2243
rect 2475 2244 2538 2245
rect 2487 2246 2502 2247
rect 2493 2248 2505 2249
rect 2477 2250 2506 2251
rect 2495 2252 2503 2253
rect 2350 2254 2497 2255
rect 2511 2254 2517 2255
rect 2513 2256 2548 2257
rect 2514 2258 2520 2259
rect 2522 2258 2539 2259
rect 2523 2260 2780 2261
rect 2529 2262 2535 2263
rect 2535 2264 2541 2265
rect 2558 2264 2563 2265
rect 2555 2266 2560 2267
rect 2549 2268 2557 2269
rect 2565 2268 2571 2269
rect 2567 2270 2578 2271
rect 2568 2272 2574 2273
rect 2582 2272 2620 2273
rect 2588 2274 2599 2275
rect 2591 2276 2602 2277
rect 2592 2278 2610 2279
rect 2604 2280 2657 2281
rect 2623 2282 2733 2283
rect 2626 2284 2631 2285
rect 2629 2286 2637 2287
rect 2632 2288 2643 2289
rect 2639 2290 2693 2291
rect 2638 2292 2667 2293
rect 2641 2294 2670 2295
rect 2644 2296 2655 2297
rect 2672 2296 2824 2297
rect 2680 2298 2718 2299
rect 2606 2300 2718 2301
rect 2684 2302 2724 2303
rect 2683 2304 2721 2305
rect 2696 2306 2814 2307
rect 2698 2308 2715 2309
rect 2701 2310 2792 2311
rect 2704 2312 2712 2313
rect 2708 2314 2739 2315
rect 2707 2316 2730 2317
rect 2720 2318 2771 2319
rect 2726 2320 2774 2321
rect 2729 2322 2753 2323
rect 2732 2324 2756 2325
rect 2735 2326 2765 2327
rect 2744 2328 2783 2329
rect 2753 2330 2786 2331
rect 2756 2332 2789 2333
rect 2759 2334 2808 2335
rect 2762 2336 2811 2337
rect 2767 2338 2791 2339
rect 2797 2338 2805 2339
rect 2807 2338 2854 2339
rect 2810 2340 2841 2341
rect 2859 2340 2864 2341
rect 2866 2340 2871 2341
rect 2281 2349 2340 2350
rect 2288 2351 2440 2352
rect 2291 2353 2306 2354
rect 2290 2355 2437 2356
rect 2295 2357 2303 2358
rect 2312 2357 2349 2358
rect 2332 2359 2512 2360
rect 2345 2361 2407 2362
rect 2353 2363 2482 2364
rect 2382 2365 2419 2366
rect 2385 2367 2545 2368
rect 2388 2369 2437 2370
rect 2430 2371 2470 2372
rect 2445 2373 2467 2374
rect 2397 2375 2467 2376
rect 2448 2377 2470 2378
rect 2350 2379 2449 2380
rect 2457 2379 2491 2380
rect 2472 2381 2479 2382
rect 2472 2383 2506 2384
rect 2475 2385 2485 2386
rect 2502 2385 2512 2386
rect 2343 2387 2503 2388
rect 2342 2389 2401 2390
rect 2514 2389 2551 2390
rect 2517 2391 2581 2392
rect 2487 2393 2518 2394
rect 2523 2393 2554 2394
rect 2523 2395 2563 2396
rect 2538 2397 2542 2398
rect 2496 2399 2539 2400
rect 2556 2399 2587 2400
rect 2547 2401 2557 2402
rect 2336 2403 2548 2404
rect 2336 2405 2786 2406
rect 2559 2407 2584 2408
rect 2592 2407 2627 2408
rect 2595 2409 2626 2410
rect 2577 2411 2596 2412
rect 2598 2411 2623 2412
rect 2571 2413 2599 2414
rect 2535 2415 2572 2416
rect 2493 2417 2536 2418
rect 2460 2419 2494 2420
rect 2601 2419 2617 2420
rect 2565 2421 2602 2422
rect 2529 2423 2566 2424
rect 2499 2425 2530 2426
rect 2329 2427 2500 2428
rect 2604 2427 2635 2428
rect 2568 2429 2605 2430
rect 2532 2431 2569 2432
rect 2319 2433 2533 2434
rect 2619 2433 2748 2434
rect 2629 2435 2659 2436
rect 2638 2437 2668 2438
rect 2670 2439 2768 2440
rect 2676 2441 2740 2442
rect 2683 2443 2718 2444
rect 2701 2445 2719 2446
rect 2680 2447 2701 2448
rect 2644 2449 2680 2450
rect 2712 2449 2733 2450
rect 2698 2451 2734 2452
rect 2697 2453 2724 2454
rect 2720 2455 2770 2456
rect 2704 2457 2722 2458
rect 2632 2459 2704 2460
rect 2729 2459 2789 2460
rect 2730 2461 2817 2462
rect 2744 2463 2813 2464
rect 2753 2465 2774 2466
rect 2726 2467 2753 2468
rect 2756 2467 2777 2468
rect 2755 2469 2763 2470
rect 2759 2471 2792 2472
rect 2735 2473 2759 2474
rect 2736 2475 2850 2476
rect 2770 2477 2780 2478
rect 2807 2477 2837 2478
rect 2810 2479 2840 2480
rect 2287 2488 2340 2489
rect 2287 2490 2295 2491
rect 2297 2490 2302 2491
rect 2305 2490 2505 2491
rect 2322 2492 2360 2493
rect 2326 2494 2494 2495
rect 2312 2496 2493 2497
rect 2327 2498 2533 2499
rect 2330 2500 2349 2501
rect 2334 2502 2530 2503
rect 2345 2504 2437 2505
rect 2353 2506 2366 2507
rect 2406 2506 2415 2507
rect 2418 2506 2427 2507
rect 2430 2506 2451 2507
rect 2432 2508 2449 2509
rect 2475 2508 2605 2509
rect 2478 2510 2508 2511
rect 2484 2512 2520 2513
rect 2499 2514 2514 2515
rect 2517 2514 2544 2515
rect 2502 2516 2517 2517
rect 2490 2518 2502 2519
rect 2531 2518 2536 2519
rect 2534 2520 2539 2521
rect 2511 2522 2538 2523
rect 2481 2524 2511 2525
rect 2553 2524 2562 2525
rect 2565 2524 2574 2525
rect 2568 2526 2577 2527
rect 2547 2528 2568 2529
rect 2320 2530 2547 2531
rect 2571 2530 2592 2531
rect 2550 2532 2571 2533
rect 2541 2534 2550 2535
rect 2586 2534 2610 2535
rect 2454 2536 2586 2537
rect 2598 2536 2637 2537
rect 2384 2538 2598 2539
rect 2601 2538 2628 2539
rect 2556 2540 2601 2541
rect 2486 2542 2556 2543
rect 2612 2542 2632 2543
rect 2472 2544 2631 2545
rect 2469 2546 2472 2547
rect 2466 2548 2469 2549
rect 2619 2548 2646 2549
rect 2583 2550 2619 2551
rect 2625 2550 2652 2551
rect 2634 2552 2683 2553
rect 2595 2554 2634 2555
rect 2342 2556 2595 2557
rect 2658 2556 2707 2557
rect 2622 2558 2658 2559
rect 2670 2558 2674 2559
rect 2654 2560 2670 2561
rect 2676 2560 2774 2561
rect 2703 2562 2707 2563
rect 2700 2564 2704 2565
rect 2712 2564 2811 2565
rect 2715 2566 2777 2567
rect 2718 2568 2770 2569
rect 2679 2570 2719 2571
rect 2667 2572 2680 2573
rect 2721 2572 2725 2573
rect 2697 2574 2722 2575
rect 2697 2576 2843 2577
rect 2730 2578 2761 2579
rect 2733 2580 2764 2581
rect 2640 2582 2734 2583
rect 2616 2584 2640 2585
rect 2580 2586 2616 2587
rect 2736 2586 2846 2587
rect 2755 2588 2792 2589
rect 2758 2590 2837 2591
rect 2766 2592 2820 2593
rect 2788 2594 2809 2595
rect 2785 2596 2808 2597
rect 2752 2598 2786 2599
rect 2788 2598 2805 2599
rect 2839 2598 2862 2599
rect 2287 2607 2326 2608
rect 2301 2609 2505 2610
rect 2313 2611 2360 2612
rect 2320 2613 2347 2614
rect 2327 2615 2514 2616
rect 2328 2617 2786 2618
rect 2334 2619 2483 2620
rect 2337 2621 2568 2622
rect 2349 2623 2354 2624
rect 2352 2625 2547 2626
rect 2358 2627 2514 2628
rect 2361 2629 2493 2630
rect 2365 2631 2535 2632
rect 2375 2633 2380 2634
rect 2387 2633 2586 2634
rect 2414 2635 2417 2636
rect 2432 2635 2435 2636
rect 2438 2635 2680 2636
rect 2446 2637 2451 2638
rect 2449 2639 2517 2640
rect 2452 2641 2565 2642
rect 2458 2643 2571 2644
rect 2471 2645 2568 2646
rect 2479 2647 2502 2648
rect 2486 2649 2604 2650
rect 2488 2651 2556 2652
rect 2498 2653 2508 2654
rect 2501 2655 2511 2656
rect 2504 2657 2538 2658
rect 2510 2659 2544 2660
rect 2516 2661 2520 2662
rect 2522 2661 2532 2662
rect 2525 2663 2634 2664
rect 2426 2665 2526 2666
rect 2537 2665 2631 2666
rect 2540 2667 2562 2668
rect 2546 2669 2574 2670
rect 2552 2671 2592 2672
rect 2549 2673 2592 2674
rect 2549 2675 2577 2676
rect 2555 2677 2595 2678
rect 2558 2679 2598 2680
rect 2561 2681 2601 2682
rect 2582 2683 2610 2684
rect 2585 2685 2613 2686
rect 2588 2687 2628 2688
rect 2594 2689 2619 2690
rect 2600 2691 2616 2692
rect 2606 2693 2646 2694
rect 2612 2695 2652 2696
rect 2615 2697 2637 2698
rect 2618 2699 2640 2700
rect 2624 2701 2683 2702
rect 2633 2703 2658 2704
rect 2636 2705 2655 2706
rect 2665 2705 2789 2706
rect 2677 2707 2722 2708
rect 2680 2709 2704 2710
rect 2683 2711 2707 2712
rect 2694 2713 2859 2714
rect 2697 2715 2798 2716
rect 2698 2717 2761 2718
rect 2701 2719 2767 2720
rect 2704 2721 2725 2722
rect 2707 2723 2725 2724
rect 2715 2725 2875 2726
rect 2718 2727 2780 2728
rect 2730 2729 2792 2730
rect 2733 2731 2770 2732
rect 2733 2733 2828 2734
rect 2736 2735 2838 2736
rect 2742 2737 2808 2738
rect 2745 2739 2811 2740
rect 2763 2741 2868 2742
rect 2782 2743 2862 2744
rect 2296 2752 2341 2753
rect 2303 2754 2309 2755
rect 2312 2754 2320 2755
rect 2306 2756 2314 2757
rect 2319 2756 2326 2757
rect 2322 2758 2329 2759
rect 2328 2760 2514 2761
rect 2343 2762 2347 2763
rect 2349 2762 2353 2763
rect 2369 2762 2550 2763
rect 2375 2764 2556 2765
rect 2386 2766 2417 2767
rect 2415 2768 2435 2769
rect 2433 2770 2447 2771
rect 2436 2772 2450 2773
rect 2442 2774 2530 2775
rect 2458 2776 2533 2777
rect 2457 2778 2468 2779
rect 2460 2780 2568 2781
rect 2463 2782 2480 2783
rect 2466 2784 2483 2785
rect 2481 2786 2499 2787
rect 2484 2788 2502 2789
rect 2362 2790 2503 2791
rect 2493 2792 2505 2793
rect 2495 2794 2604 2795
rect 2499 2796 2511 2797
rect 2505 2798 2523 2799
rect 2508 2800 2526 2801
rect 2516 2802 2539 2803
rect 2517 2804 2541 2805
rect 2382 2806 2542 2807
rect 2523 2808 2586 2809
rect 2550 2810 2559 2811
rect 2564 2810 2651 2811
rect 2473 2812 2566 2813
rect 2574 2812 2601 2813
rect 2577 2814 2589 2815
rect 2534 2816 2590 2817
rect 2535 2818 2547 2819
rect 2547 2820 2553 2821
rect 2553 2822 2562 2823
rect 2562 2824 2583 2825
rect 2580 2826 2592 2827
rect 2594 2826 2643 2827
rect 2595 2828 2607 2829
rect 2592 2830 2608 2831
rect 2601 2832 2613 2833
rect 2604 2834 2616 2835
rect 2610 2836 2625 2837
rect 2613 2838 2619 2839
rect 2625 2838 2634 2839
rect 2628 2840 2637 2841
rect 2637 2842 2684 2843
rect 2643 2844 2647 2845
rect 2668 2844 2728 2845
rect 2668 2846 2678 2847
rect 2686 2846 2699 2847
rect 2689 2848 2705 2849
rect 2661 2850 2705 2851
rect 2701 2852 2718 2853
rect 2701 2854 2737 2855
rect 2707 2856 2711 2857
rect 2680 2858 2708 2859
rect 2713 2858 2721 2859
rect 2730 2858 2740 2859
rect 2736 2860 2759 2861
rect 2742 2862 2752 2863
rect 2727 2864 2743 2865
rect 2745 2864 2755 2865
rect 2723 2866 2746 2867
rect 2782 2866 2792 2867
rect 2683 2868 2782 2869
rect 2300 2877 2341 2878
rect 2296 2879 2301 2880
rect 2309 2879 2400 2880
rect 2313 2881 2388 2882
rect 2319 2883 2384 2884
rect 2296 2885 2385 2886
rect 2321 2887 2500 2888
rect 2324 2889 2494 2890
rect 2328 2891 2334 2892
rect 2343 2891 2346 2892
rect 2349 2891 2352 2892
rect 2358 2891 2437 2892
rect 2357 2893 2515 2894
rect 2376 2895 2602 2896
rect 2390 2897 2503 2898
rect 2367 2899 2503 2900
rect 2405 2901 2560 2902
rect 2439 2903 2566 2904
rect 2415 2905 2440 2906
rect 2457 2905 2476 2906
rect 2460 2907 2470 2908
rect 2478 2907 2482 2908
rect 2481 2909 2485 2910
rect 2490 2909 2506 2910
rect 2493 2911 2509 2912
rect 2508 2913 2518 2914
rect 2355 2915 2518 2916
rect 2523 2915 2569 2916
rect 2526 2917 2536 2918
rect 2532 2919 2536 2920
rect 2529 2921 2533 2922
rect 2544 2921 2551 2922
rect 2547 2923 2551 2924
rect 2547 2925 2554 2926
rect 2562 2925 2566 2926
rect 2538 2927 2563 2928
rect 2538 2929 2542 2930
rect 2580 2929 2584 2930
rect 2577 2931 2581 2932
rect 2574 2933 2578 2934
rect 2592 2933 2792 2934
rect 2595 2935 2623 2936
rect 2607 2937 2617 2938
rect 2613 2939 2620 2940
rect 2604 2941 2614 2942
rect 2631 2941 2647 2942
rect 2634 2943 2714 2944
rect 2637 2945 2647 2946
rect 2637 2947 2699 2948
rect 2668 2949 2672 2950
rect 2683 2949 2763 2950
rect 2689 2951 2696 2952
rect 2689 2953 2770 2954
rect 2692 2955 2766 2956
rect 2710 2957 2721 2958
rect 2658 2959 2711 2960
rect 2730 2959 2734 2960
rect 2733 2961 2737 2962
rect 2628 2963 2737 2964
rect 2625 2965 2629 2966
rect 2739 2965 2761 2966
rect 2742 2967 2749 2968
rect 2751 2967 2757 2968
rect 2754 2969 2760 2970
rect 2296 2978 2301 2979
rect 2299 2980 2467 2981
rect 2307 2982 2385 2983
rect 2314 2984 2346 2985
rect 2320 2986 2334 2987
rect 2329 2988 2518 2989
rect 2349 2990 2388 2991
rect 2351 2992 2410 2993
rect 2352 2994 2391 2995
rect 2355 2996 2551 2997
rect 2357 2998 2372 2999
rect 2358 3000 2452 3001
rect 2360 3002 2400 3003
rect 2381 3004 2515 3005
rect 2381 3006 2434 3007
rect 2384 3008 2440 3009
rect 2396 3010 2539 3011
rect 2409 3012 2470 3013
rect 2412 3014 2548 3015
rect 2424 3016 2479 3017
rect 2365 3018 2479 3019
rect 2430 3020 2491 3021
rect 2433 3022 2473 3023
rect 2445 3024 2503 3025
rect 2402 3026 2503 3027
rect 2403 3028 2494 3029
rect 2460 3030 2527 3031
rect 2484 3032 2533 3033
rect 2487 3034 2536 3035
rect 2490 3036 2545 3037
rect 2493 3038 2509 3039
rect 2508 3040 2560 3041
rect 2511 3042 2563 3043
rect 2514 3044 2566 3045
rect 2517 3046 2569 3047
rect 2526 3048 2578 3049
rect 2529 3050 2581 3051
rect 2532 3052 2584 3053
rect 2541 3054 2614 3055
rect 2544 3056 2617 3057
rect 2559 3058 2611 3059
rect 2562 3060 2620 3061
rect 2565 3062 2623 3063
rect 2568 3064 2632 3065
rect 2577 3066 2638 3067
rect 2586 3068 2647 3069
rect 2610 3070 2672 3071
rect 2613 3072 2696 3073
rect 2622 3074 2690 3075
rect 2625 3076 2687 3077
rect 2628 3078 2693 3079
rect 2631 3080 2651 3081
rect 2634 3082 2644 3083
rect 2463 3084 2635 3085
rect 2637 3084 2705 3085
rect 2640 3086 2708 3087
rect 2661 3088 2666 3089
rect 2663 3090 2731 3091
rect 2666 3092 2734 3093
rect 2689 3094 2757 3095
rect 2692 3096 2760 3097
rect 2698 3098 2773 3099
rect 2299 3107 2313 3108
rect 2306 3109 2316 3110
rect 2317 3109 2353 3110
rect 2329 3111 2350 3112
rect 2332 3113 2441 3114
rect 2336 3115 2397 3116
rect 2343 3117 2512 3118
rect 2356 3119 2452 3120
rect 2362 3121 2473 3122
rect 2372 3123 2385 3124
rect 2381 3125 2444 3126
rect 2406 3127 2410 3128
rect 2419 3127 2425 3128
rect 2425 3129 2431 3130
rect 2434 3129 2446 3130
rect 2470 3129 2479 3130
rect 2473 3131 2482 3132
rect 2476 3133 2485 3134
rect 2479 3135 2488 3136
rect 2482 3137 2491 3138
rect 2485 3139 2494 3140
rect 2494 3141 2503 3142
rect 2460 3143 2504 3144
rect 2500 3145 2509 3146
rect 2506 3147 2515 3148
rect 2509 3149 2518 3150
rect 2512 3151 2533 3152
rect 2518 3153 2527 3154
rect 2521 3155 2530 3156
rect 2544 3155 2549 3156
rect 2541 3157 2546 3158
rect 2557 3157 2575 3158
rect 2568 3159 2582 3160
rect 2562 3161 2570 3162
rect 2523 3163 2564 3164
rect 2466 3165 2525 3166
rect 2577 3165 2585 3166
rect 2610 3165 2618 3166
rect 2613 3167 2645 3168
rect 2614 3169 2706 3170
rect 2620 3171 2693 3172
rect 2622 3173 2704 3174
rect 2637 3175 2647 3176
rect 2638 3177 2641 3178
rect 2586 3179 2642 3180
rect 2587 3181 2633 3182
rect 2663 3181 2682 3182
rect 2666 3183 2685 3184
rect 2689 3183 2731 3184
rect 2628 3185 2691 3186
rect 2625 3187 2630 3188
rect 2700 3187 2728 3188
rect 2299 3196 2307 3197
rect 2302 3198 2313 3199
rect 2312 3200 2326 3201
rect 2306 3202 2326 3203
rect 2315 3204 2319 3205
rect 2315 3206 2397 3207
rect 2322 3208 2441 3209
rect 2332 3210 2483 3211
rect 2335 3212 2426 3213
rect 2339 3214 2495 3215
rect 2356 3216 2388 3217
rect 2359 3218 2384 3219
rect 2368 3220 2373 3221
rect 2380 3220 2444 3221
rect 2404 3222 2410 3223
rect 2417 3222 2491 3223
rect 2419 3224 2737 3225
rect 2439 3226 2486 3227
rect 2448 3228 2513 3229
rect 2460 3230 2477 3231
rect 2463 3232 2480 3233
rect 2466 3234 2471 3235
rect 2469 3236 2474 3237
rect 2472 3238 2507 3239
rect 2484 3240 2501 3241
rect 2487 3242 2504 3243
rect 2493 3244 2510 3245
rect 2496 3246 2519 3247
rect 2505 3248 2522 3249
rect 2424 3250 2521 3251
rect 2508 3252 2525 3253
rect 2511 3254 2549 3255
rect 2514 3256 2546 3257
rect 2523 3258 2567 3259
rect 2526 3260 2582 3261
rect 2529 3262 2561 3263
rect 2539 3264 2558 3265
rect 2542 3266 2655 3267
rect 2558 3268 2639 3269
rect 2561 3270 2642 3271
rect 2563 3272 2573 3273
rect 2564 3274 2645 3275
rect 2569 3276 2609 3277
rect 2573 3278 2588 3279
rect 2584 3280 2665 3281
rect 2600 3282 2621 3283
rect 2609 3284 2679 3285
rect 2612 3286 2618 3287
rect 2614 3288 2672 3289
rect 2615 3290 2636 3291
rect 2618 3292 2625 3293
rect 2627 3292 2682 3293
rect 2629 3294 2698 3295
rect 2630 3296 2685 3297
rect 2646 3298 2691 3299
rect 2649 3300 2704 3301
rect 2676 3302 2701 3303
rect 2700 3304 2708 3305
rect 2309 3313 2316 3314
rect 2319 3313 2497 3314
rect 2321 3315 2326 3316
rect 2335 3315 2485 3316
rect 2368 3317 2378 3318
rect 2380 3317 2390 3318
rect 2383 3319 2393 3320
rect 2398 3319 2411 3320
rect 2402 3321 2650 3322
rect 2407 3323 2425 3324
rect 2404 3325 2409 3326
rect 2414 3325 2473 3326
rect 2417 3327 2506 3328
rect 2424 3329 2434 3330
rect 2436 3329 2461 3330
rect 2451 3331 2467 3332
rect 2454 3333 2470 3334
rect 2463 3335 2717 3336
rect 2448 3337 2464 3338
rect 2439 3339 2449 3340
rect 2290 3341 2440 3342
rect 2466 3341 2509 3342
rect 2475 3343 2491 3344
rect 2478 3345 2494 3346
rect 2487 3347 2635 3348
rect 2493 3349 2512 3350
rect 2487 3351 2513 3352
rect 2496 3353 2515 3354
rect 2499 3355 2524 3356
rect 2515 3357 2530 3358
rect 2517 3359 2540 3360
rect 2518 3361 2527 3362
rect 2538 3361 2562 3362
rect 2544 3363 2559 3364
rect 2547 3365 2565 3366
rect 2559 3367 2613 3368
rect 2568 3369 2625 3370
rect 2571 3371 2619 3372
rect 2573 3373 2592 3374
rect 2553 3375 2575 3376
rect 2584 3375 2601 3376
rect 2587 3377 2628 3378
rect 2609 3379 2653 3380
rect 2615 3381 2622 3382
rect 2630 3381 2663 3382
rect 2637 3383 2684 3384
rect 2646 3385 2674 3386
rect 2655 3387 2688 3388
rect 2696 3387 2701 3388
rect 2311 3396 2319 3397
rect 2320 3396 2333 3397
rect 2328 3398 2425 3399
rect 2331 3400 2346 3401
rect 2335 3402 2437 3403
rect 2334 3404 2440 3405
rect 2371 3406 2390 3407
rect 2374 3408 2393 3409
rect 2377 3410 2384 3411
rect 2392 3410 2409 3411
rect 2398 3412 2476 3413
rect 2402 3414 2464 3415
rect 2408 3416 2513 3417
rect 2411 3418 2449 3419
rect 2414 3420 2479 3421
rect 2418 3422 2467 3423
rect 2420 3424 2452 3425
rect 2430 3426 2455 3427
rect 2436 3428 2488 3429
rect 2442 3430 2494 3431
rect 2445 3432 2497 3433
rect 2495 3434 2569 3435
rect 2499 3436 2503 3437
rect 2498 3438 2572 3439
rect 2501 3440 2548 3441
rect 2504 3442 2554 3443
rect 2507 3444 2560 3445
rect 2515 3446 2529 3447
rect 2522 3448 2588 3449
rect 2525 3450 2605 3451
rect 2538 3452 2635 3453
rect 2541 3454 2619 3455
rect 2571 3456 2638 3457
rect 2287 3465 2463 3466
rect 2324 3467 2446 3468
rect 2356 3469 2372 3470
rect 2359 3471 2375 3472
rect 2379 3471 2412 3472
rect 2383 3473 2391 3474
rect 2392 3473 2536 3474
rect 2403 3475 2415 3476
rect 2406 3477 2409 3478
rect 2415 3477 2449 3478
rect 2421 3479 2437 3480
rect 2424 3481 2443 3482
rect 2474 3481 2496 3482
rect 2477 3483 2499 3484
rect 2486 3485 2508 3486
rect 2501 3487 2523 3488
rect 2504 3489 2517 3490
rect 2504 3491 2526 3492
rect 2520 3493 2542 3494
rect 2523 3495 2545 3496
rect 2550 3495 2572 3496
rect 2577 3495 2585 3496
rect 2323 3504 2360 3505
rect 2356 3506 2389 3507
rect 2391 3506 2407 3507
rect 2393 3508 2404 3509
rect 2406 3508 2428 3509
rect 2409 3510 2416 3511
rect 2418 3510 2425 3511
rect 2441 3510 2521 3511
rect 2468 3512 2475 3513
rect 2471 3514 2478 3515
rect 2480 3514 2487 3515
rect 2495 3514 2524 3515
rect 2498 3516 2502 3517
rect 2504 3516 2519 3517
rect 2550 3516 2557 3517
rect 2563 3516 2571 3517
rect 2383 3525 2392 3526
rect 2388 3527 2481 3528
rect 2392 3529 2419 3530
rect 2394 3531 2407 3532
rect 2397 3533 2410 3534
rect 2431 3533 2469 3534
rect 2437 3535 2472 3536
rect 2454 3537 2499 3538
rect 2495 3539 2519 3540
rect 2377 3548 2384 3549
rect 2389 3548 2393 3549
rect 2395 3548 2455 3549
rect 2409 3550 2432 3551
rect 2441 3550 2449 3551
<< metal2 >>
rect 2359 1121 2360 1125
rect 2372 1121 2373 1125
rect 2375 1121 2376 1125
rect 2378 1121 2379 1125
rect 2384 1121 2385 1125
rect 2387 1121 2388 1125
rect 2467 1121 2468 1125
rect 2473 1121 2474 1125
rect 2361 1131 2362 1152
rect 2399 1131 2400 1152
rect 2375 1129 2376 1134
rect 2387 1133 2388 1152
rect 2384 1129 2385 1136
rect 2409 1135 2410 1152
rect 2372 1129 2373 1138
rect 2384 1137 2385 1152
rect 2372 1139 2373 1152
rect 2396 1139 2397 1152
rect 2390 1129 2391 1142
rect 2435 1141 2436 1152
rect 2369 1129 2370 1144
rect 2390 1143 2391 1152
rect 2419 1143 2420 1152
rect 2438 1143 2439 1152
rect 2422 1129 2423 1146
rect 2464 1145 2465 1152
rect 2441 1147 2442 1152
rect 2491 1147 2492 1152
rect 2467 1129 2468 1150
rect 2526 1149 2527 1152
rect 2354 1156 2355 1159
rect 2418 1158 2419 1199
rect 2368 1156 2369 1161
rect 2477 1156 2478 1161
rect 2375 1156 2376 1163
rect 2393 1156 2394 1163
rect 2384 1156 2385 1165
rect 2430 1164 2431 1199
rect 2387 1156 2388 1167
rect 2433 1166 2434 1199
rect 2390 1156 2391 1169
rect 2424 1168 2425 1199
rect 2397 1170 2398 1199
rect 2412 1156 2413 1171
rect 2402 1156 2403 1173
rect 2412 1172 2413 1199
rect 2421 1172 2422 1199
rect 2565 1172 2566 1199
rect 2426 1156 2427 1175
rect 2438 1156 2439 1175
rect 2399 1156 2400 1177
rect 2439 1176 2440 1199
rect 2435 1156 2436 1179
rect 2472 1178 2473 1199
rect 2323 1180 2324 1199
rect 2436 1180 2437 1199
rect 2441 1156 2442 1181
rect 2478 1180 2479 1199
rect 2458 1156 2459 1183
rect 2475 1182 2476 1199
rect 2461 1156 2462 1185
rect 2466 1184 2467 1199
rect 2464 1156 2465 1187
rect 2510 1186 2511 1199
rect 2470 1156 2471 1189
rect 2513 1188 2514 1199
rect 2481 1190 2482 1199
rect 2498 1190 2499 1199
rect 2495 1156 2496 1193
rect 2525 1192 2526 1199
rect 2505 1156 2506 1195
rect 2548 1194 2549 1199
rect 2516 1196 2517 1199
rect 2596 1196 2597 1199
rect 2327 1205 2328 1236
rect 2392 1205 2393 1236
rect 2397 1203 2398 1206
rect 2401 1205 2402 1236
rect 2412 1203 2413 1206
rect 2416 1205 2417 1236
rect 2424 1203 2425 1206
rect 2428 1205 2429 1236
rect 2421 1203 2422 1208
rect 2425 1207 2426 1236
rect 2418 1203 2419 1210
rect 2422 1209 2423 1236
rect 2439 1203 2440 1210
rect 2443 1209 2444 1236
rect 2436 1203 2437 1212
rect 2440 1211 2441 1236
rect 2433 1203 2434 1214
rect 2437 1213 2438 1236
rect 2430 1203 2431 1216
rect 2434 1215 2435 1236
rect 2466 1203 2467 1216
rect 2470 1215 2471 1236
rect 2481 1203 2482 1216
rect 2485 1215 2486 1236
rect 2478 1203 2479 1218
rect 2482 1217 2483 1236
rect 2475 1203 2476 1220
rect 2479 1219 2480 1236
rect 2472 1203 2473 1222
rect 2476 1221 2477 1236
rect 2501 1221 2502 1236
rect 2501 1203 2502 1222
rect 2510 1203 2511 1222
rect 2522 1221 2523 1236
rect 2516 1203 2517 1224
rect 2534 1223 2535 1236
rect 2525 1203 2526 1226
rect 2528 1225 2529 1236
rect 2513 1203 2514 1228
rect 2525 1227 2526 1236
rect 2531 1227 2532 1236
rect 2531 1203 2532 1228
rect 2548 1203 2549 1228
rect 2553 1227 2554 1236
rect 2547 1229 2548 1236
rect 2583 1229 2584 1236
rect 2550 1231 2551 1236
rect 2568 1203 2569 1232
rect 2586 1231 2587 1236
rect 2622 1231 2623 1236
rect 2595 1233 2596 1236
rect 2619 1233 2620 1236
rect 2317 1240 2318 1243
rect 2392 1240 2393 1243
rect 2325 1244 2326 1291
rect 2339 1244 2340 1291
rect 2332 1246 2333 1291
rect 2465 1246 2466 1291
rect 2335 1248 2336 1291
rect 2459 1248 2460 1291
rect 2395 1240 2396 1251
rect 2468 1250 2469 1291
rect 2398 1240 2399 1253
rect 2401 1240 2402 1253
rect 2411 1252 2412 1291
rect 2416 1240 2417 1253
rect 2417 1254 2418 1291
rect 2428 1240 2429 1255
rect 2314 1256 2315 1291
rect 2429 1256 2430 1291
rect 2422 1240 2423 1259
rect 2423 1258 2424 1291
rect 2425 1240 2426 1259
rect 2426 1258 2427 1291
rect 2432 1258 2433 1291
rect 2437 1240 2438 1259
rect 2434 1240 2435 1261
rect 2462 1260 2463 1291
rect 2435 1262 2436 1291
rect 2440 1240 2441 1263
rect 2443 1240 2444 1263
rect 2450 1262 2451 1291
rect 2476 1240 2477 1263
rect 2489 1262 2490 1291
rect 2470 1240 2471 1265
rect 2477 1264 2478 1291
rect 2479 1240 2480 1265
rect 2492 1264 2493 1291
rect 2482 1240 2483 1267
rect 2495 1266 2496 1291
rect 2485 1240 2486 1269
rect 2498 1268 2499 1291
rect 2522 1240 2523 1269
rect 2547 1268 2548 1291
rect 2528 1240 2529 1271
rect 2544 1270 2545 1291
rect 2386 1272 2387 1291
rect 2529 1272 2530 1291
rect 2534 1240 2535 1273
rect 2556 1272 2557 1291
rect 2550 1240 2551 1275
rect 2565 1274 2566 1291
rect 2525 1240 2526 1277
rect 2550 1276 2551 1291
rect 2501 1240 2502 1279
rect 2526 1278 2527 1291
rect 2553 1240 2554 1279
rect 2574 1278 2575 1291
rect 2531 1240 2532 1281
rect 2553 1280 2554 1291
rect 2583 1240 2584 1281
rect 2662 1280 2663 1291
rect 2586 1240 2587 1283
rect 2615 1282 2616 1291
rect 2595 1240 2596 1285
rect 2633 1284 2634 1291
rect 2618 1286 2619 1291
rect 2665 1286 2666 1291
rect 2636 1288 2637 1291
rect 2649 1288 2650 1291
rect 2659 1288 2660 1291
rect 2675 1288 2676 1291
rect 2314 1295 2315 1298
rect 2318 1295 2319 1298
rect 2323 1297 2324 1366
rect 2330 1297 2331 1366
rect 2325 1295 2326 1300
rect 2429 1295 2430 1300
rect 2349 1295 2350 1302
rect 2593 1301 2594 1366
rect 2357 1303 2358 1366
rect 2642 1295 2643 1304
rect 2360 1305 2361 1366
rect 2486 1305 2487 1366
rect 2403 1307 2404 1366
rect 2411 1295 2412 1308
rect 2409 1309 2410 1366
rect 2423 1295 2424 1310
rect 2412 1311 2413 1366
rect 2426 1295 2427 1312
rect 2415 1313 2416 1366
rect 2417 1295 2418 1314
rect 2421 1313 2422 1366
rect 2432 1295 2433 1314
rect 2424 1315 2425 1366
rect 2435 1295 2436 1316
rect 2433 1317 2434 1366
rect 2450 1295 2451 1318
rect 2367 1319 2368 1366
rect 2451 1319 2452 1366
rect 2442 1321 2443 1366
rect 2465 1295 2466 1322
rect 2444 1295 2445 1324
rect 2462 1295 2463 1324
rect 2448 1325 2449 1366
rect 2459 1295 2460 1326
rect 2464 1325 2465 1366
rect 2492 1295 2493 1326
rect 2468 1295 2469 1328
rect 2477 1327 2478 1366
rect 2471 1329 2472 1366
rect 2526 1295 2527 1330
rect 2480 1295 2481 1332
rect 2498 1295 2499 1332
rect 2489 1331 2490 1366
rect 2489 1295 2490 1332
rect 2492 1333 2493 1366
rect 2495 1295 2496 1334
rect 2501 1333 2502 1366
rect 2516 1333 2517 1366
rect 2504 1335 2505 1366
rect 2529 1295 2530 1336
rect 2507 1337 2508 1366
rect 2550 1295 2551 1338
rect 2531 1339 2532 1366
rect 2544 1295 2545 1340
rect 2534 1341 2535 1366
rect 2553 1295 2554 1342
rect 2537 1343 2538 1366
rect 2556 1295 2557 1344
rect 2546 1345 2547 1366
rect 2547 1295 2548 1346
rect 2549 1345 2550 1366
rect 2559 1295 2560 1346
rect 2474 1347 2475 1366
rect 2558 1347 2559 1366
rect 2552 1349 2553 1366
rect 2565 1295 2566 1350
rect 2561 1351 2562 1366
rect 2574 1295 2575 1352
rect 2602 1351 2603 1366
rect 2636 1295 2637 1352
rect 2605 1353 2606 1366
rect 2621 1295 2622 1354
rect 2615 1295 2616 1356
rect 2665 1295 2666 1356
rect 2584 1357 2585 1366
rect 2615 1357 2616 1366
rect 2618 1295 2619 1358
rect 2642 1357 2643 1366
rect 2633 1295 2634 1360
rect 2649 1295 2650 1360
rect 2632 1361 2633 1366
rect 2659 1295 2660 1362
rect 2645 1363 2646 1366
rect 2662 1295 2663 1364
rect 2323 1370 2324 1373
rect 2381 1372 2382 1433
rect 2351 1374 2352 1433
rect 2393 1374 2394 1433
rect 2357 1370 2358 1377
rect 2378 1376 2379 1433
rect 2372 1378 2373 1433
rect 2421 1370 2422 1379
rect 2375 1380 2376 1433
rect 2415 1370 2416 1381
rect 2403 1370 2404 1383
rect 2426 1382 2427 1433
rect 2409 1370 2410 1385
rect 2414 1384 2415 1433
rect 2399 1386 2400 1433
rect 2408 1386 2409 1433
rect 2412 1370 2413 1387
rect 2417 1386 2418 1433
rect 2424 1370 2425 1387
rect 2429 1386 2430 1433
rect 2433 1370 2434 1387
rect 2438 1386 2439 1433
rect 2448 1370 2449 1387
rect 2453 1386 2454 1433
rect 2442 1370 2443 1389
rect 2447 1388 2448 1433
rect 2451 1370 2452 1389
rect 2456 1388 2457 1433
rect 2471 1388 2472 1433
rect 2498 1388 2499 1433
rect 2477 1370 2478 1391
rect 2480 1390 2481 1433
rect 2474 1370 2475 1393
rect 2477 1392 2478 1433
rect 2483 1392 2484 1433
rect 2489 1370 2490 1393
rect 2486 1370 2487 1395
rect 2489 1394 2490 1433
rect 2492 1370 2493 1395
rect 2495 1394 2496 1433
rect 2464 1370 2465 1397
rect 2492 1396 2493 1433
rect 2507 1370 2508 1397
rect 2510 1396 2511 1433
rect 2504 1370 2505 1399
rect 2507 1398 2508 1433
rect 2504 1400 2505 1433
rect 2516 1400 2517 1433
rect 2513 1370 2514 1403
rect 2587 1370 2588 1403
rect 2534 1370 2535 1405
rect 2543 1404 2544 1433
rect 2531 1370 2532 1407
rect 2534 1406 2535 1433
rect 2564 1406 2565 1433
rect 2608 1370 2609 1407
rect 2581 1370 2582 1409
rect 2630 1408 2631 1433
rect 2561 1370 2562 1411
rect 2580 1410 2581 1433
rect 2552 1370 2553 1413
rect 2561 1412 2562 1433
rect 2549 1370 2550 1415
rect 2552 1414 2553 1433
rect 2546 1370 2547 1417
rect 2549 1416 2550 1433
rect 2537 1370 2538 1419
rect 2546 1418 2547 1433
rect 2584 1370 2585 1419
rect 2615 1370 2616 1419
rect 2501 1370 2502 1421
rect 2583 1420 2584 1433
rect 2593 1370 2594 1421
rect 2608 1420 2609 1433
rect 2632 1370 2633 1421
rect 2655 1420 2656 1433
rect 2602 1370 2603 1423
rect 2633 1422 2634 1433
rect 2602 1424 2603 1433
rect 2665 1424 2666 1433
rect 2635 1370 2636 1427
rect 2649 1426 2650 1433
rect 2638 1370 2639 1429
rect 2675 1428 2676 1433
rect 2652 1430 2653 1433
rect 2668 1430 2669 1433
rect 2290 1439 2291 1514
rect 2384 1439 2385 1514
rect 2304 1441 2305 1514
rect 2308 1441 2309 1514
rect 2329 1441 2330 1514
rect 2402 1441 2403 1514
rect 2343 1443 2344 1514
rect 2486 1443 2487 1514
rect 2350 1445 2351 1514
rect 2411 1445 2412 1514
rect 2357 1447 2358 1514
rect 2417 1437 2418 1448
rect 2365 1437 2366 1450
rect 2453 1437 2454 1450
rect 2372 1437 2373 1452
rect 2426 1437 2427 1452
rect 2378 1437 2379 1454
rect 2417 1453 2418 1514
rect 2381 1437 2382 1456
rect 2399 1437 2400 1456
rect 2323 1437 2324 1458
rect 2399 1457 2400 1514
rect 2414 1437 2415 1458
rect 2435 1457 2436 1514
rect 2333 1437 2334 1460
rect 2414 1459 2415 1514
rect 2432 1459 2433 1514
rect 2456 1437 2457 1460
rect 2438 1437 2439 1462
rect 2450 1461 2451 1514
rect 2393 1437 2394 1464
rect 2438 1463 2439 1514
rect 2447 1437 2448 1464
rect 2465 1463 2466 1514
rect 2429 1437 2430 1466
rect 2447 1465 2448 1514
rect 2453 1465 2454 1514
rect 2480 1437 2481 1466
rect 2471 1467 2472 1514
rect 2555 1467 2556 1514
rect 2495 1437 2496 1470
rect 2531 1469 2532 1514
rect 2489 1437 2490 1472
rect 2495 1471 2496 1514
rect 2483 1437 2484 1474
rect 2489 1473 2490 1514
rect 2477 1437 2478 1476
rect 2483 1475 2484 1514
rect 2498 1437 2499 1476
rect 2519 1475 2520 1514
rect 2507 1437 2508 1478
rect 2528 1477 2529 1514
rect 2492 1437 2493 1480
rect 2507 1479 2508 1514
rect 2510 1437 2511 1480
rect 2522 1479 2523 1514
rect 2504 1437 2505 1482
rect 2510 1481 2511 1514
rect 2549 1437 2550 1482
rect 2597 1481 2598 1514
rect 2552 1437 2553 1484
rect 2600 1483 2601 1514
rect 2516 1437 2517 1486
rect 2552 1485 2553 1514
rect 2561 1437 2562 1486
rect 2573 1485 2574 1514
rect 2543 1437 2544 1488
rect 2561 1487 2562 1514
rect 2534 1437 2535 1490
rect 2543 1489 2544 1514
rect 2534 1491 2535 1514
rect 2549 1491 2550 1514
rect 2564 1437 2565 1492
rect 2567 1491 2568 1514
rect 2546 1437 2547 1494
rect 2564 1493 2565 1514
rect 2580 1437 2581 1494
rect 2594 1493 2595 1514
rect 2583 1437 2584 1496
rect 2590 1437 2591 1496
rect 2591 1497 2592 1514
rect 2611 1437 2612 1498
rect 2608 1437 2609 1500
rect 2615 1499 2616 1514
rect 2630 1437 2631 1500
rect 2668 1499 2669 1514
rect 2633 1437 2634 1502
rect 2671 1501 2672 1514
rect 2649 1437 2650 1504
rect 2687 1503 2688 1514
rect 2650 1505 2651 1514
rect 2684 1505 2685 1514
rect 2652 1437 2653 1508
rect 2690 1507 2691 1514
rect 2653 1509 2654 1514
rect 2659 1509 2660 1514
rect 2655 1437 2656 1512
rect 2693 1511 2694 1514
rect 2287 1518 2288 1521
rect 2301 1518 2302 1521
rect 2297 1518 2298 1523
rect 2384 1518 2385 1523
rect 2308 1518 2309 1525
rect 2423 1524 2424 1623
rect 2311 1526 2312 1623
rect 2315 1518 2316 1527
rect 2353 1526 2354 1623
rect 2411 1518 2412 1527
rect 2370 1528 2371 1623
rect 2498 1528 2499 1623
rect 2374 1530 2375 1623
rect 2447 1518 2448 1531
rect 2393 1532 2394 1623
rect 2402 1518 2403 1533
rect 2332 1518 2333 1535
rect 2402 1534 2403 1623
rect 2399 1534 2400 1623
rect 2399 1518 2400 1535
rect 2411 1534 2412 1623
rect 2471 1518 2472 1535
rect 2417 1518 2418 1537
rect 2420 1536 2421 1623
rect 2414 1518 2415 1539
rect 2417 1538 2418 1623
rect 2432 1518 2433 1539
rect 2501 1538 2502 1623
rect 2438 1518 2439 1541
rect 2456 1540 2457 1623
rect 2438 1542 2439 1623
rect 2486 1518 2487 1543
rect 2450 1518 2451 1545
rect 2486 1544 2487 1623
rect 2322 1518 2323 1547
rect 2450 1546 2451 1623
rect 2321 1548 2322 1623
rect 2471 1548 2472 1623
rect 2459 1518 2460 1551
rect 2477 1550 2478 1623
rect 2465 1518 2466 1553
rect 2480 1552 2481 1623
rect 2453 1518 2454 1555
rect 2465 1554 2466 1623
rect 2435 1518 2436 1557
rect 2453 1556 2454 1623
rect 2483 1518 2484 1557
rect 2524 1556 2525 1623
rect 2489 1518 2490 1559
rect 2504 1558 2505 1623
rect 2367 1518 2368 1561
rect 2489 1560 2490 1623
rect 2367 1562 2368 1623
rect 2492 1562 2493 1623
rect 2495 1518 2496 1563
rect 2536 1562 2537 1623
rect 2510 1518 2511 1565
rect 2513 1518 2514 1565
rect 2507 1518 2508 1567
rect 2514 1566 2515 1623
rect 2507 1568 2508 1623
rect 2706 1568 2707 1623
rect 2519 1518 2520 1571
rect 2557 1570 2558 1623
rect 2522 1518 2523 1573
rect 2569 1572 2570 1623
rect 2528 1518 2529 1575
rect 2575 1574 2576 1623
rect 2360 1576 2361 1623
rect 2527 1576 2528 1623
rect 2534 1518 2535 1577
rect 2539 1576 2540 1623
rect 2543 1518 2544 1577
rect 2696 1518 2697 1577
rect 2531 1518 2532 1579
rect 2542 1578 2543 1623
rect 2552 1518 2553 1579
rect 2581 1578 2582 1623
rect 2567 1518 2568 1581
rect 2611 1580 2612 1623
rect 2573 1518 2574 1583
rect 2617 1582 2618 1623
rect 2578 1584 2579 1623
rect 2585 1518 2586 1585
rect 2591 1518 2592 1585
rect 2608 1584 2609 1623
rect 2594 1518 2595 1587
rect 2629 1586 2630 1623
rect 2597 1518 2598 1589
rect 2623 1588 2624 1623
rect 2561 1518 2562 1591
rect 2596 1590 2597 1623
rect 2560 1592 2561 1623
rect 2625 1518 2626 1593
rect 2600 1518 2601 1595
rect 2626 1594 2627 1623
rect 2564 1518 2565 1597
rect 2599 1596 2600 1623
rect 2615 1518 2616 1597
rect 2664 1596 2665 1623
rect 2653 1518 2654 1599
rect 2658 1598 2659 1623
rect 2656 1518 2657 1601
rect 2709 1600 2710 1623
rect 2668 1518 2669 1603
rect 2700 1602 2701 1623
rect 2671 1518 2672 1605
rect 2703 1604 2704 1623
rect 2670 1606 2671 1623
rect 2697 1606 2698 1623
rect 2685 1608 2686 1623
rect 2779 1608 2780 1623
rect 2687 1518 2688 1611
rect 2718 1610 2719 1623
rect 2690 1518 2691 1613
rect 2721 1612 2722 1623
rect 2693 1518 2694 1615
rect 2744 1614 2745 1623
rect 2650 1518 2651 1617
rect 2694 1616 2695 1623
rect 2649 1618 2650 1623
rect 2667 1618 2668 1623
rect 2724 1618 2725 1623
rect 2792 1618 2793 1623
rect 2765 1620 2766 1623
rect 2772 1620 2773 1623
rect 2311 1627 2312 1630
rect 2450 1627 2451 1630
rect 2312 1631 2313 1718
rect 2423 1627 2424 1632
rect 2325 1627 2326 1634
rect 2510 1633 2511 1718
rect 2326 1635 2327 1718
rect 2646 1627 2647 1636
rect 2340 1637 2341 1718
rect 2411 1637 2412 1718
rect 2353 1627 2354 1640
rect 2367 1627 2368 1640
rect 2368 1641 2369 1718
rect 2498 1627 2499 1642
rect 2375 1643 2376 1718
rect 2489 1627 2490 1644
rect 2393 1643 2394 1718
rect 2393 1627 2394 1644
rect 2399 1643 2400 1718
rect 2399 1627 2400 1644
rect 2402 1643 2403 1718
rect 2402 1627 2403 1644
rect 2414 1645 2415 1718
rect 2516 1645 2517 1718
rect 2420 1627 2421 1648
rect 2423 1647 2424 1718
rect 2417 1627 2418 1650
rect 2420 1649 2421 1718
rect 2417 1651 2418 1718
rect 2492 1627 2493 1652
rect 2438 1627 2439 1654
rect 2450 1653 2451 1718
rect 2453 1627 2454 1654
rect 2462 1653 2463 1718
rect 2459 1627 2460 1656
rect 2581 1627 2582 1656
rect 2319 1657 2320 1718
rect 2459 1657 2460 1718
rect 2465 1627 2466 1658
rect 2474 1657 2475 1718
rect 2456 1627 2457 1660
rect 2465 1659 2466 1718
rect 2314 1627 2315 1662
rect 2456 1661 2457 1718
rect 2480 1627 2481 1662
rect 2495 1661 2496 1718
rect 2471 1627 2472 1664
rect 2480 1663 2481 1718
rect 2483 1663 2484 1718
rect 2501 1627 2502 1664
rect 2384 1627 2385 1666
rect 2501 1665 2502 1718
rect 2486 1627 2487 1668
rect 2492 1667 2493 1718
rect 2507 1667 2508 1718
rect 2778 1667 2779 1718
rect 2518 1627 2519 1670
rect 2546 1669 2547 1718
rect 2522 1671 2523 1718
rect 2524 1627 2525 1672
rect 2525 1673 2526 1718
rect 2527 1627 2528 1674
rect 2531 1673 2532 1718
rect 2534 1673 2535 1718
rect 2539 1627 2540 1674
rect 2681 1673 2682 1718
rect 2536 1627 2537 1676
rect 2540 1675 2541 1718
rect 2477 1627 2478 1678
rect 2537 1677 2538 1718
rect 2542 1627 2543 1678
rect 2543 1677 2544 1718
rect 2552 1677 2553 1718
rect 2560 1627 2561 1678
rect 2557 1627 2558 1680
rect 2567 1679 2568 1718
rect 2569 1627 2570 1680
rect 2573 1679 2574 1718
rect 2570 1681 2571 1718
rect 2575 1627 2576 1682
rect 2578 1627 2579 1682
rect 2591 1681 2592 1718
rect 2564 1683 2565 1718
rect 2579 1683 2580 1718
rect 2599 1627 2600 1684
rect 2603 1683 2604 1718
rect 2596 1627 2597 1686
rect 2600 1685 2601 1718
rect 2608 1627 2609 1686
rect 2642 1685 2643 1718
rect 2611 1627 2612 1688
rect 2612 1687 2613 1718
rect 2617 1627 2618 1688
rect 2618 1687 2619 1718
rect 2626 1627 2627 1688
rect 2633 1687 2634 1718
rect 2629 1627 2630 1690
rect 2636 1689 2637 1718
rect 2623 1627 2624 1692
rect 2630 1691 2631 1718
rect 2639 1691 2640 1718
rect 2771 1691 2772 1718
rect 2651 1693 2652 1718
rect 2721 1627 2722 1694
rect 2660 1695 2661 1718
rect 2664 1627 2665 1696
rect 2675 1695 2676 1718
rect 2730 1627 2731 1696
rect 2684 1697 2685 1718
rect 2685 1627 2686 1698
rect 2697 1627 2698 1698
rect 2740 1697 2741 1718
rect 2694 1627 2695 1700
rect 2696 1699 2697 1718
rect 2693 1701 2694 1718
rect 2755 1627 2756 1702
rect 2700 1627 2701 1704
rect 2751 1627 2752 1704
rect 2658 1627 2659 1706
rect 2699 1705 2700 1718
rect 2703 1627 2704 1706
rect 2711 1705 2712 1718
rect 2706 1627 2707 1708
rect 2720 1707 2721 1718
rect 2718 1627 2719 1710
rect 2734 1627 2735 1710
rect 2724 1627 2725 1712
rect 2786 1627 2787 1712
rect 2709 1627 2710 1714
rect 2723 1713 2724 1718
rect 2708 1715 2709 1718
rect 2748 1627 2749 1716
rect 2792 1627 2793 1716
rect 2799 1627 2800 1716
rect 2305 1722 2306 1725
rect 2306 1724 2307 1827
rect 2312 1722 2313 1725
rect 2459 1722 2460 1725
rect 2323 1726 2324 1827
rect 2330 1726 2331 1827
rect 2326 1722 2327 1729
rect 2453 1728 2454 1827
rect 2341 1730 2342 1827
rect 2444 1730 2445 1827
rect 2369 1732 2370 1827
rect 2474 1722 2475 1733
rect 2375 1722 2376 1735
rect 2426 1734 2427 1827
rect 2393 1734 2394 1827
rect 2393 1722 2394 1735
rect 2399 1734 2400 1827
rect 2399 1722 2400 1735
rect 2411 1734 2412 1827
rect 2411 1722 2412 1735
rect 2417 1722 2418 1737
rect 2501 1722 2502 1737
rect 2420 1736 2421 1827
rect 2420 1722 2421 1737
rect 2423 1736 2424 1827
rect 2423 1722 2424 1737
rect 2447 1738 2448 1827
rect 2462 1722 2463 1739
rect 2450 1722 2451 1741
rect 2462 1740 2463 1827
rect 2417 1742 2418 1827
rect 2450 1742 2451 1827
rect 2456 1722 2457 1743
rect 2459 1742 2460 1827
rect 2402 1722 2403 1745
rect 2456 1744 2457 1827
rect 2465 1722 2466 1745
rect 2468 1744 2469 1827
rect 2471 1722 2472 1745
rect 2516 1744 2517 1827
rect 2474 1746 2475 1827
rect 2480 1722 2481 1747
rect 2477 1748 2478 1827
rect 2483 1722 2484 1749
rect 2486 1748 2487 1827
rect 2495 1722 2496 1749
rect 2492 1748 2493 1827
rect 2492 1722 2493 1749
rect 2501 1748 2502 1827
rect 2510 1722 2511 1749
rect 2355 1750 2356 1827
rect 2510 1750 2511 1827
rect 2507 1722 2508 1753
rect 2513 1752 2514 1827
rect 2299 1754 2300 1827
rect 2507 1754 2508 1827
rect 2537 1722 2538 1755
rect 2549 1754 2550 1827
rect 2525 1722 2526 1757
rect 2537 1756 2538 1827
rect 2543 1722 2544 1757
rect 2561 1756 2562 1827
rect 2552 1722 2553 1759
rect 2579 1758 2580 1827
rect 2558 1760 2559 1827
rect 2760 1760 2761 1827
rect 2564 1722 2565 1763
rect 2576 1762 2577 1827
rect 2546 1722 2547 1765
rect 2564 1764 2565 1827
rect 2534 1722 2535 1767
rect 2546 1766 2547 1827
rect 2522 1722 2523 1769
rect 2534 1768 2535 1827
rect 2522 1770 2523 1827
rect 2540 1722 2541 1771
rect 2567 1722 2568 1771
rect 2582 1770 2583 1827
rect 2573 1722 2574 1773
rect 2594 1772 2595 1827
rect 2591 1722 2592 1775
rect 2606 1774 2607 1827
rect 2603 1722 2604 1777
rect 2715 1776 2716 1827
rect 2570 1722 2571 1779
rect 2603 1778 2604 1827
rect 2630 1722 2631 1779
rect 2654 1722 2655 1779
rect 2630 1780 2631 1827
rect 2657 1780 2658 1827
rect 2633 1722 2634 1783
rect 2687 1782 2688 1827
rect 2612 1722 2613 1785
rect 2633 1784 2634 1827
rect 2639 1722 2640 1785
rect 2669 1784 2670 1827
rect 2618 1722 2619 1787
rect 2639 1786 2640 1827
rect 2651 1722 2652 1787
rect 2736 1786 2737 1827
rect 2636 1722 2637 1789
rect 2651 1788 2652 1827
rect 2672 1722 2673 1789
rect 2681 1722 2682 1789
rect 2642 1722 2643 1791
rect 2672 1790 2673 1827
rect 2660 1722 2661 1793
rect 2681 1792 2682 1827
rect 2600 1722 2601 1795
rect 2660 1794 2661 1827
rect 2600 1796 2601 1827
rect 2645 1722 2646 1797
rect 2675 1722 2676 1797
rect 2705 1722 2706 1797
rect 2684 1722 2685 1799
rect 2739 1798 2740 1827
rect 2627 1800 2628 1827
rect 2684 1800 2685 1827
rect 2693 1722 2694 1801
rect 2751 1800 2752 1827
rect 2696 1722 2697 1803
rect 2766 1802 2767 1827
rect 2696 1804 2697 1827
rect 2819 1804 2820 1827
rect 2699 1722 2700 1807
rect 2769 1806 2770 1827
rect 2708 1722 2709 1809
rect 2778 1808 2779 1827
rect 2528 1810 2529 1827
rect 2708 1810 2709 1827
rect 2711 1722 2712 1811
rect 2781 1810 2782 1827
rect 2720 1722 2721 1813
rect 2796 1812 2797 1827
rect 2702 1722 2703 1815
rect 2721 1814 2722 1827
rect 2723 1722 2724 1815
rect 2784 1814 2785 1827
rect 2729 1722 2730 1817
rect 2799 1816 2800 1827
rect 2733 1818 2734 1827
rect 2771 1722 2772 1819
rect 2724 1820 2725 1827
rect 2772 1820 2773 1827
rect 2742 1822 2743 1827
rect 2747 1722 2748 1823
rect 2754 1822 2755 1827
rect 2812 1822 2813 1827
rect 2757 1824 2758 1827
rect 2809 1824 2810 1827
rect 2302 1831 2303 1834
rect 2306 1831 2307 1834
rect 2316 1831 2317 1834
rect 2459 1831 2460 1834
rect 2320 1835 2321 1942
rect 2442 1835 2443 1942
rect 2330 1831 2331 1838
rect 2406 1837 2407 1942
rect 2337 1831 2338 1840
rect 2423 1831 2424 1840
rect 2358 1831 2359 1842
rect 2687 1831 2688 1842
rect 2362 1831 2363 1844
rect 2781 1831 2782 1844
rect 2381 1831 2382 1846
rect 2393 1831 2394 1846
rect 2391 1847 2392 1942
rect 2399 1831 2400 1848
rect 2403 1847 2404 1942
rect 2411 1831 2412 1848
rect 2412 1849 2413 1942
rect 2528 1831 2529 1850
rect 2415 1851 2416 1942
rect 2532 1851 2533 1942
rect 2418 1853 2419 1942
rect 2420 1831 2421 1854
rect 2433 1853 2434 1942
rect 2462 1831 2463 1854
rect 2439 1855 2440 1942
rect 2444 1831 2445 1856
rect 2456 1831 2457 1856
rect 2460 1855 2461 1942
rect 2453 1831 2454 1858
rect 2457 1857 2458 1942
rect 2450 1831 2451 1860
rect 2454 1859 2455 1942
rect 2447 1831 2448 1862
rect 2451 1861 2452 1942
rect 2469 1861 2470 1942
rect 2523 1861 2524 1942
rect 2474 1831 2475 1864
rect 2475 1863 2476 1942
rect 2477 1831 2478 1864
rect 2478 1863 2479 1942
rect 2481 1863 2482 1942
rect 2486 1831 2487 1864
rect 2487 1865 2488 1942
rect 2501 1831 2502 1866
rect 2492 1831 2493 1868
rect 2499 1867 2500 1942
rect 2493 1869 2494 1942
rect 2516 1831 2517 1870
rect 2471 1831 2472 1872
rect 2517 1871 2518 1942
rect 2537 1831 2538 1872
rect 2541 1871 2542 1942
rect 2534 1831 2535 1874
rect 2538 1873 2539 1942
rect 2544 1873 2545 1942
rect 2561 1831 2562 1874
rect 2549 1831 2550 1876
rect 2553 1875 2554 1942
rect 2546 1831 2547 1878
rect 2550 1877 2551 1942
rect 2556 1877 2557 1942
rect 2558 1831 2559 1878
rect 2313 1831 2314 1880
rect 2559 1879 2560 1942
rect 2564 1831 2565 1880
rect 2574 1879 2575 1942
rect 2579 1831 2580 1880
rect 2580 1879 2581 1942
rect 2600 1831 2601 1880
rect 2693 1831 2694 1880
rect 2603 1831 2604 1882
rect 2613 1881 2614 1942
rect 2604 1883 2605 1942
rect 2676 1883 2677 1942
rect 2610 1885 2611 1942
rect 2690 1831 2691 1886
rect 2594 1831 2595 1888
rect 2691 1887 2692 1942
rect 2627 1831 2628 1890
rect 2631 1889 2632 1942
rect 2606 1831 2607 1892
rect 2628 1891 2629 1942
rect 2576 1831 2577 1894
rect 2607 1893 2608 1942
rect 2651 1831 2652 1894
rect 2744 1893 2745 1942
rect 2657 1831 2658 1896
rect 2658 1895 2659 1942
rect 2660 1831 2661 1896
rect 2661 1895 2662 1942
rect 2669 1831 2670 1896
rect 2670 1895 2671 1942
rect 2672 1831 2673 1896
rect 2673 1895 2674 1942
rect 2681 1831 2682 1896
rect 2694 1895 2695 1942
rect 2684 1831 2685 1898
rect 2688 1897 2689 1942
rect 2696 1831 2697 1898
rect 2781 1897 2782 1942
rect 2711 1831 2712 1900
rect 2742 1831 2743 1900
rect 2714 1901 2715 1942
rect 2763 1831 2764 1902
rect 2717 1903 2718 1942
rect 2721 1831 2722 1904
rect 2720 1905 2721 1942
rect 2733 1831 2734 1906
rect 2724 1831 2725 1908
rect 2759 1907 2760 1942
rect 2723 1909 2724 1942
rect 2736 1831 2737 1910
rect 2726 1911 2727 1942
rect 2739 1831 2740 1912
rect 2729 1913 2730 1942
rect 2833 1831 2834 1914
rect 2741 1915 2742 1942
rect 2754 1831 2755 1916
rect 2751 1831 2752 1918
rect 2771 1917 2772 1942
rect 2753 1919 2754 1942
rect 2766 1831 2767 1920
rect 2757 1831 2758 1922
rect 2762 1921 2763 1942
rect 2639 1831 2640 1924
rect 2756 1923 2757 1942
rect 2633 1831 2634 1926
rect 2640 1925 2641 1942
rect 2765 1925 2766 1942
rect 2796 1831 2797 1926
rect 2769 1831 2770 1928
rect 2816 1831 2817 1928
rect 2768 1929 2769 1942
rect 2819 1831 2820 1930
rect 2778 1831 2779 1932
rect 2847 1831 2848 1932
rect 2777 1933 2778 1942
rect 2812 1831 2813 1934
rect 2732 1935 2733 1942
rect 2812 1935 2813 1942
rect 2784 1831 2785 1938
rect 2802 1831 2803 1938
rect 2799 1831 2800 1940
rect 2805 1831 2806 1940
rect 2302 1948 2303 2077
rect 2426 1948 2427 2077
rect 2309 1950 2310 2077
rect 2429 1950 2430 2077
rect 2317 1946 2318 1953
rect 2389 1952 2390 2077
rect 2320 1946 2321 1955
rect 2445 1946 2446 1955
rect 2324 1946 2325 1957
rect 2400 1946 2401 1957
rect 2323 1958 2324 2077
rect 2495 1958 2496 2077
rect 2345 1946 2346 1961
rect 2514 1946 2515 1961
rect 2348 1946 2349 1963
rect 2691 1946 2692 1963
rect 2359 1946 2360 1965
rect 2546 1964 2547 2077
rect 2366 1946 2367 1967
rect 2391 1946 2392 1967
rect 2397 1946 2398 1967
rect 2532 1946 2533 1967
rect 2403 1946 2404 1969
rect 2501 1968 2502 2077
rect 2402 1970 2403 2077
rect 2460 1946 2461 1971
rect 2406 1946 2407 1973
rect 2420 1972 2421 2077
rect 2439 1946 2440 1973
rect 2459 1972 2460 2077
rect 2418 1946 2419 1975
rect 2438 1974 2439 2077
rect 2465 1974 2466 2077
rect 2550 1946 2551 1975
rect 2469 1946 2470 1977
rect 2622 1946 2623 1977
rect 2478 1946 2479 1979
rect 2513 1978 2514 2077
rect 2454 1946 2455 1981
rect 2477 1980 2478 2077
rect 2433 1946 2434 1983
rect 2453 1982 2454 2077
rect 2380 1984 2381 2077
rect 2432 1984 2433 2077
rect 2487 1946 2488 1985
rect 2528 1984 2529 2077
rect 2493 1946 2494 1987
rect 2534 1986 2535 2077
rect 2457 1946 2458 1989
rect 2492 1988 2493 2077
rect 2508 1946 2509 1989
rect 2549 1988 2550 2077
rect 2442 1946 2443 1991
rect 2507 1990 2508 2077
rect 2351 1992 2352 2077
rect 2441 1992 2442 2077
rect 2517 1946 2518 1993
rect 2565 1946 2566 1993
rect 2504 1994 2505 2077
rect 2516 1994 2517 2077
rect 2523 1946 2524 1995
rect 2567 1994 2568 2077
rect 2481 1946 2482 1997
rect 2522 1996 2523 2077
rect 2538 1946 2539 1997
rect 2570 1996 2571 2077
rect 2537 1998 2538 2077
rect 2553 1946 2554 1999
rect 2544 1946 2545 2001
rect 2576 2000 2577 2077
rect 2499 1946 2500 2003
rect 2543 2002 2544 2077
rect 2337 2004 2338 2077
rect 2498 2004 2499 2077
rect 2556 1946 2557 2005
rect 2582 2004 2583 2077
rect 2559 1946 2560 2007
rect 2585 2006 2586 2077
rect 2564 2008 2565 2077
rect 2697 1946 2698 2009
rect 2574 1946 2575 2011
rect 2600 2010 2601 2077
rect 2541 1946 2542 2013
rect 2573 2012 2574 2077
rect 2511 1946 2512 2015
rect 2540 2014 2541 2077
rect 2475 1946 2476 2017
rect 2510 2016 2511 2077
rect 2451 1946 2452 2019
rect 2474 2018 2475 2077
rect 2604 1946 2605 2019
rect 2625 1946 2626 2019
rect 2610 1946 2611 2021
rect 2642 2020 2643 2077
rect 2613 1946 2614 2023
rect 2645 2022 2646 2077
rect 2607 1946 2608 2025
rect 2612 2024 2613 2077
rect 2580 1946 2581 2027
rect 2606 2026 2607 2077
rect 2615 2026 2616 2077
rect 2778 2026 2779 2077
rect 2628 1946 2629 2029
rect 2654 2028 2655 2077
rect 2648 2030 2649 2077
rect 2661 1946 2662 2031
rect 2640 1946 2641 2033
rect 2660 2032 2661 2077
rect 2658 1946 2659 2035
rect 2705 2034 2706 2077
rect 2631 1946 2632 2037
rect 2657 2036 2658 2077
rect 2670 1946 2671 2037
rect 2696 2036 2697 2077
rect 2673 1946 2674 2039
rect 2699 2038 2700 2077
rect 2672 2040 2673 2077
rect 2797 2040 2798 2077
rect 2694 1946 2695 2043
rect 2714 2042 2715 2077
rect 2702 2044 2703 2077
rect 2851 2044 2852 2077
rect 2708 2046 2709 2077
rect 2723 1946 2724 2047
rect 2720 1946 2721 2049
rect 2748 2048 2749 2077
rect 2676 1946 2677 2051
rect 2720 2050 2721 2077
rect 2726 1946 2727 2051
rect 2763 2050 2764 2077
rect 2729 1946 2730 2053
rect 2760 2052 2761 2077
rect 2732 1946 2733 2055
rect 2805 1946 2806 2055
rect 2636 2056 2637 2077
rect 2732 2056 2733 2077
rect 2751 2056 2752 2077
rect 2845 2056 2846 2077
rect 2765 1946 2766 2059
rect 2794 2058 2795 2077
rect 2768 1946 2769 2061
rect 2791 2060 2792 2077
rect 2771 1946 2772 2063
rect 2774 1946 2775 2063
rect 2753 1946 2754 2065
rect 2772 2064 2773 2077
rect 2741 1946 2742 2067
rect 2754 2066 2755 2077
rect 2756 1946 2757 2067
rect 2775 2066 2776 2077
rect 2744 1946 2745 2069
rect 2757 2068 2758 2077
rect 2717 1946 2718 2071
rect 2745 2070 2746 2077
rect 2688 1946 2689 2073
rect 2717 2072 2718 2077
rect 2812 1946 2813 2073
rect 2816 1946 2817 2073
rect 2817 2074 2818 2077
rect 2824 2074 2825 2077
rect 2294 2083 2295 2200
rect 2456 2083 2457 2200
rect 2301 2085 2302 2200
rect 2426 2081 2427 2086
rect 2306 2081 2307 2088
rect 2462 2087 2463 2200
rect 2315 2089 2316 2200
rect 2429 2081 2430 2090
rect 2308 2091 2309 2200
rect 2429 2091 2430 2200
rect 2324 2093 2325 2200
rect 2516 2093 2517 2200
rect 2344 2081 2345 2096
rect 2441 2081 2442 2096
rect 2351 2081 2352 2098
rect 2432 2081 2433 2098
rect 2299 2081 2300 2100
rect 2432 2099 2433 2200
rect 2347 2081 2348 2102
rect 2350 2101 2351 2200
rect 2357 2101 2358 2200
rect 2477 2081 2478 2102
rect 2375 2103 2376 2200
rect 2495 2081 2496 2104
rect 2377 2081 2378 2106
rect 2507 2081 2508 2106
rect 2392 2081 2393 2108
rect 2567 2081 2568 2108
rect 2336 2109 2337 2200
rect 2393 2109 2394 2200
rect 2396 2081 2397 2110
rect 2537 2081 2538 2110
rect 2399 2111 2400 2200
rect 2420 2081 2421 2112
rect 2402 2081 2403 2114
rect 2486 2113 2487 2200
rect 2414 2115 2415 2200
rect 2552 2115 2553 2200
rect 2438 2081 2439 2118
rect 2519 2117 2520 2200
rect 2447 2119 2448 2200
rect 2459 2081 2460 2120
rect 2287 2121 2288 2200
rect 2459 2121 2460 2200
rect 2453 2081 2454 2124
rect 2477 2123 2478 2200
rect 2471 2125 2472 2200
rect 2474 2081 2475 2126
rect 2354 2081 2355 2128
rect 2474 2127 2475 2200
rect 2483 2127 2484 2200
rect 2492 2081 2493 2128
rect 2489 2129 2490 2200
rect 2498 2081 2499 2130
rect 2501 2081 2502 2130
rect 2507 2129 2508 2200
rect 2501 2131 2502 2200
rect 2504 2081 2505 2132
rect 2275 2133 2276 2200
rect 2504 2133 2505 2200
rect 2510 2133 2511 2200
rect 2510 2081 2511 2134
rect 2513 2133 2514 2200
rect 2513 2081 2514 2134
rect 2522 2133 2523 2200
rect 2522 2081 2523 2134
rect 2528 2081 2529 2134
rect 2558 2133 2559 2200
rect 2534 2081 2535 2136
rect 2555 2135 2556 2200
rect 2534 2137 2535 2200
rect 2543 2081 2544 2138
rect 2537 2139 2538 2200
rect 2546 2081 2547 2140
rect 2540 2139 2541 2200
rect 2540 2081 2541 2140
rect 2549 2139 2550 2200
rect 2549 2081 2550 2140
rect 2564 2081 2565 2140
rect 2567 2139 2568 2200
rect 2570 2139 2571 2200
rect 2570 2081 2571 2140
rect 2573 2139 2574 2200
rect 2573 2081 2574 2140
rect 2576 2081 2577 2140
rect 2627 2139 2628 2200
rect 2582 2139 2583 2200
rect 2582 2081 2583 2140
rect 2585 2081 2586 2142
rect 2591 2141 2592 2200
rect 2588 2143 2589 2200
rect 2879 2143 2880 2200
rect 2594 2145 2595 2200
rect 2600 2081 2601 2146
rect 2606 2081 2607 2146
rect 2630 2081 2631 2146
rect 2606 2147 2607 2200
rect 2612 2081 2613 2148
rect 2609 2149 2610 2200
rect 2615 2081 2616 2150
rect 2630 2149 2631 2200
rect 2739 2081 2740 2150
rect 2639 2151 2640 2200
rect 2645 2081 2646 2152
rect 2654 2081 2655 2152
rect 2666 2151 2667 2200
rect 2654 2153 2655 2200
rect 2660 2081 2661 2154
rect 2657 2081 2658 2156
rect 2732 2081 2733 2156
rect 2669 2157 2670 2200
rect 2723 2157 2724 2200
rect 2672 2081 2673 2160
rect 2770 2159 2771 2200
rect 2672 2161 2673 2200
rect 2817 2081 2818 2162
rect 2684 2163 2685 2200
rect 2757 2081 2758 2164
rect 2699 2081 2700 2166
rect 2711 2165 2712 2200
rect 2705 2081 2706 2168
rect 2720 2167 2721 2200
rect 2714 2167 2715 2200
rect 2714 2081 2715 2168
rect 2717 2081 2718 2170
rect 2729 2169 2730 2200
rect 2702 2081 2703 2172
rect 2717 2171 2718 2200
rect 2735 2081 2736 2172
rect 2782 2171 2783 2200
rect 2742 2171 2743 2200
rect 2742 2081 2743 2172
rect 2751 2081 2752 2174
rect 2824 2081 2825 2174
rect 2748 2081 2749 2176
rect 2752 2175 2753 2200
rect 2754 2081 2755 2176
rect 2767 2175 2768 2200
rect 2708 2081 2709 2178
rect 2755 2177 2756 2200
rect 2696 2081 2697 2180
rect 2708 2179 2709 2200
rect 2696 2181 2697 2200
rect 2807 2081 2808 2182
rect 2763 2081 2764 2184
rect 2837 2183 2838 2200
rect 2760 2081 2761 2186
rect 2764 2185 2765 2200
rect 2772 2081 2773 2186
rect 2785 2185 2786 2200
rect 2745 2081 2746 2188
rect 2773 2187 2774 2200
rect 2636 2081 2637 2190
rect 2746 2189 2747 2200
rect 2636 2191 2637 2200
rect 2642 2081 2643 2192
rect 2642 2193 2643 2200
rect 2648 2081 2649 2194
rect 2775 2081 2776 2194
rect 2788 2193 2789 2200
rect 2791 2081 2792 2194
rect 2804 2193 2805 2200
rect 2794 2081 2795 2196
rect 2807 2195 2808 2200
rect 2797 2081 2798 2198
rect 2810 2197 2811 2200
rect 2816 2197 2817 2200
rect 2820 2197 2821 2200
rect 2840 2197 2841 2200
rect 2876 2197 2877 2200
rect 2288 2206 2289 2343
rect 2456 2204 2457 2207
rect 2291 2208 2292 2343
rect 2436 2208 2437 2343
rect 2301 2204 2302 2211
rect 2429 2204 2430 2211
rect 2304 2204 2305 2213
rect 2462 2204 2463 2213
rect 2305 2214 2306 2343
rect 2457 2214 2458 2343
rect 2309 2216 2310 2343
rect 2432 2204 2433 2217
rect 2318 2218 2319 2343
rect 2499 2218 2500 2343
rect 2333 2204 2334 2221
rect 2486 2204 2487 2221
rect 2343 2222 2344 2343
rect 2489 2204 2490 2223
rect 2357 2224 2358 2343
rect 2532 2224 2533 2343
rect 2369 2226 2370 2343
rect 2510 2204 2511 2227
rect 2372 2228 2373 2343
rect 2552 2204 2553 2229
rect 2378 2204 2379 2231
rect 2474 2204 2475 2231
rect 2382 2232 2383 2343
rect 2507 2204 2508 2233
rect 2388 2234 2389 2343
rect 2393 2204 2394 2235
rect 2399 2204 2400 2235
rect 2469 2234 2470 2343
rect 2329 2236 2330 2343
rect 2400 2236 2401 2343
rect 2439 2236 2440 2343
rect 2459 2204 2460 2237
rect 2322 2238 2323 2343
rect 2460 2238 2461 2343
rect 2445 2240 2446 2343
rect 2544 2240 2545 2343
rect 2447 2204 2448 2243
rect 2448 2242 2449 2343
rect 2466 2242 2467 2343
rect 2483 2204 2484 2243
rect 2471 2204 2472 2245
rect 2472 2244 2473 2343
rect 2475 2244 2476 2343
rect 2537 2204 2538 2245
rect 2487 2246 2488 2343
rect 2501 2204 2502 2247
rect 2493 2248 2494 2343
rect 2504 2204 2505 2249
rect 2477 2204 2478 2251
rect 2505 2250 2506 2343
rect 2495 2204 2496 2253
rect 2502 2252 2503 2343
rect 2350 2204 2351 2255
rect 2496 2254 2497 2343
rect 2511 2254 2512 2343
rect 2516 2204 2517 2255
rect 2513 2204 2514 2257
rect 2547 2256 2548 2343
rect 2514 2258 2515 2343
rect 2519 2204 2520 2259
rect 2522 2204 2523 2259
rect 2538 2258 2539 2343
rect 2523 2260 2524 2343
rect 2779 2260 2780 2343
rect 2529 2262 2530 2343
rect 2534 2204 2535 2263
rect 2535 2264 2536 2343
rect 2540 2204 2541 2265
rect 2558 2204 2559 2265
rect 2562 2264 2563 2343
rect 2555 2204 2556 2267
rect 2559 2266 2560 2343
rect 2549 2204 2550 2269
rect 2556 2268 2557 2343
rect 2565 2268 2566 2343
rect 2570 2204 2571 2269
rect 2567 2204 2568 2271
rect 2577 2270 2578 2343
rect 2568 2272 2569 2343
rect 2573 2204 2574 2273
rect 2582 2204 2583 2273
rect 2619 2272 2620 2343
rect 2588 2204 2589 2275
rect 2598 2274 2599 2343
rect 2591 2204 2592 2277
rect 2601 2276 2602 2343
rect 2592 2278 2593 2343
rect 2609 2204 2610 2279
rect 2594 2204 2595 2281
rect 2595 2280 2596 2343
rect 2604 2280 2605 2343
rect 2656 2280 2657 2343
rect 2623 2282 2624 2343
rect 2732 2204 2733 2283
rect 2626 2284 2627 2343
rect 2630 2204 2631 2285
rect 2629 2286 2630 2343
rect 2636 2204 2637 2287
rect 2632 2288 2633 2343
rect 2642 2204 2643 2289
rect 2639 2204 2640 2291
rect 2692 2290 2693 2343
rect 2638 2292 2639 2343
rect 2666 2204 2667 2293
rect 2641 2294 2642 2343
rect 2669 2204 2670 2295
rect 2644 2296 2645 2343
rect 2654 2204 2655 2297
rect 2672 2204 2673 2297
rect 2823 2204 2824 2297
rect 2680 2298 2681 2343
rect 2717 2204 2718 2299
rect 2606 2204 2607 2301
rect 2717 2300 2718 2343
rect 2684 2204 2685 2303
rect 2723 2302 2724 2343
rect 2683 2304 2684 2343
rect 2720 2204 2721 2305
rect 2696 2204 2697 2307
rect 2813 2204 2814 2307
rect 2698 2308 2699 2343
rect 2714 2204 2715 2309
rect 2701 2310 2702 2343
rect 2791 2204 2792 2311
rect 2704 2312 2705 2343
rect 2711 2204 2712 2313
rect 2708 2204 2709 2315
rect 2738 2314 2739 2343
rect 2707 2316 2708 2343
rect 2729 2204 2730 2317
rect 2720 2318 2721 2343
rect 2770 2204 2771 2319
rect 2726 2320 2727 2343
rect 2773 2204 2774 2321
rect 2729 2322 2730 2343
rect 2752 2204 2753 2323
rect 2732 2324 2733 2343
rect 2755 2204 2756 2325
rect 2735 2326 2736 2343
rect 2764 2204 2765 2327
rect 2744 2328 2745 2343
rect 2782 2204 2783 2329
rect 2753 2330 2754 2343
rect 2785 2204 2786 2331
rect 2756 2332 2757 2343
rect 2788 2204 2789 2333
rect 2759 2334 2760 2343
rect 2807 2204 2808 2335
rect 2762 2336 2763 2343
rect 2810 2204 2811 2337
rect 2767 2204 2768 2339
rect 2790 2338 2791 2343
rect 2797 2338 2798 2343
rect 2804 2204 2805 2339
rect 2807 2338 2808 2343
rect 2853 2204 2854 2339
rect 2810 2340 2811 2343
rect 2840 2204 2841 2341
rect 2859 2204 2860 2341
rect 2863 2204 2864 2341
rect 2866 2204 2867 2341
rect 2870 2204 2871 2341
rect 2281 2347 2282 2350
rect 2339 2349 2340 2482
rect 2288 2347 2289 2352
rect 2439 2347 2440 2352
rect 2291 2347 2292 2354
rect 2305 2347 2306 2354
rect 2290 2355 2291 2482
rect 2436 2347 2437 2356
rect 2295 2347 2296 2358
rect 2302 2347 2303 2358
rect 2312 2347 2313 2358
rect 2348 2357 2349 2482
rect 2332 2347 2333 2360
rect 2511 2347 2512 2360
rect 2345 2361 2346 2482
rect 2406 2361 2407 2482
rect 2353 2347 2354 2364
rect 2481 2363 2482 2482
rect 2382 2347 2383 2366
rect 2418 2365 2419 2482
rect 2385 2367 2386 2482
rect 2544 2347 2545 2368
rect 2388 2347 2389 2370
rect 2436 2369 2437 2482
rect 2430 2371 2431 2482
rect 2469 2347 2470 2372
rect 2445 2347 2446 2374
rect 2466 2347 2467 2374
rect 2397 2375 2398 2482
rect 2466 2375 2467 2482
rect 2448 2347 2449 2378
rect 2469 2377 2470 2482
rect 2350 2347 2351 2380
rect 2448 2379 2449 2482
rect 2457 2347 2458 2380
rect 2490 2379 2491 2482
rect 2472 2347 2473 2382
rect 2478 2381 2479 2482
rect 2472 2383 2473 2482
rect 2505 2347 2506 2384
rect 2475 2347 2476 2386
rect 2484 2385 2485 2482
rect 2502 2347 2503 2386
rect 2511 2385 2512 2482
rect 2343 2347 2344 2388
rect 2502 2387 2503 2482
rect 2342 2389 2343 2482
rect 2400 2347 2401 2390
rect 2514 2347 2515 2390
rect 2550 2389 2551 2482
rect 2517 2347 2518 2392
rect 2580 2391 2581 2482
rect 2487 2347 2488 2394
rect 2517 2393 2518 2482
rect 2523 2347 2524 2394
rect 2553 2393 2554 2482
rect 2523 2395 2524 2482
rect 2562 2347 2563 2396
rect 2538 2347 2539 2398
rect 2541 2397 2542 2482
rect 2496 2347 2497 2400
rect 2538 2399 2539 2482
rect 2556 2347 2557 2400
rect 2586 2399 2587 2482
rect 2547 2347 2548 2402
rect 2556 2401 2557 2482
rect 2336 2347 2337 2404
rect 2547 2403 2548 2482
rect 2336 2405 2337 2482
rect 2785 2405 2786 2482
rect 2559 2347 2560 2408
rect 2583 2407 2584 2482
rect 2592 2347 2593 2408
rect 2626 2347 2627 2408
rect 2595 2347 2596 2410
rect 2625 2409 2626 2482
rect 2577 2347 2578 2412
rect 2595 2411 2596 2482
rect 2598 2347 2599 2412
rect 2622 2411 2623 2482
rect 2571 2347 2572 2414
rect 2598 2413 2599 2482
rect 2535 2347 2536 2416
rect 2571 2415 2572 2482
rect 2493 2347 2494 2418
rect 2535 2417 2536 2482
rect 2460 2347 2461 2420
rect 2493 2419 2494 2482
rect 2601 2347 2602 2420
rect 2616 2419 2617 2482
rect 2565 2347 2566 2422
rect 2601 2421 2602 2482
rect 2529 2347 2530 2424
rect 2565 2423 2566 2482
rect 2499 2347 2500 2426
rect 2529 2425 2530 2482
rect 2329 2427 2330 2482
rect 2499 2427 2500 2482
rect 2604 2347 2605 2428
rect 2634 2427 2635 2482
rect 2568 2347 2569 2430
rect 2604 2429 2605 2482
rect 2532 2347 2533 2432
rect 2568 2431 2569 2482
rect 2319 2433 2320 2482
rect 2532 2433 2533 2482
rect 2619 2433 2620 2482
rect 2747 2347 2748 2434
rect 2629 2347 2630 2436
rect 2658 2435 2659 2482
rect 2638 2347 2639 2438
rect 2667 2437 2668 2482
rect 2640 2439 2641 2482
rect 2641 2347 2642 2440
rect 2670 2439 2671 2482
rect 2767 2439 2768 2482
rect 2676 2441 2677 2482
rect 2739 2441 2740 2482
rect 2683 2347 2684 2444
rect 2717 2347 2718 2444
rect 2701 2347 2702 2446
rect 2718 2445 2719 2482
rect 2680 2347 2681 2448
rect 2700 2447 2701 2482
rect 2644 2347 2645 2450
rect 2679 2449 2680 2482
rect 2712 2449 2713 2482
rect 2732 2347 2733 2450
rect 2698 2347 2699 2452
rect 2733 2451 2734 2482
rect 2697 2453 2698 2482
rect 2723 2347 2724 2454
rect 2720 2347 2721 2456
rect 2769 2347 2770 2456
rect 2704 2347 2705 2458
rect 2721 2457 2722 2482
rect 2632 2347 2633 2460
rect 2703 2459 2704 2482
rect 2729 2347 2730 2460
rect 2788 2459 2789 2482
rect 2730 2461 2731 2482
rect 2816 2347 2817 2462
rect 2744 2347 2745 2464
rect 2812 2463 2813 2482
rect 2753 2347 2754 2466
rect 2773 2465 2774 2482
rect 2726 2347 2727 2468
rect 2752 2467 2753 2482
rect 2756 2347 2757 2468
rect 2776 2467 2777 2482
rect 2755 2469 2756 2482
rect 2762 2347 2763 2470
rect 2759 2347 2760 2472
rect 2791 2471 2792 2482
rect 2735 2347 2736 2474
rect 2758 2473 2759 2482
rect 2736 2475 2737 2482
rect 2849 2475 2850 2482
rect 2770 2477 2771 2482
rect 2779 2477 2780 2482
rect 2807 2347 2808 2478
rect 2836 2477 2837 2482
rect 2810 2347 2811 2480
rect 2839 2479 2840 2482
rect 2287 2486 2288 2489
rect 2339 2486 2340 2489
rect 2287 2490 2288 2601
rect 2294 2490 2295 2601
rect 2297 2490 2298 2601
rect 2301 2490 2302 2601
rect 2305 2486 2306 2491
rect 2504 2490 2505 2601
rect 2322 2486 2323 2493
rect 2359 2492 2360 2601
rect 2326 2486 2327 2495
rect 2493 2486 2494 2495
rect 2312 2486 2313 2497
rect 2492 2496 2493 2601
rect 2327 2498 2328 2601
rect 2532 2486 2533 2499
rect 2330 2500 2331 2601
rect 2348 2486 2349 2501
rect 2334 2502 2335 2601
rect 2529 2486 2530 2503
rect 2345 2486 2346 2505
rect 2436 2486 2437 2505
rect 2353 2506 2354 2601
rect 2365 2506 2366 2601
rect 2406 2486 2407 2507
rect 2414 2506 2415 2601
rect 2418 2486 2419 2507
rect 2426 2506 2427 2601
rect 2430 2486 2431 2507
rect 2450 2506 2451 2601
rect 2432 2508 2433 2601
rect 2448 2486 2449 2509
rect 2475 2486 2476 2509
rect 2604 2486 2605 2509
rect 2478 2486 2479 2511
rect 2507 2510 2508 2601
rect 2484 2486 2485 2513
rect 2519 2512 2520 2601
rect 2499 2486 2500 2515
rect 2513 2514 2514 2601
rect 2517 2486 2518 2515
rect 2543 2514 2544 2601
rect 2502 2486 2503 2517
rect 2516 2516 2517 2601
rect 2490 2486 2491 2519
rect 2501 2518 2502 2601
rect 2531 2518 2532 2601
rect 2535 2486 2536 2519
rect 2534 2520 2535 2601
rect 2538 2486 2539 2521
rect 2511 2486 2512 2523
rect 2537 2522 2538 2601
rect 2481 2486 2482 2525
rect 2510 2524 2511 2601
rect 2553 2486 2554 2525
rect 2561 2524 2562 2601
rect 2565 2486 2566 2525
rect 2573 2524 2574 2601
rect 2568 2486 2569 2527
rect 2576 2526 2577 2601
rect 2547 2486 2548 2529
rect 2567 2528 2568 2601
rect 2320 2530 2321 2601
rect 2546 2530 2547 2601
rect 2571 2486 2572 2531
rect 2591 2530 2592 2601
rect 2550 2486 2551 2533
rect 2570 2532 2571 2601
rect 2541 2486 2542 2535
rect 2549 2534 2550 2601
rect 2586 2486 2587 2535
rect 2609 2534 2610 2601
rect 2454 2486 2455 2537
rect 2585 2536 2586 2601
rect 2598 2486 2599 2537
rect 2636 2536 2637 2601
rect 2384 2538 2385 2601
rect 2597 2538 2598 2601
rect 2601 2486 2602 2539
rect 2627 2538 2628 2601
rect 2556 2486 2557 2541
rect 2600 2540 2601 2601
rect 2486 2542 2487 2601
rect 2555 2542 2556 2601
rect 2612 2542 2613 2601
rect 2631 2486 2632 2543
rect 2472 2486 2473 2545
rect 2630 2544 2631 2601
rect 2469 2486 2470 2547
rect 2471 2546 2472 2601
rect 2466 2486 2467 2549
rect 2468 2548 2469 2601
rect 2619 2486 2620 2549
rect 2645 2548 2646 2601
rect 2583 2486 2584 2551
rect 2618 2550 2619 2601
rect 2625 2486 2626 2551
rect 2651 2550 2652 2601
rect 2634 2486 2635 2553
rect 2682 2552 2683 2601
rect 2595 2486 2596 2555
rect 2633 2554 2634 2601
rect 2342 2486 2343 2557
rect 2594 2556 2595 2601
rect 2658 2486 2659 2557
rect 2706 2486 2707 2557
rect 2622 2486 2623 2559
rect 2657 2558 2658 2601
rect 2670 2486 2671 2559
rect 2673 2486 2674 2559
rect 2654 2560 2655 2601
rect 2669 2560 2670 2601
rect 2676 2560 2677 2601
rect 2773 2486 2774 2561
rect 2703 2486 2704 2563
rect 2706 2562 2707 2601
rect 2700 2486 2701 2565
rect 2703 2564 2704 2601
rect 2712 2486 2713 2565
rect 2810 2564 2811 2601
rect 2715 2566 2716 2601
rect 2776 2486 2777 2567
rect 2718 2486 2719 2569
rect 2769 2568 2770 2601
rect 2679 2486 2680 2571
rect 2718 2570 2719 2601
rect 2667 2486 2668 2573
rect 2679 2572 2680 2601
rect 2721 2486 2722 2573
rect 2724 2572 2725 2601
rect 2697 2486 2698 2575
rect 2721 2574 2722 2601
rect 2697 2576 2698 2601
rect 2842 2486 2843 2577
rect 2730 2486 2731 2579
rect 2760 2578 2761 2601
rect 2733 2486 2734 2581
rect 2763 2580 2764 2601
rect 2640 2486 2641 2583
rect 2733 2582 2734 2601
rect 2616 2486 2617 2585
rect 2639 2584 2640 2601
rect 2580 2486 2581 2587
rect 2615 2586 2616 2601
rect 2736 2486 2737 2587
rect 2845 2486 2846 2587
rect 2755 2486 2756 2589
rect 2791 2588 2792 2601
rect 2758 2486 2759 2591
rect 2836 2486 2837 2591
rect 2766 2592 2767 2601
rect 2819 2486 2820 2593
rect 2788 2486 2789 2595
rect 2808 2486 2809 2595
rect 2785 2486 2786 2597
rect 2807 2596 2808 2601
rect 2752 2486 2753 2599
rect 2785 2598 2786 2601
rect 2788 2598 2789 2601
rect 2804 2598 2805 2601
rect 2839 2486 2840 2599
rect 2861 2598 2862 2601
rect 2287 2605 2288 2608
rect 2325 2607 2326 2746
rect 2301 2605 2302 2610
rect 2504 2605 2505 2610
rect 2313 2605 2314 2612
rect 2359 2605 2360 2612
rect 2320 2605 2321 2614
rect 2346 2613 2347 2746
rect 2327 2605 2328 2616
rect 2513 2605 2514 2616
rect 2328 2617 2329 2746
rect 2785 2605 2786 2618
rect 2334 2605 2335 2620
rect 2482 2619 2483 2746
rect 2337 2605 2338 2622
rect 2567 2605 2568 2622
rect 2349 2605 2350 2624
rect 2353 2605 2354 2624
rect 2352 2625 2353 2746
rect 2546 2605 2547 2626
rect 2358 2627 2359 2746
rect 2513 2627 2514 2746
rect 2361 2629 2362 2746
rect 2492 2605 2493 2630
rect 2365 2631 2366 2746
rect 2534 2605 2535 2632
rect 2375 2633 2376 2746
rect 2379 2633 2380 2746
rect 2387 2605 2388 2634
rect 2585 2605 2586 2634
rect 2414 2605 2415 2636
rect 2416 2635 2417 2746
rect 2432 2605 2433 2636
rect 2434 2635 2435 2746
rect 2438 2605 2439 2636
rect 2679 2605 2680 2636
rect 2446 2637 2447 2746
rect 2450 2605 2451 2638
rect 2449 2639 2450 2746
rect 2516 2605 2517 2640
rect 2452 2641 2453 2746
rect 2564 2641 2565 2746
rect 2458 2643 2459 2746
rect 2570 2605 2571 2644
rect 2467 2645 2468 2746
rect 2468 2605 2469 2646
rect 2471 2605 2472 2646
rect 2567 2645 2568 2746
rect 2479 2647 2480 2746
rect 2501 2605 2502 2648
rect 2486 2605 2487 2650
rect 2603 2649 2604 2746
rect 2488 2651 2489 2746
rect 2555 2605 2556 2652
rect 2498 2653 2499 2746
rect 2507 2605 2508 2654
rect 2501 2655 2502 2746
rect 2510 2605 2511 2656
rect 2504 2657 2505 2746
rect 2537 2605 2538 2658
rect 2510 2659 2511 2746
rect 2543 2605 2544 2660
rect 2516 2661 2517 2746
rect 2519 2605 2520 2662
rect 2522 2661 2523 2746
rect 2531 2605 2532 2662
rect 2525 2605 2526 2664
rect 2633 2605 2634 2664
rect 2426 2605 2427 2666
rect 2525 2665 2526 2746
rect 2537 2665 2538 2746
rect 2630 2605 2631 2666
rect 2540 2667 2541 2746
rect 2561 2605 2562 2668
rect 2546 2669 2547 2746
rect 2573 2605 2574 2670
rect 2552 2671 2553 2746
rect 2591 2605 2592 2672
rect 2549 2605 2550 2674
rect 2591 2673 2592 2746
rect 2549 2675 2550 2746
rect 2576 2605 2577 2676
rect 2555 2677 2556 2746
rect 2594 2605 2595 2678
rect 2558 2679 2559 2746
rect 2597 2605 2598 2680
rect 2561 2681 2562 2746
rect 2600 2605 2601 2682
rect 2582 2683 2583 2746
rect 2609 2605 2610 2684
rect 2585 2685 2586 2746
rect 2612 2605 2613 2686
rect 2588 2687 2589 2746
rect 2627 2605 2628 2688
rect 2594 2689 2595 2746
rect 2618 2605 2619 2690
rect 2600 2691 2601 2746
rect 2615 2605 2616 2692
rect 2606 2693 2607 2746
rect 2645 2605 2646 2694
rect 2612 2695 2613 2746
rect 2651 2605 2652 2696
rect 2615 2697 2616 2746
rect 2636 2605 2637 2698
rect 2618 2699 2619 2746
rect 2639 2605 2640 2700
rect 2624 2701 2625 2746
rect 2682 2605 2683 2702
rect 2633 2703 2634 2746
rect 2657 2605 2658 2704
rect 2636 2705 2637 2746
rect 2654 2605 2655 2706
rect 2665 2705 2666 2746
rect 2788 2605 2789 2706
rect 2677 2707 2678 2746
rect 2721 2605 2722 2708
rect 2680 2709 2681 2746
rect 2703 2605 2704 2710
rect 2683 2711 2684 2746
rect 2706 2605 2707 2712
rect 2694 2605 2695 2714
rect 2858 2605 2859 2714
rect 2697 2605 2698 2716
rect 2797 2605 2798 2716
rect 2698 2717 2699 2746
rect 2760 2605 2761 2718
rect 2701 2719 2702 2746
rect 2766 2605 2767 2720
rect 2704 2721 2705 2746
rect 2724 2605 2725 2722
rect 2707 2723 2708 2746
rect 2724 2723 2725 2746
rect 2715 2605 2716 2726
rect 2874 2605 2875 2726
rect 2718 2605 2719 2728
rect 2779 2727 2780 2746
rect 2730 2729 2731 2746
rect 2791 2605 2792 2730
rect 2733 2605 2734 2732
rect 2769 2605 2770 2732
rect 2733 2733 2734 2746
rect 2827 2605 2828 2734
rect 2736 2735 2737 2746
rect 2837 2605 2838 2736
rect 2742 2737 2743 2746
rect 2807 2605 2808 2738
rect 2745 2739 2746 2746
rect 2810 2605 2811 2740
rect 2763 2605 2764 2742
rect 2867 2605 2868 2742
rect 2782 2743 2783 2746
rect 2861 2605 2862 2744
rect 2296 2752 2297 2871
rect 2340 2752 2341 2871
rect 2303 2754 2304 2871
rect 2308 2750 2309 2755
rect 2312 2750 2313 2755
rect 2319 2750 2320 2755
rect 2306 2756 2307 2871
rect 2313 2756 2314 2871
rect 2319 2756 2320 2871
rect 2325 2750 2326 2757
rect 2322 2750 2323 2759
rect 2328 2750 2329 2759
rect 2328 2760 2329 2871
rect 2513 2750 2514 2761
rect 2343 2762 2344 2871
rect 2346 2750 2347 2763
rect 2349 2762 2350 2871
rect 2352 2750 2353 2763
rect 2369 2762 2370 2871
rect 2549 2750 2550 2763
rect 2375 2750 2376 2765
rect 2555 2750 2556 2765
rect 2386 2750 2387 2767
rect 2416 2750 2417 2767
rect 2415 2768 2416 2871
rect 2434 2750 2435 2769
rect 2433 2770 2434 2871
rect 2446 2750 2447 2771
rect 2436 2772 2437 2871
rect 2449 2750 2450 2773
rect 2442 2774 2443 2871
rect 2529 2774 2530 2871
rect 2458 2750 2459 2777
rect 2532 2776 2533 2871
rect 2457 2778 2458 2871
rect 2467 2750 2468 2779
rect 2460 2780 2461 2871
rect 2567 2750 2568 2781
rect 2463 2782 2464 2871
rect 2479 2750 2480 2783
rect 2466 2784 2467 2871
rect 2482 2750 2483 2785
rect 2481 2786 2482 2871
rect 2498 2750 2499 2787
rect 2484 2788 2485 2871
rect 2501 2750 2502 2789
rect 2362 2790 2363 2871
rect 2502 2790 2503 2871
rect 2493 2792 2494 2871
rect 2504 2750 2505 2793
rect 2495 2750 2496 2795
rect 2603 2750 2604 2795
rect 2499 2796 2500 2871
rect 2510 2750 2511 2797
rect 2505 2798 2506 2871
rect 2522 2750 2523 2799
rect 2508 2800 2509 2871
rect 2525 2750 2526 2801
rect 2516 2750 2517 2803
rect 2538 2802 2539 2871
rect 2517 2804 2518 2871
rect 2540 2750 2541 2805
rect 2382 2750 2383 2807
rect 2541 2806 2542 2871
rect 2523 2808 2524 2871
rect 2585 2750 2586 2809
rect 2550 2810 2551 2871
rect 2558 2750 2559 2811
rect 2564 2750 2565 2811
rect 2650 2810 2651 2871
rect 2473 2750 2474 2813
rect 2565 2812 2566 2871
rect 2574 2812 2575 2871
rect 2600 2750 2601 2813
rect 2577 2814 2578 2871
rect 2588 2750 2589 2815
rect 2534 2750 2535 2817
rect 2589 2816 2590 2871
rect 2535 2818 2536 2871
rect 2546 2750 2547 2819
rect 2547 2820 2548 2871
rect 2552 2750 2553 2821
rect 2553 2822 2554 2871
rect 2561 2750 2562 2823
rect 2562 2824 2563 2871
rect 2582 2750 2583 2825
rect 2580 2826 2581 2871
rect 2591 2750 2592 2827
rect 2594 2750 2595 2827
rect 2642 2750 2643 2827
rect 2595 2828 2596 2871
rect 2606 2750 2607 2829
rect 2592 2830 2593 2871
rect 2607 2830 2608 2871
rect 2601 2832 2602 2871
rect 2612 2750 2613 2833
rect 2604 2834 2605 2871
rect 2615 2750 2616 2835
rect 2610 2836 2611 2871
rect 2624 2750 2625 2837
rect 2613 2838 2614 2871
rect 2618 2750 2619 2839
rect 2625 2838 2626 2871
rect 2633 2750 2634 2839
rect 2628 2840 2629 2871
rect 2636 2750 2637 2841
rect 2637 2842 2638 2871
rect 2683 2750 2684 2843
rect 2643 2844 2644 2871
rect 2646 2750 2647 2845
rect 2668 2750 2669 2845
rect 2727 2750 2728 2845
rect 2668 2846 2669 2871
rect 2677 2750 2678 2847
rect 2686 2846 2687 2871
rect 2698 2750 2699 2847
rect 2689 2848 2690 2871
rect 2704 2750 2705 2849
rect 2661 2750 2662 2851
rect 2704 2850 2705 2871
rect 2701 2750 2702 2853
rect 2717 2750 2718 2853
rect 2701 2854 2702 2871
rect 2736 2750 2737 2855
rect 2707 2750 2708 2857
rect 2710 2856 2711 2871
rect 2680 2750 2681 2859
rect 2707 2858 2708 2871
rect 2713 2858 2714 2871
rect 2720 2858 2721 2871
rect 2730 2750 2731 2859
rect 2739 2858 2740 2871
rect 2733 2858 2734 2871
rect 2733 2750 2734 2859
rect 2736 2860 2737 2871
rect 2758 2750 2759 2861
rect 2742 2750 2743 2863
rect 2751 2862 2752 2871
rect 2727 2864 2728 2871
rect 2742 2864 2743 2871
rect 2745 2750 2746 2865
rect 2754 2864 2755 2871
rect 2723 2866 2724 2871
rect 2745 2866 2746 2871
rect 2782 2750 2783 2867
rect 2791 2866 2792 2871
rect 2683 2868 2684 2871
rect 2781 2868 2782 2871
rect 2300 2875 2301 2878
rect 2340 2875 2341 2878
rect 2296 2875 2297 2880
rect 2300 2879 2301 2972
rect 2309 2875 2310 2880
rect 2399 2879 2400 2972
rect 2313 2875 2314 2882
rect 2387 2881 2388 2972
rect 2319 2875 2320 2884
rect 2383 2875 2384 2884
rect 2296 2885 2297 2972
rect 2384 2885 2385 2972
rect 2321 2887 2322 2972
rect 2499 2875 2500 2888
rect 2324 2889 2325 2972
rect 2493 2875 2494 2890
rect 2328 2875 2329 2892
rect 2333 2891 2334 2972
rect 2343 2875 2344 2892
rect 2345 2891 2346 2972
rect 2349 2875 2350 2892
rect 2351 2891 2352 2972
rect 2358 2875 2359 2892
rect 2436 2875 2437 2892
rect 2357 2893 2358 2972
rect 2514 2893 2515 2972
rect 2364 2895 2365 2972
rect 2365 2875 2366 2896
rect 2376 2875 2377 2896
rect 2601 2875 2602 2896
rect 2390 2897 2391 2972
rect 2502 2875 2503 2898
rect 2367 2899 2368 2972
rect 2502 2899 2503 2972
rect 2405 2901 2406 2972
rect 2559 2901 2560 2972
rect 2433 2901 2434 2972
rect 2433 2875 2434 2902
rect 2439 2875 2440 2904
rect 2565 2875 2566 2904
rect 2415 2875 2416 2906
rect 2439 2905 2440 2972
rect 2457 2875 2458 2906
rect 2475 2905 2476 2972
rect 2460 2875 2461 2908
rect 2469 2907 2470 2972
rect 2463 2907 2464 2972
rect 2463 2875 2464 2908
rect 2466 2907 2467 2972
rect 2466 2875 2467 2908
rect 2478 2907 2479 2972
rect 2481 2875 2482 2908
rect 2481 2909 2482 2972
rect 2484 2875 2485 2910
rect 2490 2909 2491 2972
rect 2505 2875 2506 2910
rect 2493 2911 2494 2972
rect 2508 2875 2509 2912
rect 2508 2913 2509 2972
rect 2517 2875 2518 2914
rect 2355 2875 2356 2916
rect 2517 2915 2518 2972
rect 2523 2875 2524 2916
rect 2568 2915 2569 2972
rect 2526 2917 2527 2972
rect 2535 2875 2536 2918
rect 2532 2875 2533 2920
rect 2535 2919 2536 2972
rect 2529 2875 2530 2922
rect 2532 2921 2533 2972
rect 2544 2921 2545 2972
rect 2550 2875 2551 2922
rect 2547 2875 2548 2924
rect 2550 2923 2551 2972
rect 2547 2925 2548 2972
rect 2553 2875 2554 2926
rect 2562 2875 2563 2926
rect 2565 2925 2566 2972
rect 2538 2875 2539 2928
rect 2562 2927 2563 2972
rect 2538 2929 2539 2972
rect 2541 2875 2542 2930
rect 2580 2875 2581 2930
rect 2583 2929 2584 2972
rect 2577 2875 2578 2932
rect 2580 2931 2581 2972
rect 2574 2875 2575 2934
rect 2577 2933 2578 2972
rect 2592 2933 2593 2972
rect 2791 2875 2792 2934
rect 2595 2875 2596 2936
rect 2622 2935 2623 2972
rect 2607 2875 2608 2938
rect 2616 2937 2617 2972
rect 2610 2937 2611 2972
rect 2610 2875 2611 2938
rect 2613 2875 2614 2940
rect 2619 2939 2620 2972
rect 2604 2875 2605 2942
rect 2613 2941 2614 2972
rect 2631 2941 2632 2972
rect 2646 2875 2647 2942
rect 2634 2943 2635 2972
rect 2713 2875 2714 2944
rect 2637 2875 2638 2946
rect 2646 2945 2647 2972
rect 2637 2947 2638 2972
rect 2698 2875 2699 2948
rect 2668 2875 2669 2950
rect 2671 2949 2672 2972
rect 2683 2875 2684 2950
rect 2762 2949 2763 2972
rect 2686 2949 2687 2972
rect 2686 2875 2687 2950
rect 2689 2875 2690 2952
rect 2695 2951 2696 2972
rect 2689 2953 2690 2972
rect 2769 2953 2770 2972
rect 2692 2955 2693 2972
rect 2765 2955 2766 2972
rect 2704 2955 2705 2972
rect 2704 2875 2705 2956
rect 2707 2955 2708 2972
rect 2707 2875 2708 2956
rect 2710 2875 2711 2958
rect 2720 2957 2721 2972
rect 2658 2959 2659 2972
rect 2710 2959 2711 2972
rect 2730 2959 2731 2972
rect 2733 2875 2734 2960
rect 2733 2961 2734 2972
rect 2736 2875 2737 2962
rect 2628 2875 2629 2964
rect 2736 2963 2737 2972
rect 2625 2875 2626 2966
rect 2628 2965 2629 2972
rect 2739 2875 2740 2966
rect 2760 2875 2761 2966
rect 2742 2875 2743 2968
rect 2748 2875 2749 2968
rect 2751 2875 2752 2968
rect 2756 2967 2757 2972
rect 2754 2875 2755 2970
rect 2759 2969 2760 2972
rect 2296 2976 2297 2979
rect 2300 2976 2301 2979
rect 2299 2980 2300 3101
rect 2466 2976 2467 2981
rect 2307 2976 2308 2983
rect 2384 2976 2385 2983
rect 2314 2976 2315 2985
rect 2345 2976 2346 2985
rect 2320 2986 2321 3101
rect 2333 2976 2334 2987
rect 2329 2988 2330 3101
rect 2517 2976 2518 2989
rect 2349 2990 2350 3101
rect 2387 2976 2388 2991
rect 2351 2976 2352 2993
rect 2409 2976 2410 2993
rect 2352 2994 2353 3101
rect 2390 2976 2391 2995
rect 2355 2996 2356 3101
rect 2550 2976 2551 2997
rect 2357 2976 2358 2999
rect 2371 2976 2372 2999
rect 2358 3000 2359 3101
rect 2451 3000 2452 3101
rect 2360 2976 2361 3003
rect 2399 2976 2400 3003
rect 2381 2976 2382 3005
rect 2514 2976 2515 3005
rect 2381 3006 2382 3101
rect 2433 2976 2434 3007
rect 2384 3008 2385 3101
rect 2439 2976 2440 3009
rect 2396 3010 2397 3101
rect 2538 2976 2539 3011
rect 2409 3012 2410 3101
rect 2469 2976 2470 3013
rect 2412 3014 2413 3101
rect 2547 2976 2548 3015
rect 2424 3016 2425 3101
rect 2478 2976 2479 3017
rect 2365 3018 2366 3101
rect 2478 3018 2479 3101
rect 2430 3020 2431 3101
rect 2490 2976 2491 3021
rect 2433 3022 2434 3101
rect 2472 3022 2473 3101
rect 2445 3024 2446 3101
rect 2502 2976 2503 3025
rect 2402 2976 2403 3027
rect 2502 3026 2503 3101
rect 2403 3028 2404 3101
rect 2493 2976 2494 3029
rect 2460 3030 2461 3101
rect 2526 2976 2527 3031
rect 2481 3030 2482 3101
rect 2481 2976 2482 3031
rect 2484 3032 2485 3101
rect 2532 2976 2533 3033
rect 2487 3034 2488 3101
rect 2535 2976 2536 3035
rect 2490 3036 2491 3101
rect 2544 2976 2545 3037
rect 2493 3038 2494 3101
rect 2508 2976 2509 3039
rect 2508 3040 2509 3101
rect 2559 2976 2560 3041
rect 2511 3042 2512 3101
rect 2562 2976 2563 3043
rect 2514 3044 2515 3101
rect 2565 2976 2566 3045
rect 2517 3046 2518 3101
rect 2568 2976 2569 3047
rect 2526 3048 2527 3101
rect 2577 2976 2578 3049
rect 2529 3050 2530 3101
rect 2580 2976 2581 3051
rect 2532 3052 2533 3101
rect 2583 2976 2584 3053
rect 2541 3054 2542 3101
rect 2613 2976 2614 3055
rect 2544 3056 2545 3101
rect 2616 2976 2617 3057
rect 2559 3058 2560 3101
rect 2610 2976 2611 3059
rect 2562 3060 2563 3101
rect 2619 2976 2620 3061
rect 2565 3062 2566 3101
rect 2622 2976 2623 3063
rect 2568 3064 2569 3101
rect 2631 2976 2632 3065
rect 2577 3066 2578 3101
rect 2637 2976 2638 3067
rect 2586 3068 2587 3101
rect 2646 2976 2647 3069
rect 2610 3070 2611 3101
rect 2671 2976 2672 3071
rect 2613 3072 2614 3101
rect 2695 2976 2696 3073
rect 2622 3074 2623 3101
rect 2689 2976 2690 3075
rect 2625 3076 2626 3101
rect 2686 2976 2687 3077
rect 2628 3078 2629 3101
rect 2692 2976 2693 3079
rect 2631 3080 2632 3101
rect 2650 3080 2651 3101
rect 2634 2976 2635 3083
rect 2643 2976 2644 3083
rect 2463 2976 2464 3085
rect 2634 3084 2635 3101
rect 2637 3084 2638 3101
rect 2704 2976 2705 3085
rect 2640 3086 2641 3101
rect 2707 2976 2708 3087
rect 2661 2976 2662 3089
rect 2665 2976 2666 3089
rect 2663 3090 2664 3101
rect 2730 2976 2731 3091
rect 2666 3092 2667 3101
rect 2733 2976 2734 3093
rect 2689 3094 2690 3101
rect 2756 2976 2757 3095
rect 2692 3096 2693 3101
rect 2759 2976 2760 3097
rect 2698 3098 2699 3101
rect 2772 2976 2773 3099
rect 2299 3105 2300 3108
rect 2312 3107 2313 3190
rect 2306 3109 2307 3190
rect 2315 3109 2316 3190
rect 2317 3105 2318 3110
rect 2352 3105 2353 3110
rect 2329 3105 2330 3112
rect 2349 3105 2350 3112
rect 2332 3113 2333 3190
rect 2440 3113 2441 3190
rect 2336 3105 2337 3116
rect 2396 3115 2397 3190
rect 2343 3105 2344 3118
rect 2511 3105 2512 3118
rect 2356 3119 2357 3190
rect 2451 3105 2452 3120
rect 2362 3105 2363 3122
rect 2472 3105 2473 3122
rect 2372 3123 2373 3190
rect 2384 3105 2385 3124
rect 2381 3105 2382 3126
rect 2443 3125 2444 3190
rect 2406 3127 2407 3190
rect 2409 3105 2410 3128
rect 2419 3127 2420 3190
rect 2424 3105 2425 3128
rect 2425 3129 2426 3190
rect 2430 3105 2431 3130
rect 2434 3129 2435 3190
rect 2445 3105 2446 3130
rect 2470 3129 2471 3190
rect 2478 3105 2479 3130
rect 2473 3131 2474 3190
rect 2481 3105 2482 3132
rect 2476 3133 2477 3190
rect 2484 3105 2485 3134
rect 2479 3135 2480 3190
rect 2487 3105 2488 3136
rect 2482 3137 2483 3190
rect 2490 3105 2491 3138
rect 2485 3139 2486 3190
rect 2493 3105 2494 3140
rect 2494 3141 2495 3190
rect 2502 3105 2503 3142
rect 2460 3105 2461 3144
rect 2503 3143 2504 3190
rect 2500 3145 2501 3190
rect 2508 3105 2509 3146
rect 2506 3147 2507 3190
rect 2514 3105 2515 3148
rect 2509 3149 2510 3190
rect 2517 3105 2518 3150
rect 2512 3151 2513 3190
rect 2532 3105 2533 3152
rect 2518 3153 2519 3190
rect 2526 3105 2527 3154
rect 2521 3155 2522 3190
rect 2529 3105 2530 3156
rect 2544 3105 2545 3156
rect 2548 3155 2549 3190
rect 2541 3105 2542 3158
rect 2545 3157 2546 3190
rect 2557 3157 2558 3190
rect 2574 3105 2575 3158
rect 2559 3105 2560 3160
rect 2560 3159 2561 3190
rect 2565 3105 2566 3160
rect 2566 3159 2567 3190
rect 2568 3105 2569 3160
rect 2581 3159 2582 3190
rect 2562 3105 2563 3162
rect 2569 3161 2570 3190
rect 2523 3105 2524 3164
rect 2563 3163 2564 3190
rect 2466 3105 2467 3166
rect 2524 3165 2525 3190
rect 2577 3105 2578 3166
rect 2584 3165 2585 3190
rect 2610 3105 2611 3166
rect 2617 3165 2618 3190
rect 2613 3105 2614 3168
rect 2644 3167 2645 3190
rect 2614 3169 2615 3190
rect 2705 3105 2706 3170
rect 2620 3171 2621 3190
rect 2692 3105 2693 3172
rect 2622 3105 2623 3174
rect 2703 3173 2704 3190
rect 2637 3105 2638 3176
rect 2646 3105 2647 3176
rect 2638 3177 2639 3190
rect 2640 3105 2641 3178
rect 2586 3105 2587 3180
rect 2641 3179 2642 3190
rect 2587 3181 2588 3190
rect 2632 3181 2633 3190
rect 2663 3105 2664 3182
rect 2681 3181 2682 3190
rect 2666 3105 2667 3184
rect 2684 3183 2685 3190
rect 2689 3105 2690 3184
rect 2730 3183 2731 3190
rect 2628 3105 2629 3186
rect 2690 3185 2691 3190
rect 2625 3105 2626 3188
rect 2629 3187 2630 3190
rect 2700 3187 2701 3190
rect 2727 3187 2728 3190
rect 2299 3194 2300 3197
rect 2306 3194 2307 3197
rect 2302 3198 2303 3307
rect 2312 3194 2313 3199
rect 2312 3200 2313 3307
rect 2325 3194 2326 3201
rect 2306 3202 2307 3307
rect 2325 3202 2326 3307
rect 2315 3194 2316 3205
rect 2318 3194 2319 3205
rect 2315 3206 2316 3307
rect 2396 3194 2397 3207
rect 2322 3208 2323 3307
rect 2440 3194 2441 3209
rect 2332 3194 2333 3211
rect 2482 3194 2483 3211
rect 2335 3212 2336 3307
rect 2425 3194 2426 3213
rect 2339 3194 2340 3215
rect 2494 3194 2495 3215
rect 2356 3216 2357 3307
rect 2387 3194 2388 3217
rect 2359 3218 2360 3307
rect 2383 3218 2384 3307
rect 2368 3220 2369 3307
rect 2372 3194 2373 3221
rect 2380 3220 2381 3307
rect 2443 3194 2444 3221
rect 2404 3222 2405 3307
rect 2409 3194 2410 3223
rect 2417 3222 2418 3307
rect 2490 3222 2491 3307
rect 2419 3194 2420 3225
rect 2736 3194 2737 3225
rect 2433 3226 2434 3307
rect 2434 3194 2435 3227
rect 2439 3226 2440 3307
rect 2485 3194 2486 3227
rect 2448 3228 2449 3307
rect 2512 3194 2513 3229
rect 2460 3230 2461 3307
rect 2476 3194 2477 3231
rect 2463 3232 2464 3307
rect 2479 3194 2480 3233
rect 2466 3234 2467 3307
rect 2470 3194 2471 3235
rect 2469 3236 2470 3307
rect 2473 3194 2474 3237
rect 2472 3238 2473 3307
rect 2506 3194 2507 3239
rect 2484 3240 2485 3307
rect 2500 3194 2501 3241
rect 2487 3242 2488 3307
rect 2503 3194 2504 3243
rect 2493 3244 2494 3307
rect 2509 3194 2510 3245
rect 2496 3246 2497 3307
rect 2518 3194 2519 3247
rect 2505 3248 2506 3307
rect 2521 3194 2522 3249
rect 2424 3250 2425 3307
rect 2520 3250 2521 3307
rect 2508 3252 2509 3307
rect 2524 3194 2525 3253
rect 2511 3254 2512 3307
rect 2548 3194 2549 3255
rect 2514 3256 2515 3307
rect 2545 3194 2546 3257
rect 2523 3258 2524 3307
rect 2566 3194 2567 3259
rect 2526 3260 2527 3307
rect 2581 3194 2582 3261
rect 2529 3262 2530 3307
rect 2560 3194 2561 3263
rect 2539 3264 2540 3307
rect 2557 3194 2558 3265
rect 2542 3266 2543 3307
rect 2654 3194 2655 3267
rect 2558 3268 2559 3307
rect 2638 3194 2639 3269
rect 2561 3270 2562 3307
rect 2641 3194 2642 3271
rect 2563 3194 2564 3273
rect 2572 3194 2573 3273
rect 2564 3274 2565 3307
rect 2644 3194 2645 3275
rect 2569 3194 2570 3277
rect 2608 3194 2609 3277
rect 2573 3278 2574 3307
rect 2587 3194 2588 3279
rect 2584 3194 2585 3281
rect 2664 3194 2665 3281
rect 2600 3282 2601 3307
rect 2620 3194 2621 3283
rect 2609 3284 2610 3307
rect 2678 3194 2679 3285
rect 2612 3286 2613 3307
rect 2617 3194 2618 3287
rect 2614 3194 2615 3289
rect 2671 3194 2672 3289
rect 2615 3290 2616 3307
rect 2635 3194 2636 3291
rect 2618 3292 2619 3307
rect 2624 3292 2625 3307
rect 2627 3292 2628 3307
rect 2681 3194 2682 3293
rect 2629 3194 2630 3295
rect 2697 3194 2698 3295
rect 2630 3296 2631 3307
rect 2684 3194 2685 3297
rect 2646 3298 2647 3307
rect 2690 3298 2691 3307
rect 2649 3300 2650 3307
rect 2703 3194 2704 3301
rect 2676 3302 2677 3307
rect 2700 3194 2701 3303
rect 2700 3304 2701 3307
rect 2707 3304 2708 3307
rect 2309 3311 2310 3314
rect 2315 3311 2316 3314
rect 2319 3311 2320 3314
rect 2496 3311 2497 3314
rect 2321 3315 2322 3390
rect 2325 3311 2326 3316
rect 2335 3315 2336 3390
rect 2484 3311 2485 3316
rect 2368 3311 2369 3318
rect 2377 3317 2378 3390
rect 2380 3311 2381 3318
rect 2389 3317 2390 3390
rect 2383 3311 2384 3320
rect 2392 3319 2393 3390
rect 2398 3311 2399 3320
rect 2410 3311 2411 3320
rect 2402 3321 2403 3390
rect 2649 3311 2650 3322
rect 2407 3311 2408 3324
rect 2424 3311 2425 3324
rect 2404 3311 2405 3326
rect 2408 3325 2409 3390
rect 2414 3325 2415 3390
rect 2472 3311 2473 3326
rect 2417 3311 2418 3328
rect 2505 3311 2506 3328
rect 2424 3329 2425 3390
rect 2433 3311 2434 3330
rect 2436 3329 2437 3390
rect 2460 3311 2461 3330
rect 2451 3331 2452 3390
rect 2466 3311 2467 3332
rect 2454 3333 2455 3390
rect 2469 3311 2470 3334
rect 2463 3311 2464 3336
rect 2716 3311 2717 3336
rect 2448 3311 2449 3338
rect 2463 3337 2464 3390
rect 2439 3311 2440 3340
rect 2448 3339 2449 3390
rect 2290 3341 2291 3390
rect 2439 3341 2440 3390
rect 2466 3341 2467 3390
rect 2508 3311 2509 3342
rect 2475 3343 2476 3390
rect 2490 3311 2491 3344
rect 2478 3345 2479 3390
rect 2493 3311 2494 3346
rect 2487 3311 2488 3348
rect 2634 3347 2635 3390
rect 2493 3349 2494 3390
rect 2511 3311 2512 3350
rect 2487 3351 2488 3390
rect 2512 3351 2513 3390
rect 2496 3353 2497 3390
rect 2514 3311 2515 3354
rect 2499 3355 2500 3390
rect 2523 3311 2524 3356
rect 2515 3357 2516 3390
rect 2529 3311 2530 3358
rect 2517 3311 2518 3360
rect 2539 3311 2540 3360
rect 2518 3361 2519 3390
rect 2526 3311 2527 3362
rect 2538 3361 2539 3390
rect 2561 3311 2562 3362
rect 2544 3363 2545 3390
rect 2558 3311 2559 3364
rect 2547 3365 2548 3390
rect 2564 3311 2565 3366
rect 2559 3367 2560 3390
rect 2612 3311 2613 3368
rect 2568 3369 2569 3390
rect 2624 3311 2625 3370
rect 2571 3371 2572 3390
rect 2618 3311 2619 3372
rect 2573 3311 2574 3374
rect 2591 3311 2592 3374
rect 2553 3375 2554 3390
rect 2574 3375 2575 3390
rect 2584 3375 2585 3390
rect 2600 3311 2601 3376
rect 2587 3377 2588 3390
rect 2627 3311 2628 3378
rect 2609 3311 2610 3380
rect 2652 3311 2653 3380
rect 2615 3311 2616 3382
rect 2621 3311 2622 3382
rect 2630 3311 2631 3382
rect 2662 3311 2663 3382
rect 2637 3383 2638 3390
rect 2683 3311 2684 3384
rect 2646 3311 2647 3386
rect 2673 3311 2674 3386
rect 2655 3311 2656 3388
rect 2687 3311 2688 3388
rect 2696 3311 2697 3388
rect 2700 3311 2701 3388
rect 2311 3394 2312 3397
rect 2318 3394 2319 3397
rect 2320 3396 2321 3459
rect 2332 3394 2333 3397
rect 2328 3394 2329 3399
rect 2424 3394 2425 3399
rect 2331 3400 2332 3459
rect 2345 3400 2346 3459
rect 2335 3394 2336 3403
rect 2436 3394 2437 3403
rect 2334 3404 2335 3459
rect 2439 3394 2440 3405
rect 2371 3406 2372 3459
rect 2389 3394 2390 3407
rect 2374 3408 2375 3459
rect 2392 3394 2393 3409
rect 2377 3394 2378 3411
rect 2383 3410 2384 3459
rect 2392 3410 2393 3459
rect 2408 3394 2409 3411
rect 2398 3412 2399 3459
rect 2475 3394 2476 3413
rect 2402 3414 2403 3459
rect 2463 3394 2464 3415
rect 2408 3416 2409 3459
rect 2512 3394 2513 3417
rect 2411 3418 2412 3459
rect 2448 3394 2449 3419
rect 2414 3420 2415 3459
rect 2478 3394 2479 3421
rect 2418 3394 2419 3423
rect 2466 3394 2467 3423
rect 2420 3424 2421 3459
rect 2451 3394 2452 3425
rect 2430 3394 2431 3427
rect 2454 3394 2455 3427
rect 2436 3428 2437 3459
rect 2487 3394 2488 3429
rect 2442 3430 2443 3459
rect 2493 3394 2494 3431
rect 2445 3432 2446 3459
rect 2496 3394 2497 3433
rect 2495 3434 2496 3459
rect 2568 3394 2569 3435
rect 2499 3394 2500 3437
rect 2502 3394 2503 3437
rect 2498 3438 2499 3459
rect 2571 3394 2572 3439
rect 2501 3440 2502 3459
rect 2547 3394 2548 3441
rect 2504 3442 2505 3459
rect 2553 3394 2554 3443
rect 2507 3444 2508 3459
rect 2559 3394 2560 3445
rect 2515 3394 2516 3447
rect 2528 3446 2529 3459
rect 2522 3448 2523 3459
rect 2587 3394 2588 3449
rect 2525 3450 2526 3459
rect 2604 3394 2605 3451
rect 2538 3394 2539 3453
rect 2634 3394 2635 3453
rect 2541 3454 2542 3459
rect 2618 3394 2619 3455
rect 2571 3456 2572 3459
rect 2637 3394 2638 3457
rect 2287 3463 2288 3466
rect 2462 3463 2463 3466
rect 2324 3463 2325 3468
rect 2445 3463 2446 3468
rect 2356 3469 2357 3498
rect 2371 3463 2372 3470
rect 2359 3471 2360 3498
rect 2374 3463 2375 3472
rect 2379 3471 2380 3498
rect 2411 3463 2412 3472
rect 2383 3463 2384 3474
rect 2390 3473 2391 3498
rect 2392 3463 2393 3474
rect 2535 3463 2536 3474
rect 2403 3475 2404 3498
rect 2414 3463 2415 3476
rect 2406 3477 2407 3498
rect 2408 3463 2409 3478
rect 2415 3477 2416 3498
rect 2448 3463 2449 3478
rect 2421 3479 2422 3498
rect 2436 3463 2437 3480
rect 2424 3481 2425 3498
rect 2442 3463 2443 3482
rect 2474 3481 2475 3498
rect 2495 3463 2496 3482
rect 2477 3483 2478 3498
rect 2498 3463 2499 3484
rect 2486 3485 2487 3498
rect 2507 3463 2508 3486
rect 2501 3487 2502 3498
rect 2522 3463 2523 3488
rect 2504 3463 2505 3490
rect 2516 3463 2517 3490
rect 2504 3491 2505 3498
rect 2525 3463 2526 3492
rect 2520 3493 2521 3498
rect 2541 3463 2542 3494
rect 2523 3495 2524 3498
rect 2544 3463 2545 3496
rect 2550 3495 2551 3498
rect 2571 3463 2572 3496
rect 2577 3463 2578 3496
rect 2584 3463 2585 3496
rect 2323 3502 2324 3505
rect 2359 3502 2360 3505
rect 2356 3502 2357 3507
rect 2388 3506 2389 3519
rect 2391 3506 2392 3519
rect 2406 3502 2407 3507
rect 2393 3502 2394 3509
rect 2403 3502 2404 3509
rect 2406 3508 2407 3519
rect 2427 3502 2428 3509
rect 2409 3510 2410 3519
rect 2415 3502 2416 3511
rect 2418 3510 2419 3519
rect 2424 3502 2425 3511
rect 2441 3502 2442 3511
rect 2520 3502 2521 3511
rect 2468 3512 2469 3519
rect 2474 3502 2475 3513
rect 2471 3514 2472 3519
rect 2477 3502 2478 3515
rect 2480 3514 2481 3519
rect 2486 3502 2487 3515
rect 2495 3514 2496 3519
rect 2523 3502 2524 3515
rect 2498 3516 2499 3519
rect 2501 3502 2502 3517
rect 2504 3502 2505 3517
rect 2518 3516 2519 3519
rect 2550 3502 2551 3517
rect 2556 3502 2557 3517
rect 2563 3502 2564 3517
rect 2570 3502 2571 3517
rect 2383 3525 2384 3542
rect 2391 3523 2392 3526
rect 2388 3523 2389 3528
rect 2480 3523 2481 3528
rect 2392 3529 2393 3542
rect 2418 3523 2419 3530
rect 2394 3523 2395 3532
rect 2406 3523 2407 3532
rect 2397 3523 2398 3534
rect 2409 3523 2410 3534
rect 2431 3533 2432 3542
rect 2468 3523 2469 3534
rect 2437 3535 2438 3542
rect 2471 3523 2472 3536
rect 2454 3537 2455 3542
rect 2498 3523 2499 3538
rect 2495 3523 2496 3540
rect 2518 3523 2519 3540
rect 2377 3546 2378 3549
rect 2383 3546 2384 3549
rect 2389 3546 2390 3549
rect 2392 3546 2393 3549
rect 2395 3546 2396 3549
rect 2454 3546 2455 3549
rect 2409 3546 2410 3551
rect 2431 3546 2432 3551
rect 2441 3546 2442 3551
rect 2448 3546 2449 3551
<< via >>
rect 2359 1121 2360 1122
rect 2372 1121 2373 1122
rect 2375 1121 2376 1122
rect 2378 1121 2379 1122
rect 2384 1121 2385 1122
rect 2387 1121 2388 1122
rect 2467 1121 2468 1122
rect 2473 1121 2474 1122
rect 2361 1131 2362 1132
rect 2399 1131 2400 1132
rect 2375 1133 2376 1134
rect 2387 1133 2388 1134
rect 2384 1135 2385 1136
rect 2409 1135 2410 1136
rect 2372 1137 2373 1138
rect 2384 1137 2385 1138
rect 2372 1139 2373 1140
rect 2396 1139 2397 1140
rect 2390 1141 2391 1142
rect 2435 1141 2436 1142
rect 2369 1143 2370 1144
rect 2390 1143 2391 1144
rect 2419 1143 2420 1144
rect 2438 1143 2439 1144
rect 2422 1145 2423 1146
rect 2464 1145 2465 1146
rect 2441 1147 2442 1148
rect 2491 1147 2492 1148
rect 2467 1149 2468 1150
rect 2526 1149 2527 1150
rect 2354 1158 2355 1159
rect 2418 1158 2419 1159
rect 2368 1160 2369 1161
rect 2477 1160 2478 1161
rect 2375 1162 2376 1163
rect 2393 1162 2394 1163
rect 2384 1164 2385 1165
rect 2430 1164 2431 1165
rect 2387 1166 2388 1167
rect 2433 1166 2434 1167
rect 2390 1168 2391 1169
rect 2424 1168 2425 1169
rect 2397 1170 2398 1171
rect 2412 1170 2413 1171
rect 2402 1172 2403 1173
rect 2412 1172 2413 1173
rect 2421 1172 2422 1173
rect 2565 1172 2566 1173
rect 2426 1174 2427 1175
rect 2438 1174 2439 1175
rect 2399 1176 2400 1177
rect 2439 1176 2440 1177
rect 2435 1178 2436 1179
rect 2472 1178 2473 1179
rect 2323 1180 2324 1181
rect 2436 1180 2437 1181
rect 2441 1180 2442 1181
rect 2478 1180 2479 1181
rect 2458 1182 2459 1183
rect 2475 1182 2476 1183
rect 2461 1184 2462 1185
rect 2466 1184 2467 1185
rect 2464 1186 2465 1187
rect 2510 1186 2511 1187
rect 2470 1188 2471 1189
rect 2513 1188 2514 1189
rect 2481 1190 2482 1191
rect 2498 1190 2499 1191
rect 2495 1192 2496 1193
rect 2525 1192 2526 1193
rect 2505 1194 2506 1195
rect 2548 1194 2549 1195
rect 2516 1196 2517 1197
rect 2596 1196 2597 1197
rect 2327 1205 2328 1206
rect 2392 1205 2393 1206
rect 2397 1205 2398 1206
rect 2401 1205 2402 1206
rect 2412 1205 2413 1206
rect 2416 1205 2417 1206
rect 2424 1205 2425 1206
rect 2428 1205 2429 1206
rect 2421 1207 2422 1208
rect 2425 1207 2426 1208
rect 2418 1209 2419 1210
rect 2422 1209 2423 1210
rect 2439 1209 2440 1210
rect 2443 1209 2444 1210
rect 2436 1211 2437 1212
rect 2440 1211 2441 1212
rect 2433 1213 2434 1214
rect 2437 1213 2438 1214
rect 2430 1215 2431 1216
rect 2434 1215 2435 1216
rect 2466 1215 2467 1216
rect 2470 1215 2471 1216
rect 2481 1215 2482 1216
rect 2485 1215 2486 1216
rect 2478 1217 2479 1218
rect 2482 1217 2483 1218
rect 2475 1219 2476 1220
rect 2479 1219 2480 1220
rect 2472 1221 2473 1222
rect 2476 1221 2477 1222
rect 2510 1221 2511 1222
rect 2522 1221 2523 1222
rect 2516 1223 2517 1224
rect 2534 1223 2535 1224
rect 2525 1225 2526 1226
rect 2528 1225 2529 1226
rect 2513 1227 2514 1228
rect 2525 1227 2526 1228
rect 2548 1227 2549 1228
rect 2553 1227 2554 1228
rect 2547 1229 2548 1230
rect 2583 1229 2584 1230
rect 2550 1231 2551 1232
rect 2568 1231 2569 1232
rect 2586 1231 2587 1232
rect 2622 1231 2623 1232
rect 2595 1233 2596 1234
rect 2619 1233 2620 1234
rect 2317 1242 2318 1243
rect 2392 1242 2393 1243
rect 2325 1244 2326 1245
rect 2339 1244 2340 1245
rect 2332 1246 2333 1247
rect 2465 1246 2466 1247
rect 2335 1248 2336 1249
rect 2459 1248 2460 1249
rect 2395 1250 2396 1251
rect 2468 1250 2469 1251
rect 2398 1252 2399 1253
rect 2401 1252 2402 1253
rect 2411 1252 2412 1253
rect 2416 1252 2417 1253
rect 2417 1254 2418 1255
rect 2428 1254 2429 1255
rect 2314 1256 2315 1257
rect 2429 1256 2430 1257
rect 2432 1258 2433 1259
rect 2437 1258 2438 1259
rect 2434 1260 2435 1261
rect 2462 1260 2463 1261
rect 2435 1262 2436 1263
rect 2440 1262 2441 1263
rect 2443 1262 2444 1263
rect 2450 1262 2451 1263
rect 2476 1262 2477 1263
rect 2489 1262 2490 1263
rect 2470 1264 2471 1265
rect 2477 1264 2478 1265
rect 2479 1264 2480 1265
rect 2492 1264 2493 1265
rect 2482 1266 2483 1267
rect 2495 1266 2496 1267
rect 2485 1268 2486 1269
rect 2498 1268 2499 1269
rect 2522 1268 2523 1269
rect 2547 1268 2548 1269
rect 2528 1270 2529 1271
rect 2544 1270 2545 1271
rect 2386 1272 2387 1273
rect 2529 1272 2530 1273
rect 2534 1272 2535 1273
rect 2556 1272 2557 1273
rect 2550 1274 2551 1275
rect 2565 1274 2566 1275
rect 2525 1276 2526 1277
rect 2550 1276 2551 1277
rect 2501 1278 2502 1279
rect 2526 1278 2527 1279
rect 2553 1278 2554 1279
rect 2574 1278 2575 1279
rect 2531 1280 2532 1281
rect 2553 1280 2554 1281
rect 2583 1280 2584 1281
rect 2662 1280 2663 1281
rect 2586 1282 2587 1283
rect 2615 1282 2616 1283
rect 2595 1284 2596 1285
rect 2633 1284 2634 1285
rect 2618 1286 2619 1287
rect 2665 1286 2666 1287
rect 2636 1288 2637 1289
rect 2649 1288 2650 1289
rect 2659 1288 2660 1289
rect 2675 1288 2676 1289
rect 2314 1297 2315 1298
rect 2318 1297 2319 1298
rect 2323 1297 2324 1298
rect 2330 1297 2331 1298
rect 2325 1299 2326 1300
rect 2429 1299 2430 1300
rect 2349 1301 2350 1302
rect 2593 1301 2594 1302
rect 2357 1303 2358 1304
rect 2642 1303 2643 1304
rect 2360 1305 2361 1306
rect 2486 1305 2487 1306
rect 2403 1307 2404 1308
rect 2411 1307 2412 1308
rect 2409 1309 2410 1310
rect 2423 1309 2424 1310
rect 2412 1311 2413 1312
rect 2426 1311 2427 1312
rect 2415 1313 2416 1314
rect 2417 1313 2418 1314
rect 2421 1313 2422 1314
rect 2432 1313 2433 1314
rect 2424 1315 2425 1316
rect 2435 1315 2436 1316
rect 2433 1317 2434 1318
rect 2450 1317 2451 1318
rect 2367 1319 2368 1320
rect 2451 1319 2452 1320
rect 2442 1321 2443 1322
rect 2465 1321 2466 1322
rect 2444 1323 2445 1324
rect 2462 1323 2463 1324
rect 2448 1325 2449 1326
rect 2459 1325 2460 1326
rect 2464 1325 2465 1326
rect 2492 1325 2493 1326
rect 2468 1327 2469 1328
rect 2477 1327 2478 1328
rect 2471 1329 2472 1330
rect 2526 1329 2527 1330
rect 2480 1331 2481 1332
rect 2498 1331 2499 1332
rect 2492 1333 2493 1334
rect 2495 1333 2496 1334
rect 2501 1333 2502 1334
rect 2516 1333 2517 1334
rect 2504 1335 2505 1336
rect 2529 1335 2530 1336
rect 2507 1337 2508 1338
rect 2550 1337 2551 1338
rect 2531 1339 2532 1340
rect 2544 1339 2545 1340
rect 2534 1341 2535 1342
rect 2553 1341 2554 1342
rect 2537 1343 2538 1344
rect 2556 1343 2557 1344
rect 2549 1345 2550 1346
rect 2559 1345 2560 1346
rect 2474 1347 2475 1348
rect 2558 1347 2559 1348
rect 2552 1349 2553 1350
rect 2565 1349 2566 1350
rect 2561 1351 2562 1352
rect 2574 1351 2575 1352
rect 2602 1351 2603 1352
rect 2636 1351 2637 1352
rect 2605 1353 2606 1354
rect 2621 1353 2622 1354
rect 2615 1355 2616 1356
rect 2665 1355 2666 1356
rect 2584 1357 2585 1358
rect 2615 1357 2616 1358
rect 2618 1357 2619 1358
rect 2642 1357 2643 1358
rect 2633 1359 2634 1360
rect 2649 1359 2650 1360
rect 2632 1361 2633 1362
rect 2659 1361 2660 1362
rect 2645 1363 2646 1364
rect 2662 1363 2663 1364
rect 2323 1372 2324 1373
rect 2381 1372 2382 1373
rect 2351 1374 2352 1375
rect 2393 1374 2394 1375
rect 2357 1376 2358 1377
rect 2378 1376 2379 1377
rect 2372 1378 2373 1379
rect 2421 1378 2422 1379
rect 2375 1380 2376 1381
rect 2415 1380 2416 1381
rect 2403 1382 2404 1383
rect 2426 1382 2427 1383
rect 2409 1384 2410 1385
rect 2414 1384 2415 1385
rect 2399 1386 2400 1387
rect 2408 1386 2409 1387
rect 2412 1386 2413 1387
rect 2417 1386 2418 1387
rect 2424 1386 2425 1387
rect 2429 1386 2430 1387
rect 2433 1386 2434 1387
rect 2438 1386 2439 1387
rect 2448 1386 2449 1387
rect 2453 1386 2454 1387
rect 2442 1388 2443 1389
rect 2447 1388 2448 1389
rect 2451 1388 2452 1389
rect 2456 1388 2457 1389
rect 2471 1388 2472 1389
rect 2498 1388 2499 1389
rect 2477 1390 2478 1391
rect 2480 1390 2481 1391
rect 2474 1392 2475 1393
rect 2477 1392 2478 1393
rect 2483 1392 2484 1393
rect 2489 1392 2490 1393
rect 2486 1394 2487 1395
rect 2489 1394 2490 1395
rect 2492 1394 2493 1395
rect 2495 1394 2496 1395
rect 2464 1396 2465 1397
rect 2492 1396 2493 1397
rect 2507 1396 2508 1397
rect 2510 1396 2511 1397
rect 2504 1398 2505 1399
rect 2507 1398 2508 1399
rect 2504 1400 2505 1401
rect 2516 1400 2517 1401
rect 2513 1402 2514 1403
rect 2587 1402 2588 1403
rect 2534 1404 2535 1405
rect 2543 1404 2544 1405
rect 2531 1406 2532 1407
rect 2534 1406 2535 1407
rect 2564 1406 2565 1407
rect 2608 1406 2609 1407
rect 2581 1408 2582 1409
rect 2630 1408 2631 1409
rect 2561 1410 2562 1411
rect 2580 1410 2581 1411
rect 2552 1412 2553 1413
rect 2561 1412 2562 1413
rect 2549 1414 2550 1415
rect 2552 1414 2553 1415
rect 2546 1416 2547 1417
rect 2549 1416 2550 1417
rect 2537 1418 2538 1419
rect 2546 1418 2547 1419
rect 2584 1418 2585 1419
rect 2615 1418 2616 1419
rect 2501 1420 2502 1421
rect 2583 1420 2584 1421
rect 2593 1420 2594 1421
rect 2608 1420 2609 1421
rect 2632 1420 2633 1421
rect 2655 1420 2656 1421
rect 2602 1422 2603 1423
rect 2633 1422 2634 1423
rect 2602 1424 2603 1425
rect 2665 1424 2666 1425
rect 2635 1426 2636 1427
rect 2649 1426 2650 1427
rect 2638 1428 2639 1429
rect 2675 1428 2676 1429
rect 2652 1430 2653 1431
rect 2668 1430 2669 1431
rect 2290 1439 2291 1440
rect 2384 1439 2385 1440
rect 2304 1441 2305 1442
rect 2308 1441 2309 1442
rect 2329 1441 2330 1442
rect 2402 1441 2403 1442
rect 2343 1443 2344 1444
rect 2486 1443 2487 1444
rect 2350 1445 2351 1446
rect 2411 1445 2412 1446
rect 2357 1447 2358 1448
rect 2417 1447 2418 1448
rect 2365 1449 2366 1450
rect 2453 1449 2454 1450
rect 2372 1451 2373 1452
rect 2426 1451 2427 1452
rect 2378 1453 2379 1454
rect 2417 1453 2418 1454
rect 2381 1455 2382 1456
rect 2399 1455 2400 1456
rect 2323 1457 2324 1458
rect 2399 1457 2400 1458
rect 2414 1457 2415 1458
rect 2435 1457 2436 1458
rect 2333 1459 2334 1460
rect 2414 1459 2415 1460
rect 2432 1459 2433 1460
rect 2456 1459 2457 1460
rect 2438 1461 2439 1462
rect 2450 1461 2451 1462
rect 2393 1463 2394 1464
rect 2438 1463 2439 1464
rect 2447 1463 2448 1464
rect 2465 1463 2466 1464
rect 2429 1465 2430 1466
rect 2447 1465 2448 1466
rect 2453 1465 2454 1466
rect 2480 1465 2481 1466
rect 2471 1467 2472 1468
rect 2555 1467 2556 1468
rect 2495 1469 2496 1470
rect 2531 1469 2532 1470
rect 2489 1471 2490 1472
rect 2495 1471 2496 1472
rect 2483 1473 2484 1474
rect 2489 1473 2490 1474
rect 2477 1475 2478 1476
rect 2483 1475 2484 1476
rect 2498 1475 2499 1476
rect 2519 1475 2520 1476
rect 2507 1477 2508 1478
rect 2528 1477 2529 1478
rect 2492 1479 2493 1480
rect 2507 1479 2508 1480
rect 2510 1479 2511 1480
rect 2522 1479 2523 1480
rect 2504 1481 2505 1482
rect 2510 1481 2511 1482
rect 2549 1481 2550 1482
rect 2597 1481 2598 1482
rect 2552 1483 2553 1484
rect 2600 1483 2601 1484
rect 2516 1485 2517 1486
rect 2552 1485 2553 1486
rect 2561 1485 2562 1486
rect 2573 1485 2574 1486
rect 2543 1487 2544 1488
rect 2561 1487 2562 1488
rect 2534 1489 2535 1490
rect 2543 1489 2544 1490
rect 2534 1491 2535 1492
rect 2549 1491 2550 1492
rect 2564 1491 2565 1492
rect 2567 1491 2568 1492
rect 2546 1493 2547 1494
rect 2564 1493 2565 1494
rect 2580 1493 2581 1494
rect 2594 1493 2595 1494
rect 2583 1495 2584 1496
rect 2590 1495 2591 1496
rect 2591 1497 2592 1498
rect 2611 1497 2612 1498
rect 2608 1499 2609 1500
rect 2615 1499 2616 1500
rect 2630 1499 2631 1500
rect 2668 1499 2669 1500
rect 2633 1501 2634 1502
rect 2671 1501 2672 1502
rect 2649 1503 2650 1504
rect 2687 1503 2688 1504
rect 2650 1505 2651 1506
rect 2684 1505 2685 1506
rect 2652 1507 2653 1508
rect 2690 1507 2691 1508
rect 2653 1509 2654 1510
rect 2659 1509 2660 1510
rect 2655 1511 2656 1512
rect 2693 1511 2694 1512
rect 2287 1520 2288 1521
rect 2301 1520 2302 1521
rect 2297 1522 2298 1523
rect 2384 1522 2385 1523
rect 2308 1524 2309 1525
rect 2423 1524 2424 1525
rect 2311 1526 2312 1527
rect 2315 1526 2316 1527
rect 2353 1526 2354 1527
rect 2411 1526 2412 1527
rect 2370 1528 2371 1529
rect 2498 1528 2499 1529
rect 2374 1530 2375 1531
rect 2447 1530 2448 1531
rect 2393 1532 2394 1533
rect 2402 1532 2403 1533
rect 2332 1534 2333 1535
rect 2402 1534 2403 1535
rect 2411 1534 2412 1535
rect 2471 1534 2472 1535
rect 2417 1536 2418 1537
rect 2420 1536 2421 1537
rect 2414 1538 2415 1539
rect 2417 1538 2418 1539
rect 2432 1538 2433 1539
rect 2501 1538 2502 1539
rect 2438 1540 2439 1541
rect 2456 1540 2457 1541
rect 2438 1542 2439 1543
rect 2486 1542 2487 1543
rect 2450 1544 2451 1545
rect 2486 1544 2487 1545
rect 2322 1546 2323 1547
rect 2450 1546 2451 1547
rect 2321 1548 2322 1549
rect 2471 1548 2472 1549
rect 2459 1550 2460 1551
rect 2477 1550 2478 1551
rect 2465 1552 2466 1553
rect 2480 1552 2481 1553
rect 2453 1554 2454 1555
rect 2465 1554 2466 1555
rect 2435 1556 2436 1557
rect 2453 1556 2454 1557
rect 2483 1556 2484 1557
rect 2524 1556 2525 1557
rect 2489 1558 2490 1559
rect 2504 1558 2505 1559
rect 2367 1560 2368 1561
rect 2489 1560 2490 1561
rect 2367 1562 2368 1563
rect 2492 1562 2493 1563
rect 2495 1562 2496 1563
rect 2536 1562 2537 1563
rect 2510 1564 2511 1565
rect 2513 1564 2514 1565
rect 2507 1566 2508 1567
rect 2514 1566 2515 1567
rect 2507 1568 2508 1569
rect 2706 1568 2707 1569
rect 2519 1570 2520 1571
rect 2557 1570 2558 1571
rect 2522 1572 2523 1573
rect 2569 1572 2570 1573
rect 2528 1574 2529 1575
rect 2575 1574 2576 1575
rect 2360 1576 2361 1577
rect 2527 1576 2528 1577
rect 2534 1576 2535 1577
rect 2539 1576 2540 1577
rect 2543 1576 2544 1577
rect 2696 1576 2697 1577
rect 2531 1578 2532 1579
rect 2542 1578 2543 1579
rect 2552 1578 2553 1579
rect 2581 1578 2582 1579
rect 2567 1580 2568 1581
rect 2611 1580 2612 1581
rect 2573 1582 2574 1583
rect 2617 1582 2618 1583
rect 2578 1584 2579 1585
rect 2585 1584 2586 1585
rect 2591 1584 2592 1585
rect 2608 1584 2609 1585
rect 2594 1586 2595 1587
rect 2629 1586 2630 1587
rect 2597 1588 2598 1589
rect 2623 1588 2624 1589
rect 2561 1590 2562 1591
rect 2596 1590 2597 1591
rect 2560 1592 2561 1593
rect 2625 1592 2626 1593
rect 2600 1594 2601 1595
rect 2626 1594 2627 1595
rect 2564 1596 2565 1597
rect 2599 1596 2600 1597
rect 2615 1596 2616 1597
rect 2664 1596 2665 1597
rect 2653 1598 2654 1599
rect 2658 1598 2659 1599
rect 2656 1600 2657 1601
rect 2709 1600 2710 1601
rect 2668 1602 2669 1603
rect 2700 1602 2701 1603
rect 2671 1604 2672 1605
rect 2703 1604 2704 1605
rect 2670 1606 2671 1607
rect 2697 1606 2698 1607
rect 2685 1608 2686 1609
rect 2779 1608 2780 1609
rect 2687 1610 2688 1611
rect 2718 1610 2719 1611
rect 2690 1612 2691 1613
rect 2721 1612 2722 1613
rect 2693 1614 2694 1615
rect 2744 1614 2745 1615
rect 2650 1616 2651 1617
rect 2694 1616 2695 1617
rect 2649 1618 2650 1619
rect 2667 1618 2668 1619
rect 2724 1618 2725 1619
rect 2792 1618 2793 1619
rect 2765 1620 2766 1621
rect 2772 1620 2773 1621
rect 2311 1629 2312 1630
rect 2450 1629 2451 1630
rect 2312 1631 2313 1632
rect 2423 1631 2424 1632
rect 2325 1633 2326 1634
rect 2510 1633 2511 1634
rect 2326 1635 2327 1636
rect 2646 1635 2647 1636
rect 2340 1637 2341 1638
rect 2411 1637 2412 1638
rect 2353 1639 2354 1640
rect 2367 1639 2368 1640
rect 2368 1641 2369 1642
rect 2498 1641 2499 1642
rect 2375 1643 2376 1644
rect 2489 1643 2490 1644
rect 2414 1645 2415 1646
rect 2516 1645 2517 1646
rect 2420 1647 2421 1648
rect 2423 1647 2424 1648
rect 2417 1649 2418 1650
rect 2420 1649 2421 1650
rect 2417 1651 2418 1652
rect 2492 1651 2493 1652
rect 2438 1653 2439 1654
rect 2450 1653 2451 1654
rect 2453 1653 2454 1654
rect 2462 1653 2463 1654
rect 2459 1655 2460 1656
rect 2581 1655 2582 1656
rect 2319 1657 2320 1658
rect 2459 1657 2460 1658
rect 2465 1657 2466 1658
rect 2474 1657 2475 1658
rect 2456 1659 2457 1660
rect 2465 1659 2466 1660
rect 2314 1661 2315 1662
rect 2456 1661 2457 1662
rect 2480 1661 2481 1662
rect 2495 1661 2496 1662
rect 2471 1663 2472 1664
rect 2480 1663 2481 1664
rect 2483 1663 2484 1664
rect 2501 1663 2502 1664
rect 2384 1665 2385 1666
rect 2501 1665 2502 1666
rect 2486 1667 2487 1668
rect 2492 1667 2493 1668
rect 2507 1667 2508 1668
rect 2778 1667 2779 1668
rect 2518 1669 2519 1670
rect 2546 1669 2547 1670
rect 2522 1671 2523 1672
rect 2524 1671 2525 1672
rect 2525 1673 2526 1674
rect 2527 1673 2528 1674
rect 2531 1673 2532 1674
rect 2534 1673 2535 1674
rect 2539 1673 2540 1674
rect 2681 1673 2682 1674
rect 2536 1675 2537 1676
rect 2540 1675 2541 1676
rect 2477 1677 2478 1678
rect 2537 1677 2538 1678
rect 2552 1677 2553 1678
rect 2560 1677 2561 1678
rect 2557 1679 2558 1680
rect 2567 1679 2568 1680
rect 2569 1679 2570 1680
rect 2573 1679 2574 1680
rect 2570 1681 2571 1682
rect 2575 1681 2576 1682
rect 2578 1681 2579 1682
rect 2591 1681 2592 1682
rect 2564 1683 2565 1684
rect 2579 1683 2580 1684
rect 2599 1683 2600 1684
rect 2603 1683 2604 1684
rect 2596 1685 2597 1686
rect 2600 1685 2601 1686
rect 2608 1685 2609 1686
rect 2642 1685 2643 1686
rect 2626 1687 2627 1688
rect 2633 1687 2634 1688
rect 2629 1689 2630 1690
rect 2636 1689 2637 1690
rect 2623 1691 2624 1692
rect 2630 1691 2631 1692
rect 2639 1691 2640 1692
rect 2771 1691 2772 1692
rect 2651 1693 2652 1694
rect 2721 1693 2722 1694
rect 2660 1695 2661 1696
rect 2664 1695 2665 1696
rect 2675 1695 2676 1696
rect 2730 1695 2731 1696
rect 2697 1697 2698 1698
rect 2740 1697 2741 1698
rect 2694 1699 2695 1700
rect 2696 1699 2697 1700
rect 2693 1701 2694 1702
rect 2755 1701 2756 1702
rect 2700 1703 2701 1704
rect 2751 1703 2752 1704
rect 2658 1705 2659 1706
rect 2699 1705 2700 1706
rect 2703 1705 2704 1706
rect 2711 1705 2712 1706
rect 2706 1707 2707 1708
rect 2720 1707 2721 1708
rect 2718 1709 2719 1710
rect 2734 1709 2735 1710
rect 2724 1711 2725 1712
rect 2786 1711 2787 1712
rect 2709 1713 2710 1714
rect 2723 1713 2724 1714
rect 2708 1715 2709 1716
rect 2748 1715 2749 1716
rect 2792 1715 2793 1716
rect 2799 1715 2800 1716
rect 2312 1724 2313 1725
rect 2459 1724 2460 1725
rect 2323 1726 2324 1727
rect 2330 1726 2331 1727
rect 2326 1728 2327 1729
rect 2453 1728 2454 1729
rect 2341 1730 2342 1731
rect 2444 1730 2445 1731
rect 2369 1732 2370 1733
rect 2474 1732 2475 1733
rect 2375 1734 2376 1735
rect 2426 1734 2427 1735
rect 2417 1736 2418 1737
rect 2501 1736 2502 1737
rect 2447 1738 2448 1739
rect 2462 1738 2463 1739
rect 2450 1740 2451 1741
rect 2462 1740 2463 1741
rect 2417 1742 2418 1743
rect 2450 1742 2451 1743
rect 2456 1742 2457 1743
rect 2459 1742 2460 1743
rect 2402 1744 2403 1745
rect 2456 1744 2457 1745
rect 2465 1744 2466 1745
rect 2468 1744 2469 1745
rect 2471 1744 2472 1745
rect 2516 1744 2517 1745
rect 2474 1746 2475 1747
rect 2480 1746 2481 1747
rect 2477 1748 2478 1749
rect 2483 1748 2484 1749
rect 2486 1748 2487 1749
rect 2495 1748 2496 1749
rect 2501 1748 2502 1749
rect 2510 1748 2511 1749
rect 2355 1750 2356 1751
rect 2510 1750 2511 1751
rect 2507 1752 2508 1753
rect 2513 1752 2514 1753
rect 2299 1754 2300 1755
rect 2507 1754 2508 1755
rect 2537 1754 2538 1755
rect 2549 1754 2550 1755
rect 2525 1756 2526 1757
rect 2537 1756 2538 1757
rect 2543 1756 2544 1757
rect 2561 1756 2562 1757
rect 2552 1758 2553 1759
rect 2579 1758 2580 1759
rect 2558 1760 2559 1761
rect 2760 1760 2761 1761
rect 2564 1762 2565 1763
rect 2576 1762 2577 1763
rect 2546 1764 2547 1765
rect 2564 1764 2565 1765
rect 2534 1766 2535 1767
rect 2546 1766 2547 1767
rect 2522 1768 2523 1769
rect 2534 1768 2535 1769
rect 2522 1770 2523 1771
rect 2540 1770 2541 1771
rect 2567 1770 2568 1771
rect 2582 1770 2583 1771
rect 2573 1772 2574 1773
rect 2594 1772 2595 1773
rect 2591 1774 2592 1775
rect 2606 1774 2607 1775
rect 2603 1776 2604 1777
rect 2715 1776 2716 1777
rect 2570 1778 2571 1779
rect 2603 1778 2604 1779
rect 2630 1778 2631 1779
rect 2654 1778 2655 1779
rect 2630 1780 2631 1781
rect 2657 1780 2658 1781
rect 2633 1782 2634 1783
rect 2687 1782 2688 1783
rect 2612 1784 2613 1785
rect 2633 1784 2634 1785
rect 2639 1784 2640 1785
rect 2669 1784 2670 1785
rect 2618 1786 2619 1787
rect 2639 1786 2640 1787
rect 2651 1786 2652 1787
rect 2736 1786 2737 1787
rect 2636 1788 2637 1789
rect 2651 1788 2652 1789
rect 2672 1788 2673 1789
rect 2681 1788 2682 1789
rect 2642 1790 2643 1791
rect 2672 1790 2673 1791
rect 2660 1792 2661 1793
rect 2681 1792 2682 1793
rect 2600 1794 2601 1795
rect 2660 1794 2661 1795
rect 2600 1796 2601 1797
rect 2645 1796 2646 1797
rect 2675 1796 2676 1797
rect 2705 1796 2706 1797
rect 2684 1798 2685 1799
rect 2739 1798 2740 1799
rect 2627 1800 2628 1801
rect 2684 1800 2685 1801
rect 2693 1800 2694 1801
rect 2751 1800 2752 1801
rect 2696 1802 2697 1803
rect 2766 1802 2767 1803
rect 2696 1804 2697 1805
rect 2819 1804 2820 1805
rect 2699 1806 2700 1807
rect 2769 1806 2770 1807
rect 2708 1808 2709 1809
rect 2778 1808 2779 1809
rect 2528 1810 2529 1811
rect 2708 1810 2709 1811
rect 2711 1810 2712 1811
rect 2781 1810 2782 1811
rect 2720 1812 2721 1813
rect 2796 1812 2797 1813
rect 2702 1814 2703 1815
rect 2721 1814 2722 1815
rect 2723 1814 2724 1815
rect 2784 1814 2785 1815
rect 2729 1816 2730 1817
rect 2799 1816 2800 1817
rect 2733 1818 2734 1819
rect 2771 1818 2772 1819
rect 2724 1820 2725 1821
rect 2772 1820 2773 1821
rect 2742 1822 2743 1823
rect 2747 1822 2748 1823
rect 2754 1822 2755 1823
rect 2812 1822 2813 1823
rect 2757 1824 2758 1825
rect 2809 1824 2810 1825
rect 2302 1833 2303 1834
rect 2306 1833 2307 1834
rect 2316 1833 2317 1834
rect 2459 1833 2460 1834
rect 2320 1835 2321 1836
rect 2442 1835 2443 1836
rect 2330 1837 2331 1838
rect 2406 1837 2407 1838
rect 2337 1839 2338 1840
rect 2423 1839 2424 1840
rect 2358 1841 2359 1842
rect 2687 1841 2688 1842
rect 2362 1843 2363 1844
rect 2781 1843 2782 1844
rect 2381 1845 2382 1846
rect 2393 1845 2394 1846
rect 2391 1847 2392 1848
rect 2399 1847 2400 1848
rect 2403 1847 2404 1848
rect 2411 1847 2412 1848
rect 2412 1849 2413 1850
rect 2528 1849 2529 1850
rect 2415 1851 2416 1852
rect 2532 1851 2533 1852
rect 2418 1853 2419 1854
rect 2420 1853 2421 1854
rect 2433 1853 2434 1854
rect 2462 1853 2463 1854
rect 2439 1855 2440 1856
rect 2444 1855 2445 1856
rect 2456 1855 2457 1856
rect 2460 1855 2461 1856
rect 2453 1857 2454 1858
rect 2457 1857 2458 1858
rect 2450 1859 2451 1860
rect 2454 1859 2455 1860
rect 2447 1861 2448 1862
rect 2451 1861 2452 1862
rect 2469 1861 2470 1862
rect 2523 1861 2524 1862
rect 2481 1863 2482 1864
rect 2486 1863 2487 1864
rect 2487 1865 2488 1866
rect 2501 1865 2502 1866
rect 2492 1867 2493 1868
rect 2499 1867 2500 1868
rect 2493 1869 2494 1870
rect 2516 1869 2517 1870
rect 2471 1871 2472 1872
rect 2517 1871 2518 1872
rect 2537 1871 2538 1872
rect 2541 1871 2542 1872
rect 2534 1873 2535 1874
rect 2538 1873 2539 1874
rect 2544 1873 2545 1874
rect 2561 1873 2562 1874
rect 2549 1875 2550 1876
rect 2553 1875 2554 1876
rect 2546 1877 2547 1878
rect 2550 1877 2551 1878
rect 2556 1877 2557 1878
rect 2558 1877 2559 1878
rect 2313 1879 2314 1880
rect 2559 1879 2560 1880
rect 2564 1879 2565 1880
rect 2574 1879 2575 1880
rect 2600 1879 2601 1880
rect 2693 1879 2694 1880
rect 2603 1881 2604 1882
rect 2613 1881 2614 1882
rect 2604 1883 2605 1884
rect 2676 1883 2677 1884
rect 2610 1885 2611 1886
rect 2690 1885 2691 1886
rect 2594 1887 2595 1888
rect 2691 1887 2692 1888
rect 2627 1889 2628 1890
rect 2631 1889 2632 1890
rect 2606 1891 2607 1892
rect 2628 1891 2629 1892
rect 2576 1893 2577 1894
rect 2607 1893 2608 1894
rect 2651 1893 2652 1894
rect 2744 1893 2745 1894
rect 2681 1895 2682 1896
rect 2694 1895 2695 1896
rect 2684 1897 2685 1898
rect 2688 1897 2689 1898
rect 2696 1897 2697 1898
rect 2781 1897 2782 1898
rect 2711 1899 2712 1900
rect 2742 1899 2743 1900
rect 2714 1901 2715 1902
rect 2763 1901 2764 1902
rect 2717 1903 2718 1904
rect 2721 1903 2722 1904
rect 2720 1905 2721 1906
rect 2733 1905 2734 1906
rect 2724 1907 2725 1908
rect 2759 1907 2760 1908
rect 2723 1909 2724 1910
rect 2736 1909 2737 1910
rect 2726 1911 2727 1912
rect 2739 1911 2740 1912
rect 2729 1913 2730 1914
rect 2833 1913 2834 1914
rect 2741 1915 2742 1916
rect 2754 1915 2755 1916
rect 2751 1917 2752 1918
rect 2771 1917 2772 1918
rect 2753 1919 2754 1920
rect 2766 1919 2767 1920
rect 2757 1921 2758 1922
rect 2762 1921 2763 1922
rect 2639 1923 2640 1924
rect 2756 1923 2757 1924
rect 2633 1925 2634 1926
rect 2640 1925 2641 1926
rect 2765 1925 2766 1926
rect 2796 1925 2797 1926
rect 2769 1927 2770 1928
rect 2816 1927 2817 1928
rect 2768 1929 2769 1930
rect 2819 1929 2820 1930
rect 2778 1931 2779 1932
rect 2847 1931 2848 1932
rect 2777 1933 2778 1934
rect 2812 1933 2813 1934
rect 2732 1935 2733 1936
rect 2812 1935 2813 1936
rect 2784 1937 2785 1938
rect 2802 1937 2803 1938
rect 2799 1939 2800 1940
rect 2805 1939 2806 1940
rect 2302 1948 2303 1949
rect 2426 1948 2427 1949
rect 2309 1950 2310 1951
rect 2429 1950 2430 1951
rect 2317 1952 2318 1953
rect 2389 1952 2390 1953
rect 2320 1954 2321 1955
rect 2445 1954 2446 1955
rect 2324 1956 2325 1957
rect 2400 1956 2401 1957
rect 2323 1958 2324 1959
rect 2495 1958 2496 1959
rect 2345 1960 2346 1961
rect 2514 1960 2515 1961
rect 2348 1962 2349 1963
rect 2691 1962 2692 1963
rect 2359 1964 2360 1965
rect 2546 1964 2547 1965
rect 2366 1966 2367 1967
rect 2391 1966 2392 1967
rect 2397 1966 2398 1967
rect 2532 1966 2533 1967
rect 2403 1968 2404 1969
rect 2501 1968 2502 1969
rect 2402 1970 2403 1971
rect 2460 1970 2461 1971
rect 2406 1972 2407 1973
rect 2420 1972 2421 1973
rect 2439 1972 2440 1973
rect 2459 1972 2460 1973
rect 2418 1974 2419 1975
rect 2438 1974 2439 1975
rect 2465 1974 2466 1975
rect 2550 1974 2551 1975
rect 2469 1976 2470 1977
rect 2622 1976 2623 1977
rect 2478 1978 2479 1979
rect 2513 1978 2514 1979
rect 2454 1980 2455 1981
rect 2477 1980 2478 1981
rect 2433 1982 2434 1983
rect 2453 1982 2454 1983
rect 2380 1984 2381 1985
rect 2432 1984 2433 1985
rect 2487 1984 2488 1985
rect 2528 1984 2529 1985
rect 2493 1986 2494 1987
rect 2534 1986 2535 1987
rect 2457 1988 2458 1989
rect 2492 1988 2493 1989
rect 2508 1988 2509 1989
rect 2549 1988 2550 1989
rect 2442 1990 2443 1991
rect 2507 1990 2508 1991
rect 2351 1992 2352 1993
rect 2441 1992 2442 1993
rect 2517 1992 2518 1993
rect 2565 1992 2566 1993
rect 2504 1994 2505 1995
rect 2516 1994 2517 1995
rect 2523 1994 2524 1995
rect 2567 1994 2568 1995
rect 2481 1996 2482 1997
rect 2522 1996 2523 1997
rect 2538 1996 2539 1997
rect 2570 1996 2571 1997
rect 2537 1998 2538 1999
rect 2553 1998 2554 1999
rect 2544 2000 2545 2001
rect 2576 2000 2577 2001
rect 2499 2002 2500 2003
rect 2543 2002 2544 2003
rect 2337 2004 2338 2005
rect 2498 2004 2499 2005
rect 2556 2004 2557 2005
rect 2582 2004 2583 2005
rect 2559 2006 2560 2007
rect 2585 2006 2586 2007
rect 2564 2008 2565 2009
rect 2697 2008 2698 2009
rect 2574 2010 2575 2011
rect 2600 2010 2601 2011
rect 2541 2012 2542 2013
rect 2573 2012 2574 2013
rect 2511 2014 2512 2015
rect 2540 2014 2541 2015
rect 2475 2016 2476 2017
rect 2510 2016 2511 2017
rect 2451 2018 2452 2019
rect 2474 2018 2475 2019
rect 2604 2018 2605 2019
rect 2625 2018 2626 2019
rect 2610 2020 2611 2021
rect 2642 2020 2643 2021
rect 2613 2022 2614 2023
rect 2645 2022 2646 2023
rect 2607 2024 2608 2025
rect 2612 2024 2613 2025
rect 2580 2026 2581 2027
rect 2606 2026 2607 2027
rect 2615 2026 2616 2027
rect 2778 2026 2779 2027
rect 2628 2028 2629 2029
rect 2654 2028 2655 2029
rect 2648 2030 2649 2031
rect 2661 2030 2662 2031
rect 2640 2032 2641 2033
rect 2660 2032 2661 2033
rect 2658 2034 2659 2035
rect 2705 2034 2706 2035
rect 2631 2036 2632 2037
rect 2657 2036 2658 2037
rect 2670 2036 2671 2037
rect 2696 2036 2697 2037
rect 2673 2038 2674 2039
rect 2699 2038 2700 2039
rect 2672 2040 2673 2041
rect 2797 2040 2798 2041
rect 2694 2042 2695 2043
rect 2714 2042 2715 2043
rect 2702 2044 2703 2045
rect 2851 2044 2852 2045
rect 2708 2046 2709 2047
rect 2723 2046 2724 2047
rect 2720 2048 2721 2049
rect 2748 2048 2749 2049
rect 2676 2050 2677 2051
rect 2720 2050 2721 2051
rect 2726 2050 2727 2051
rect 2763 2050 2764 2051
rect 2729 2052 2730 2053
rect 2760 2052 2761 2053
rect 2732 2054 2733 2055
rect 2805 2054 2806 2055
rect 2636 2056 2637 2057
rect 2732 2056 2733 2057
rect 2751 2056 2752 2057
rect 2845 2056 2846 2057
rect 2765 2058 2766 2059
rect 2794 2058 2795 2059
rect 2768 2060 2769 2061
rect 2791 2060 2792 2061
rect 2771 2062 2772 2063
rect 2774 2062 2775 2063
rect 2753 2064 2754 2065
rect 2772 2064 2773 2065
rect 2741 2066 2742 2067
rect 2754 2066 2755 2067
rect 2756 2066 2757 2067
rect 2775 2066 2776 2067
rect 2744 2068 2745 2069
rect 2757 2068 2758 2069
rect 2717 2070 2718 2071
rect 2745 2070 2746 2071
rect 2688 2072 2689 2073
rect 2717 2072 2718 2073
rect 2812 2072 2813 2073
rect 2816 2072 2817 2073
rect 2817 2074 2818 2075
rect 2824 2074 2825 2075
rect 2294 2083 2295 2084
rect 2456 2083 2457 2084
rect 2301 2085 2302 2086
rect 2426 2085 2427 2086
rect 2306 2087 2307 2088
rect 2462 2087 2463 2088
rect 2315 2089 2316 2090
rect 2429 2089 2430 2090
rect 2308 2091 2309 2092
rect 2429 2091 2430 2092
rect 2324 2093 2325 2094
rect 2516 2093 2517 2094
rect 2344 2095 2345 2096
rect 2441 2095 2442 2096
rect 2351 2097 2352 2098
rect 2432 2097 2433 2098
rect 2299 2099 2300 2100
rect 2432 2099 2433 2100
rect 2347 2101 2348 2102
rect 2350 2101 2351 2102
rect 2357 2101 2358 2102
rect 2477 2101 2478 2102
rect 2375 2103 2376 2104
rect 2495 2103 2496 2104
rect 2377 2105 2378 2106
rect 2507 2105 2508 2106
rect 2392 2107 2393 2108
rect 2567 2107 2568 2108
rect 2336 2109 2337 2110
rect 2393 2109 2394 2110
rect 2396 2109 2397 2110
rect 2537 2109 2538 2110
rect 2399 2111 2400 2112
rect 2420 2111 2421 2112
rect 2402 2113 2403 2114
rect 2486 2113 2487 2114
rect 2414 2115 2415 2116
rect 2552 2115 2553 2116
rect 2438 2117 2439 2118
rect 2519 2117 2520 2118
rect 2447 2119 2448 2120
rect 2459 2119 2460 2120
rect 2287 2121 2288 2122
rect 2459 2121 2460 2122
rect 2453 2123 2454 2124
rect 2477 2123 2478 2124
rect 2471 2125 2472 2126
rect 2474 2125 2475 2126
rect 2354 2127 2355 2128
rect 2474 2127 2475 2128
rect 2483 2127 2484 2128
rect 2492 2127 2493 2128
rect 2489 2129 2490 2130
rect 2498 2129 2499 2130
rect 2501 2129 2502 2130
rect 2507 2129 2508 2130
rect 2501 2131 2502 2132
rect 2504 2131 2505 2132
rect 2275 2133 2276 2134
rect 2504 2133 2505 2134
rect 2528 2133 2529 2134
rect 2558 2133 2559 2134
rect 2534 2135 2535 2136
rect 2555 2135 2556 2136
rect 2534 2137 2535 2138
rect 2543 2137 2544 2138
rect 2537 2139 2538 2140
rect 2546 2139 2547 2140
rect 2564 2139 2565 2140
rect 2567 2139 2568 2140
rect 2576 2139 2577 2140
rect 2627 2139 2628 2140
rect 2585 2141 2586 2142
rect 2591 2141 2592 2142
rect 2588 2143 2589 2144
rect 2879 2143 2880 2144
rect 2594 2145 2595 2146
rect 2600 2145 2601 2146
rect 2606 2145 2607 2146
rect 2630 2145 2631 2146
rect 2606 2147 2607 2148
rect 2612 2147 2613 2148
rect 2609 2149 2610 2150
rect 2615 2149 2616 2150
rect 2630 2149 2631 2150
rect 2739 2149 2740 2150
rect 2639 2151 2640 2152
rect 2645 2151 2646 2152
rect 2654 2151 2655 2152
rect 2666 2151 2667 2152
rect 2654 2153 2655 2154
rect 2660 2153 2661 2154
rect 2657 2155 2658 2156
rect 2732 2155 2733 2156
rect 2669 2157 2670 2158
rect 2723 2157 2724 2158
rect 2672 2159 2673 2160
rect 2770 2159 2771 2160
rect 2672 2161 2673 2162
rect 2817 2161 2818 2162
rect 2684 2163 2685 2164
rect 2757 2163 2758 2164
rect 2699 2165 2700 2166
rect 2711 2165 2712 2166
rect 2705 2167 2706 2168
rect 2720 2167 2721 2168
rect 2717 2169 2718 2170
rect 2729 2169 2730 2170
rect 2702 2171 2703 2172
rect 2717 2171 2718 2172
rect 2735 2171 2736 2172
rect 2782 2171 2783 2172
rect 2751 2173 2752 2174
rect 2824 2173 2825 2174
rect 2748 2175 2749 2176
rect 2752 2175 2753 2176
rect 2754 2175 2755 2176
rect 2767 2175 2768 2176
rect 2708 2177 2709 2178
rect 2755 2177 2756 2178
rect 2696 2179 2697 2180
rect 2708 2179 2709 2180
rect 2696 2181 2697 2182
rect 2807 2181 2808 2182
rect 2763 2183 2764 2184
rect 2837 2183 2838 2184
rect 2760 2185 2761 2186
rect 2764 2185 2765 2186
rect 2772 2185 2773 2186
rect 2785 2185 2786 2186
rect 2745 2187 2746 2188
rect 2773 2187 2774 2188
rect 2636 2189 2637 2190
rect 2746 2189 2747 2190
rect 2636 2191 2637 2192
rect 2642 2191 2643 2192
rect 2642 2193 2643 2194
rect 2648 2193 2649 2194
rect 2775 2193 2776 2194
rect 2788 2193 2789 2194
rect 2791 2193 2792 2194
rect 2804 2193 2805 2194
rect 2794 2195 2795 2196
rect 2807 2195 2808 2196
rect 2797 2197 2798 2198
rect 2810 2197 2811 2198
rect 2816 2197 2817 2198
rect 2820 2197 2821 2198
rect 2840 2197 2841 2198
rect 2876 2197 2877 2198
rect 2288 2206 2289 2207
rect 2456 2206 2457 2207
rect 2291 2208 2292 2209
rect 2436 2208 2437 2209
rect 2301 2210 2302 2211
rect 2429 2210 2430 2211
rect 2304 2212 2305 2213
rect 2462 2212 2463 2213
rect 2305 2214 2306 2215
rect 2457 2214 2458 2215
rect 2309 2216 2310 2217
rect 2432 2216 2433 2217
rect 2318 2218 2319 2219
rect 2499 2218 2500 2219
rect 2333 2220 2334 2221
rect 2486 2220 2487 2221
rect 2343 2222 2344 2223
rect 2489 2222 2490 2223
rect 2357 2224 2358 2225
rect 2532 2224 2533 2225
rect 2369 2226 2370 2227
rect 2510 2226 2511 2227
rect 2372 2228 2373 2229
rect 2552 2228 2553 2229
rect 2378 2230 2379 2231
rect 2474 2230 2475 2231
rect 2382 2232 2383 2233
rect 2507 2232 2508 2233
rect 2388 2234 2389 2235
rect 2393 2234 2394 2235
rect 2399 2234 2400 2235
rect 2469 2234 2470 2235
rect 2329 2236 2330 2237
rect 2400 2236 2401 2237
rect 2439 2236 2440 2237
rect 2459 2236 2460 2237
rect 2322 2238 2323 2239
rect 2460 2238 2461 2239
rect 2445 2240 2446 2241
rect 2544 2240 2545 2241
rect 2466 2242 2467 2243
rect 2483 2242 2484 2243
rect 2475 2244 2476 2245
rect 2537 2244 2538 2245
rect 2487 2246 2488 2247
rect 2501 2246 2502 2247
rect 2493 2248 2494 2249
rect 2504 2248 2505 2249
rect 2477 2250 2478 2251
rect 2505 2250 2506 2251
rect 2495 2252 2496 2253
rect 2502 2252 2503 2253
rect 2350 2254 2351 2255
rect 2496 2254 2497 2255
rect 2511 2254 2512 2255
rect 2516 2254 2517 2255
rect 2513 2256 2514 2257
rect 2547 2256 2548 2257
rect 2514 2258 2515 2259
rect 2519 2258 2520 2259
rect 2522 2258 2523 2259
rect 2538 2258 2539 2259
rect 2523 2260 2524 2261
rect 2779 2260 2780 2261
rect 2529 2262 2530 2263
rect 2534 2262 2535 2263
rect 2535 2264 2536 2265
rect 2540 2264 2541 2265
rect 2558 2264 2559 2265
rect 2562 2264 2563 2265
rect 2555 2266 2556 2267
rect 2559 2266 2560 2267
rect 2549 2268 2550 2269
rect 2556 2268 2557 2269
rect 2565 2268 2566 2269
rect 2570 2268 2571 2269
rect 2567 2270 2568 2271
rect 2577 2270 2578 2271
rect 2568 2272 2569 2273
rect 2573 2272 2574 2273
rect 2582 2272 2583 2273
rect 2619 2272 2620 2273
rect 2588 2274 2589 2275
rect 2598 2274 2599 2275
rect 2591 2276 2592 2277
rect 2601 2276 2602 2277
rect 2592 2278 2593 2279
rect 2609 2278 2610 2279
rect 2604 2280 2605 2281
rect 2656 2280 2657 2281
rect 2623 2282 2624 2283
rect 2732 2282 2733 2283
rect 2626 2284 2627 2285
rect 2630 2284 2631 2285
rect 2629 2286 2630 2287
rect 2636 2286 2637 2287
rect 2632 2288 2633 2289
rect 2642 2288 2643 2289
rect 2639 2290 2640 2291
rect 2692 2290 2693 2291
rect 2638 2292 2639 2293
rect 2666 2292 2667 2293
rect 2641 2294 2642 2295
rect 2669 2294 2670 2295
rect 2644 2296 2645 2297
rect 2654 2296 2655 2297
rect 2672 2296 2673 2297
rect 2823 2296 2824 2297
rect 2680 2298 2681 2299
rect 2717 2298 2718 2299
rect 2606 2300 2607 2301
rect 2717 2300 2718 2301
rect 2684 2302 2685 2303
rect 2723 2302 2724 2303
rect 2683 2304 2684 2305
rect 2720 2304 2721 2305
rect 2696 2306 2697 2307
rect 2813 2306 2814 2307
rect 2698 2308 2699 2309
rect 2714 2308 2715 2309
rect 2701 2310 2702 2311
rect 2791 2310 2792 2311
rect 2704 2312 2705 2313
rect 2711 2312 2712 2313
rect 2708 2314 2709 2315
rect 2738 2314 2739 2315
rect 2707 2316 2708 2317
rect 2729 2316 2730 2317
rect 2720 2318 2721 2319
rect 2770 2318 2771 2319
rect 2726 2320 2727 2321
rect 2773 2320 2774 2321
rect 2729 2322 2730 2323
rect 2752 2322 2753 2323
rect 2732 2324 2733 2325
rect 2755 2324 2756 2325
rect 2735 2326 2736 2327
rect 2764 2326 2765 2327
rect 2744 2328 2745 2329
rect 2782 2328 2783 2329
rect 2753 2330 2754 2331
rect 2785 2330 2786 2331
rect 2756 2332 2757 2333
rect 2788 2332 2789 2333
rect 2759 2334 2760 2335
rect 2807 2334 2808 2335
rect 2762 2336 2763 2337
rect 2810 2336 2811 2337
rect 2767 2338 2768 2339
rect 2790 2338 2791 2339
rect 2797 2338 2798 2339
rect 2804 2338 2805 2339
rect 2807 2338 2808 2339
rect 2853 2338 2854 2339
rect 2810 2340 2811 2341
rect 2840 2340 2841 2341
rect 2859 2340 2860 2341
rect 2863 2340 2864 2341
rect 2866 2340 2867 2341
rect 2870 2340 2871 2341
rect 2281 2349 2282 2350
rect 2339 2349 2340 2350
rect 2288 2351 2289 2352
rect 2439 2351 2440 2352
rect 2291 2353 2292 2354
rect 2305 2353 2306 2354
rect 2290 2355 2291 2356
rect 2436 2355 2437 2356
rect 2295 2357 2296 2358
rect 2302 2357 2303 2358
rect 2312 2357 2313 2358
rect 2348 2357 2349 2358
rect 2332 2359 2333 2360
rect 2511 2359 2512 2360
rect 2345 2361 2346 2362
rect 2406 2361 2407 2362
rect 2353 2363 2354 2364
rect 2481 2363 2482 2364
rect 2382 2365 2383 2366
rect 2418 2365 2419 2366
rect 2385 2367 2386 2368
rect 2544 2367 2545 2368
rect 2388 2369 2389 2370
rect 2436 2369 2437 2370
rect 2430 2371 2431 2372
rect 2469 2371 2470 2372
rect 2445 2373 2446 2374
rect 2466 2373 2467 2374
rect 2397 2375 2398 2376
rect 2466 2375 2467 2376
rect 2448 2377 2449 2378
rect 2469 2377 2470 2378
rect 2350 2379 2351 2380
rect 2448 2379 2449 2380
rect 2457 2379 2458 2380
rect 2490 2379 2491 2380
rect 2472 2381 2473 2382
rect 2478 2381 2479 2382
rect 2472 2383 2473 2384
rect 2505 2383 2506 2384
rect 2475 2385 2476 2386
rect 2484 2385 2485 2386
rect 2502 2385 2503 2386
rect 2511 2385 2512 2386
rect 2343 2387 2344 2388
rect 2502 2387 2503 2388
rect 2342 2389 2343 2390
rect 2400 2389 2401 2390
rect 2514 2389 2515 2390
rect 2550 2389 2551 2390
rect 2517 2391 2518 2392
rect 2580 2391 2581 2392
rect 2487 2393 2488 2394
rect 2517 2393 2518 2394
rect 2523 2393 2524 2394
rect 2553 2393 2554 2394
rect 2523 2395 2524 2396
rect 2562 2395 2563 2396
rect 2538 2397 2539 2398
rect 2541 2397 2542 2398
rect 2496 2399 2497 2400
rect 2538 2399 2539 2400
rect 2556 2399 2557 2400
rect 2586 2399 2587 2400
rect 2547 2401 2548 2402
rect 2556 2401 2557 2402
rect 2336 2403 2337 2404
rect 2547 2403 2548 2404
rect 2336 2405 2337 2406
rect 2785 2405 2786 2406
rect 2559 2407 2560 2408
rect 2583 2407 2584 2408
rect 2592 2407 2593 2408
rect 2626 2407 2627 2408
rect 2595 2409 2596 2410
rect 2625 2409 2626 2410
rect 2577 2411 2578 2412
rect 2595 2411 2596 2412
rect 2598 2411 2599 2412
rect 2622 2411 2623 2412
rect 2571 2413 2572 2414
rect 2598 2413 2599 2414
rect 2535 2415 2536 2416
rect 2571 2415 2572 2416
rect 2493 2417 2494 2418
rect 2535 2417 2536 2418
rect 2460 2419 2461 2420
rect 2493 2419 2494 2420
rect 2601 2419 2602 2420
rect 2616 2419 2617 2420
rect 2565 2421 2566 2422
rect 2601 2421 2602 2422
rect 2529 2423 2530 2424
rect 2565 2423 2566 2424
rect 2499 2425 2500 2426
rect 2529 2425 2530 2426
rect 2329 2427 2330 2428
rect 2499 2427 2500 2428
rect 2604 2427 2605 2428
rect 2634 2427 2635 2428
rect 2568 2429 2569 2430
rect 2604 2429 2605 2430
rect 2532 2431 2533 2432
rect 2568 2431 2569 2432
rect 2319 2433 2320 2434
rect 2532 2433 2533 2434
rect 2619 2433 2620 2434
rect 2747 2433 2748 2434
rect 2629 2435 2630 2436
rect 2658 2435 2659 2436
rect 2638 2437 2639 2438
rect 2667 2437 2668 2438
rect 2670 2439 2671 2440
rect 2767 2439 2768 2440
rect 2676 2441 2677 2442
rect 2739 2441 2740 2442
rect 2683 2443 2684 2444
rect 2717 2443 2718 2444
rect 2701 2445 2702 2446
rect 2718 2445 2719 2446
rect 2680 2447 2681 2448
rect 2700 2447 2701 2448
rect 2644 2449 2645 2450
rect 2679 2449 2680 2450
rect 2712 2449 2713 2450
rect 2732 2449 2733 2450
rect 2698 2451 2699 2452
rect 2733 2451 2734 2452
rect 2697 2453 2698 2454
rect 2723 2453 2724 2454
rect 2720 2455 2721 2456
rect 2769 2455 2770 2456
rect 2704 2457 2705 2458
rect 2721 2457 2722 2458
rect 2632 2459 2633 2460
rect 2703 2459 2704 2460
rect 2729 2459 2730 2460
rect 2788 2459 2789 2460
rect 2730 2461 2731 2462
rect 2816 2461 2817 2462
rect 2744 2463 2745 2464
rect 2812 2463 2813 2464
rect 2753 2465 2754 2466
rect 2773 2465 2774 2466
rect 2726 2467 2727 2468
rect 2752 2467 2753 2468
rect 2756 2467 2757 2468
rect 2776 2467 2777 2468
rect 2755 2469 2756 2470
rect 2762 2469 2763 2470
rect 2759 2471 2760 2472
rect 2791 2471 2792 2472
rect 2735 2473 2736 2474
rect 2758 2473 2759 2474
rect 2736 2475 2737 2476
rect 2849 2475 2850 2476
rect 2770 2477 2771 2478
rect 2779 2477 2780 2478
rect 2807 2477 2808 2478
rect 2836 2477 2837 2478
rect 2810 2479 2811 2480
rect 2839 2479 2840 2480
rect 2287 2488 2288 2489
rect 2339 2488 2340 2489
rect 2287 2490 2288 2491
rect 2294 2490 2295 2491
rect 2297 2490 2298 2491
rect 2301 2490 2302 2491
rect 2305 2490 2306 2491
rect 2504 2490 2505 2491
rect 2322 2492 2323 2493
rect 2359 2492 2360 2493
rect 2326 2494 2327 2495
rect 2493 2494 2494 2495
rect 2312 2496 2313 2497
rect 2492 2496 2493 2497
rect 2327 2498 2328 2499
rect 2532 2498 2533 2499
rect 2330 2500 2331 2501
rect 2348 2500 2349 2501
rect 2334 2502 2335 2503
rect 2529 2502 2530 2503
rect 2345 2504 2346 2505
rect 2436 2504 2437 2505
rect 2353 2506 2354 2507
rect 2365 2506 2366 2507
rect 2406 2506 2407 2507
rect 2414 2506 2415 2507
rect 2418 2506 2419 2507
rect 2426 2506 2427 2507
rect 2430 2506 2431 2507
rect 2450 2506 2451 2507
rect 2432 2508 2433 2509
rect 2448 2508 2449 2509
rect 2475 2508 2476 2509
rect 2604 2508 2605 2509
rect 2478 2510 2479 2511
rect 2507 2510 2508 2511
rect 2484 2512 2485 2513
rect 2519 2512 2520 2513
rect 2499 2514 2500 2515
rect 2513 2514 2514 2515
rect 2517 2514 2518 2515
rect 2543 2514 2544 2515
rect 2502 2516 2503 2517
rect 2516 2516 2517 2517
rect 2490 2518 2491 2519
rect 2501 2518 2502 2519
rect 2531 2518 2532 2519
rect 2535 2518 2536 2519
rect 2534 2520 2535 2521
rect 2538 2520 2539 2521
rect 2511 2522 2512 2523
rect 2537 2522 2538 2523
rect 2481 2524 2482 2525
rect 2510 2524 2511 2525
rect 2553 2524 2554 2525
rect 2561 2524 2562 2525
rect 2565 2524 2566 2525
rect 2573 2524 2574 2525
rect 2568 2526 2569 2527
rect 2576 2526 2577 2527
rect 2547 2528 2548 2529
rect 2567 2528 2568 2529
rect 2320 2530 2321 2531
rect 2546 2530 2547 2531
rect 2571 2530 2572 2531
rect 2591 2530 2592 2531
rect 2550 2532 2551 2533
rect 2570 2532 2571 2533
rect 2541 2534 2542 2535
rect 2549 2534 2550 2535
rect 2586 2534 2587 2535
rect 2609 2534 2610 2535
rect 2454 2536 2455 2537
rect 2585 2536 2586 2537
rect 2598 2536 2599 2537
rect 2636 2536 2637 2537
rect 2384 2538 2385 2539
rect 2597 2538 2598 2539
rect 2601 2538 2602 2539
rect 2627 2538 2628 2539
rect 2556 2540 2557 2541
rect 2600 2540 2601 2541
rect 2486 2542 2487 2543
rect 2555 2542 2556 2543
rect 2612 2542 2613 2543
rect 2631 2542 2632 2543
rect 2472 2544 2473 2545
rect 2630 2544 2631 2545
rect 2469 2546 2470 2547
rect 2471 2546 2472 2547
rect 2466 2548 2467 2549
rect 2468 2548 2469 2549
rect 2619 2548 2620 2549
rect 2645 2548 2646 2549
rect 2583 2550 2584 2551
rect 2618 2550 2619 2551
rect 2625 2550 2626 2551
rect 2651 2550 2652 2551
rect 2634 2552 2635 2553
rect 2682 2552 2683 2553
rect 2595 2554 2596 2555
rect 2633 2554 2634 2555
rect 2342 2556 2343 2557
rect 2594 2556 2595 2557
rect 2658 2556 2659 2557
rect 2706 2556 2707 2557
rect 2622 2558 2623 2559
rect 2657 2558 2658 2559
rect 2670 2558 2671 2559
rect 2673 2558 2674 2559
rect 2654 2560 2655 2561
rect 2669 2560 2670 2561
rect 2676 2560 2677 2561
rect 2773 2560 2774 2561
rect 2703 2562 2704 2563
rect 2706 2562 2707 2563
rect 2700 2564 2701 2565
rect 2703 2564 2704 2565
rect 2712 2564 2713 2565
rect 2810 2564 2811 2565
rect 2715 2566 2716 2567
rect 2776 2566 2777 2567
rect 2718 2568 2719 2569
rect 2769 2568 2770 2569
rect 2679 2570 2680 2571
rect 2718 2570 2719 2571
rect 2667 2572 2668 2573
rect 2679 2572 2680 2573
rect 2721 2572 2722 2573
rect 2724 2572 2725 2573
rect 2697 2574 2698 2575
rect 2721 2574 2722 2575
rect 2697 2576 2698 2577
rect 2842 2576 2843 2577
rect 2730 2578 2731 2579
rect 2760 2578 2761 2579
rect 2733 2580 2734 2581
rect 2763 2580 2764 2581
rect 2640 2582 2641 2583
rect 2733 2582 2734 2583
rect 2616 2584 2617 2585
rect 2639 2584 2640 2585
rect 2580 2586 2581 2587
rect 2615 2586 2616 2587
rect 2736 2586 2737 2587
rect 2845 2586 2846 2587
rect 2755 2588 2756 2589
rect 2791 2588 2792 2589
rect 2758 2590 2759 2591
rect 2836 2590 2837 2591
rect 2766 2592 2767 2593
rect 2819 2592 2820 2593
rect 2788 2594 2789 2595
rect 2808 2594 2809 2595
rect 2785 2596 2786 2597
rect 2807 2596 2808 2597
rect 2752 2598 2753 2599
rect 2785 2598 2786 2599
rect 2788 2598 2789 2599
rect 2804 2598 2805 2599
rect 2839 2598 2840 2599
rect 2861 2598 2862 2599
rect 2287 2607 2288 2608
rect 2325 2607 2326 2608
rect 2301 2609 2302 2610
rect 2504 2609 2505 2610
rect 2313 2611 2314 2612
rect 2359 2611 2360 2612
rect 2320 2613 2321 2614
rect 2346 2613 2347 2614
rect 2327 2615 2328 2616
rect 2513 2615 2514 2616
rect 2328 2617 2329 2618
rect 2785 2617 2786 2618
rect 2334 2619 2335 2620
rect 2482 2619 2483 2620
rect 2337 2621 2338 2622
rect 2567 2621 2568 2622
rect 2349 2623 2350 2624
rect 2353 2623 2354 2624
rect 2352 2625 2353 2626
rect 2546 2625 2547 2626
rect 2358 2627 2359 2628
rect 2513 2627 2514 2628
rect 2361 2629 2362 2630
rect 2492 2629 2493 2630
rect 2365 2631 2366 2632
rect 2534 2631 2535 2632
rect 2375 2633 2376 2634
rect 2379 2633 2380 2634
rect 2387 2633 2388 2634
rect 2585 2633 2586 2634
rect 2414 2635 2415 2636
rect 2416 2635 2417 2636
rect 2432 2635 2433 2636
rect 2434 2635 2435 2636
rect 2438 2635 2439 2636
rect 2679 2635 2680 2636
rect 2446 2637 2447 2638
rect 2450 2637 2451 2638
rect 2449 2639 2450 2640
rect 2516 2639 2517 2640
rect 2452 2641 2453 2642
rect 2564 2641 2565 2642
rect 2458 2643 2459 2644
rect 2570 2643 2571 2644
rect 2471 2645 2472 2646
rect 2567 2645 2568 2646
rect 2479 2647 2480 2648
rect 2501 2647 2502 2648
rect 2486 2649 2487 2650
rect 2603 2649 2604 2650
rect 2488 2651 2489 2652
rect 2555 2651 2556 2652
rect 2498 2653 2499 2654
rect 2507 2653 2508 2654
rect 2501 2655 2502 2656
rect 2510 2655 2511 2656
rect 2504 2657 2505 2658
rect 2537 2657 2538 2658
rect 2510 2659 2511 2660
rect 2543 2659 2544 2660
rect 2516 2661 2517 2662
rect 2519 2661 2520 2662
rect 2522 2661 2523 2662
rect 2531 2661 2532 2662
rect 2525 2663 2526 2664
rect 2633 2663 2634 2664
rect 2426 2665 2427 2666
rect 2525 2665 2526 2666
rect 2537 2665 2538 2666
rect 2630 2665 2631 2666
rect 2540 2667 2541 2668
rect 2561 2667 2562 2668
rect 2546 2669 2547 2670
rect 2573 2669 2574 2670
rect 2552 2671 2553 2672
rect 2591 2671 2592 2672
rect 2549 2673 2550 2674
rect 2591 2673 2592 2674
rect 2549 2675 2550 2676
rect 2576 2675 2577 2676
rect 2555 2677 2556 2678
rect 2594 2677 2595 2678
rect 2558 2679 2559 2680
rect 2597 2679 2598 2680
rect 2561 2681 2562 2682
rect 2600 2681 2601 2682
rect 2582 2683 2583 2684
rect 2609 2683 2610 2684
rect 2585 2685 2586 2686
rect 2612 2685 2613 2686
rect 2588 2687 2589 2688
rect 2627 2687 2628 2688
rect 2594 2689 2595 2690
rect 2618 2689 2619 2690
rect 2600 2691 2601 2692
rect 2615 2691 2616 2692
rect 2606 2693 2607 2694
rect 2645 2693 2646 2694
rect 2612 2695 2613 2696
rect 2651 2695 2652 2696
rect 2615 2697 2616 2698
rect 2636 2697 2637 2698
rect 2618 2699 2619 2700
rect 2639 2699 2640 2700
rect 2624 2701 2625 2702
rect 2682 2701 2683 2702
rect 2633 2703 2634 2704
rect 2657 2703 2658 2704
rect 2636 2705 2637 2706
rect 2654 2705 2655 2706
rect 2665 2705 2666 2706
rect 2788 2705 2789 2706
rect 2677 2707 2678 2708
rect 2721 2707 2722 2708
rect 2680 2709 2681 2710
rect 2703 2709 2704 2710
rect 2683 2711 2684 2712
rect 2706 2711 2707 2712
rect 2694 2713 2695 2714
rect 2858 2713 2859 2714
rect 2697 2715 2698 2716
rect 2797 2715 2798 2716
rect 2698 2717 2699 2718
rect 2760 2717 2761 2718
rect 2701 2719 2702 2720
rect 2766 2719 2767 2720
rect 2704 2721 2705 2722
rect 2724 2721 2725 2722
rect 2707 2723 2708 2724
rect 2724 2723 2725 2724
rect 2715 2725 2716 2726
rect 2874 2725 2875 2726
rect 2718 2727 2719 2728
rect 2779 2727 2780 2728
rect 2730 2729 2731 2730
rect 2791 2729 2792 2730
rect 2733 2731 2734 2732
rect 2769 2731 2770 2732
rect 2733 2733 2734 2734
rect 2827 2733 2828 2734
rect 2736 2735 2737 2736
rect 2837 2735 2838 2736
rect 2742 2737 2743 2738
rect 2807 2737 2808 2738
rect 2745 2739 2746 2740
rect 2810 2739 2811 2740
rect 2763 2741 2764 2742
rect 2867 2741 2868 2742
rect 2782 2743 2783 2744
rect 2861 2743 2862 2744
rect 2296 2752 2297 2753
rect 2340 2752 2341 2753
rect 2303 2754 2304 2755
rect 2308 2754 2309 2755
rect 2312 2754 2313 2755
rect 2319 2754 2320 2755
rect 2306 2756 2307 2757
rect 2313 2756 2314 2757
rect 2319 2756 2320 2757
rect 2325 2756 2326 2757
rect 2322 2758 2323 2759
rect 2328 2758 2329 2759
rect 2328 2760 2329 2761
rect 2513 2760 2514 2761
rect 2343 2762 2344 2763
rect 2346 2762 2347 2763
rect 2349 2762 2350 2763
rect 2352 2762 2353 2763
rect 2369 2762 2370 2763
rect 2549 2762 2550 2763
rect 2375 2764 2376 2765
rect 2555 2764 2556 2765
rect 2386 2766 2387 2767
rect 2416 2766 2417 2767
rect 2415 2768 2416 2769
rect 2434 2768 2435 2769
rect 2433 2770 2434 2771
rect 2446 2770 2447 2771
rect 2436 2772 2437 2773
rect 2449 2772 2450 2773
rect 2442 2774 2443 2775
rect 2529 2774 2530 2775
rect 2458 2776 2459 2777
rect 2532 2776 2533 2777
rect 2457 2778 2458 2779
rect 2467 2778 2468 2779
rect 2460 2780 2461 2781
rect 2567 2780 2568 2781
rect 2463 2782 2464 2783
rect 2479 2782 2480 2783
rect 2466 2784 2467 2785
rect 2482 2784 2483 2785
rect 2481 2786 2482 2787
rect 2498 2786 2499 2787
rect 2484 2788 2485 2789
rect 2501 2788 2502 2789
rect 2362 2790 2363 2791
rect 2502 2790 2503 2791
rect 2493 2792 2494 2793
rect 2504 2792 2505 2793
rect 2495 2794 2496 2795
rect 2603 2794 2604 2795
rect 2499 2796 2500 2797
rect 2510 2796 2511 2797
rect 2505 2798 2506 2799
rect 2522 2798 2523 2799
rect 2508 2800 2509 2801
rect 2525 2800 2526 2801
rect 2516 2802 2517 2803
rect 2538 2802 2539 2803
rect 2517 2804 2518 2805
rect 2540 2804 2541 2805
rect 2382 2806 2383 2807
rect 2541 2806 2542 2807
rect 2523 2808 2524 2809
rect 2585 2808 2586 2809
rect 2550 2810 2551 2811
rect 2558 2810 2559 2811
rect 2564 2810 2565 2811
rect 2650 2810 2651 2811
rect 2473 2812 2474 2813
rect 2565 2812 2566 2813
rect 2574 2812 2575 2813
rect 2600 2812 2601 2813
rect 2577 2814 2578 2815
rect 2588 2814 2589 2815
rect 2534 2816 2535 2817
rect 2589 2816 2590 2817
rect 2535 2818 2536 2819
rect 2546 2818 2547 2819
rect 2547 2820 2548 2821
rect 2552 2820 2553 2821
rect 2553 2822 2554 2823
rect 2561 2822 2562 2823
rect 2562 2824 2563 2825
rect 2582 2824 2583 2825
rect 2580 2826 2581 2827
rect 2591 2826 2592 2827
rect 2594 2826 2595 2827
rect 2642 2826 2643 2827
rect 2595 2828 2596 2829
rect 2606 2828 2607 2829
rect 2592 2830 2593 2831
rect 2607 2830 2608 2831
rect 2601 2832 2602 2833
rect 2612 2832 2613 2833
rect 2604 2834 2605 2835
rect 2615 2834 2616 2835
rect 2610 2836 2611 2837
rect 2624 2836 2625 2837
rect 2613 2838 2614 2839
rect 2618 2838 2619 2839
rect 2625 2838 2626 2839
rect 2633 2838 2634 2839
rect 2628 2840 2629 2841
rect 2636 2840 2637 2841
rect 2637 2842 2638 2843
rect 2683 2842 2684 2843
rect 2643 2844 2644 2845
rect 2646 2844 2647 2845
rect 2668 2844 2669 2845
rect 2727 2844 2728 2845
rect 2668 2846 2669 2847
rect 2677 2846 2678 2847
rect 2686 2846 2687 2847
rect 2698 2846 2699 2847
rect 2689 2848 2690 2849
rect 2704 2848 2705 2849
rect 2661 2850 2662 2851
rect 2704 2850 2705 2851
rect 2701 2852 2702 2853
rect 2717 2852 2718 2853
rect 2701 2854 2702 2855
rect 2736 2854 2737 2855
rect 2707 2856 2708 2857
rect 2710 2856 2711 2857
rect 2680 2858 2681 2859
rect 2707 2858 2708 2859
rect 2713 2858 2714 2859
rect 2720 2858 2721 2859
rect 2730 2858 2731 2859
rect 2739 2858 2740 2859
rect 2736 2860 2737 2861
rect 2758 2860 2759 2861
rect 2742 2862 2743 2863
rect 2751 2862 2752 2863
rect 2727 2864 2728 2865
rect 2742 2864 2743 2865
rect 2745 2864 2746 2865
rect 2754 2864 2755 2865
rect 2723 2866 2724 2867
rect 2745 2866 2746 2867
rect 2782 2866 2783 2867
rect 2791 2866 2792 2867
rect 2683 2868 2684 2869
rect 2781 2868 2782 2869
rect 2300 2877 2301 2878
rect 2340 2877 2341 2878
rect 2296 2879 2297 2880
rect 2300 2879 2301 2880
rect 2309 2879 2310 2880
rect 2399 2879 2400 2880
rect 2313 2881 2314 2882
rect 2387 2881 2388 2882
rect 2319 2883 2320 2884
rect 2383 2883 2384 2884
rect 2296 2885 2297 2886
rect 2384 2885 2385 2886
rect 2321 2887 2322 2888
rect 2499 2887 2500 2888
rect 2324 2889 2325 2890
rect 2493 2889 2494 2890
rect 2328 2891 2329 2892
rect 2333 2891 2334 2892
rect 2343 2891 2344 2892
rect 2345 2891 2346 2892
rect 2349 2891 2350 2892
rect 2351 2891 2352 2892
rect 2358 2891 2359 2892
rect 2436 2891 2437 2892
rect 2357 2893 2358 2894
rect 2514 2893 2515 2894
rect 2376 2895 2377 2896
rect 2601 2895 2602 2896
rect 2390 2897 2391 2898
rect 2502 2897 2503 2898
rect 2367 2899 2368 2900
rect 2502 2899 2503 2900
rect 2405 2901 2406 2902
rect 2559 2901 2560 2902
rect 2439 2903 2440 2904
rect 2565 2903 2566 2904
rect 2415 2905 2416 2906
rect 2439 2905 2440 2906
rect 2457 2905 2458 2906
rect 2475 2905 2476 2906
rect 2460 2907 2461 2908
rect 2469 2907 2470 2908
rect 2478 2907 2479 2908
rect 2481 2907 2482 2908
rect 2481 2909 2482 2910
rect 2484 2909 2485 2910
rect 2490 2909 2491 2910
rect 2505 2909 2506 2910
rect 2493 2911 2494 2912
rect 2508 2911 2509 2912
rect 2508 2913 2509 2914
rect 2517 2913 2518 2914
rect 2355 2915 2356 2916
rect 2517 2915 2518 2916
rect 2523 2915 2524 2916
rect 2568 2915 2569 2916
rect 2526 2917 2527 2918
rect 2535 2917 2536 2918
rect 2532 2919 2533 2920
rect 2535 2919 2536 2920
rect 2529 2921 2530 2922
rect 2532 2921 2533 2922
rect 2544 2921 2545 2922
rect 2550 2921 2551 2922
rect 2547 2923 2548 2924
rect 2550 2923 2551 2924
rect 2547 2925 2548 2926
rect 2553 2925 2554 2926
rect 2562 2925 2563 2926
rect 2565 2925 2566 2926
rect 2538 2927 2539 2928
rect 2562 2927 2563 2928
rect 2538 2929 2539 2930
rect 2541 2929 2542 2930
rect 2580 2929 2581 2930
rect 2583 2929 2584 2930
rect 2577 2931 2578 2932
rect 2580 2931 2581 2932
rect 2574 2933 2575 2934
rect 2577 2933 2578 2934
rect 2592 2933 2593 2934
rect 2791 2933 2792 2934
rect 2595 2935 2596 2936
rect 2622 2935 2623 2936
rect 2607 2937 2608 2938
rect 2616 2937 2617 2938
rect 2613 2939 2614 2940
rect 2619 2939 2620 2940
rect 2604 2941 2605 2942
rect 2613 2941 2614 2942
rect 2631 2941 2632 2942
rect 2646 2941 2647 2942
rect 2634 2943 2635 2944
rect 2713 2943 2714 2944
rect 2637 2945 2638 2946
rect 2646 2945 2647 2946
rect 2637 2947 2638 2948
rect 2698 2947 2699 2948
rect 2668 2949 2669 2950
rect 2671 2949 2672 2950
rect 2683 2949 2684 2950
rect 2762 2949 2763 2950
rect 2689 2951 2690 2952
rect 2695 2951 2696 2952
rect 2689 2953 2690 2954
rect 2769 2953 2770 2954
rect 2692 2955 2693 2956
rect 2765 2955 2766 2956
rect 2710 2957 2711 2958
rect 2720 2957 2721 2958
rect 2658 2959 2659 2960
rect 2710 2959 2711 2960
rect 2730 2959 2731 2960
rect 2733 2959 2734 2960
rect 2733 2961 2734 2962
rect 2736 2961 2737 2962
rect 2628 2963 2629 2964
rect 2736 2963 2737 2964
rect 2625 2965 2626 2966
rect 2628 2965 2629 2966
rect 2739 2965 2740 2966
rect 2760 2965 2761 2966
rect 2742 2967 2743 2968
rect 2748 2967 2749 2968
rect 2751 2967 2752 2968
rect 2756 2967 2757 2968
rect 2754 2969 2755 2970
rect 2759 2969 2760 2970
rect 2296 2978 2297 2979
rect 2300 2978 2301 2979
rect 2299 2980 2300 2981
rect 2466 2980 2467 2981
rect 2307 2982 2308 2983
rect 2384 2982 2385 2983
rect 2314 2984 2315 2985
rect 2345 2984 2346 2985
rect 2320 2986 2321 2987
rect 2333 2986 2334 2987
rect 2329 2988 2330 2989
rect 2517 2988 2518 2989
rect 2349 2990 2350 2991
rect 2387 2990 2388 2991
rect 2351 2992 2352 2993
rect 2409 2992 2410 2993
rect 2352 2994 2353 2995
rect 2390 2994 2391 2995
rect 2355 2996 2356 2997
rect 2550 2996 2551 2997
rect 2357 2998 2358 2999
rect 2371 2998 2372 2999
rect 2358 3000 2359 3001
rect 2451 3000 2452 3001
rect 2360 3002 2361 3003
rect 2399 3002 2400 3003
rect 2381 3004 2382 3005
rect 2514 3004 2515 3005
rect 2381 3006 2382 3007
rect 2433 3006 2434 3007
rect 2384 3008 2385 3009
rect 2439 3008 2440 3009
rect 2396 3010 2397 3011
rect 2538 3010 2539 3011
rect 2409 3012 2410 3013
rect 2469 3012 2470 3013
rect 2412 3014 2413 3015
rect 2547 3014 2548 3015
rect 2424 3016 2425 3017
rect 2478 3016 2479 3017
rect 2365 3018 2366 3019
rect 2478 3018 2479 3019
rect 2430 3020 2431 3021
rect 2490 3020 2491 3021
rect 2433 3022 2434 3023
rect 2472 3022 2473 3023
rect 2445 3024 2446 3025
rect 2502 3024 2503 3025
rect 2402 3026 2403 3027
rect 2502 3026 2503 3027
rect 2403 3028 2404 3029
rect 2493 3028 2494 3029
rect 2460 3030 2461 3031
rect 2526 3030 2527 3031
rect 2484 3032 2485 3033
rect 2532 3032 2533 3033
rect 2487 3034 2488 3035
rect 2535 3034 2536 3035
rect 2490 3036 2491 3037
rect 2544 3036 2545 3037
rect 2493 3038 2494 3039
rect 2508 3038 2509 3039
rect 2508 3040 2509 3041
rect 2559 3040 2560 3041
rect 2511 3042 2512 3043
rect 2562 3042 2563 3043
rect 2514 3044 2515 3045
rect 2565 3044 2566 3045
rect 2517 3046 2518 3047
rect 2568 3046 2569 3047
rect 2526 3048 2527 3049
rect 2577 3048 2578 3049
rect 2529 3050 2530 3051
rect 2580 3050 2581 3051
rect 2532 3052 2533 3053
rect 2583 3052 2584 3053
rect 2541 3054 2542 3055
rect 2613 3054 2614 3055
rect 2544 3056 2545 3057
rect 2616 3056 2617 3057
rect 2559 3058 2560 3059
rect 2610 3058 2611 3059
rect 2562 3060 2563 3061
rect 2619 3060 2620 3061
rect 2565 3062 2566 3063
rect 2622 3062 2623 3063
rect 2568 3064 2569 3065
rect 2631 3064 2632 3065
rect 2577 3066 2578 3067
rect 2637 3066 2638 3067
rect 2586 3068 2587 3069
rect 2646 3068 2647 3069
rect 2610 3070 2611 3071
rect 2671 3070 2672 3071
rect 2613 3072 2614 3073
rect 2695 3072 2696 3073
rect 2622 3074 2623 3075
rect 2689 3074 2690 3075
rect 2625 3076 2626 3077
rect 2686 3076 2687 3077
rect 2628 3078 2629 3079
rect 2692 3078 2693 3079
rect 2631 3080 2632 3081
rect 2650 3080 2651 3081
rect 2634 3082 2635 3083
rect 2643 3082 2644 3083
rect 2463 3084 2464 3085
rect 2634 3084 2635 3085
rect 2637 3084 2638 3085
rect 2704 3084 2705 3085
rect 2640 3086 2641 3087
rect 2707 3086 2708 3087
rect 2661 3088 2662 3089
rect 2665 3088 2666 3089
rect 2663 3090 2664 3091
rect 2730 3090 2731 3091
rect 2666 3092 2667 3093
rect 2733 3092 2734 3093
rect 2689 3094 2690 3095
rect 2756 3094 2757 3095
rect 2692 3096 2693 3097
rect 2759 3096 2760 3097
rect 2698 3098 2699 3099
rect 2772 3098 2773 3099
rect 2299 3107 2300 3108
rect 2312 3107 2313 3108
rect 2306 3109 2307 3110
rect 2315 3109 2316 3110
rect 2317 3109 2318 3110
rect 2352 3109 2353 3110
rect 2329 3111 2330 3112
rect 2349 3111 2350 3112
rect 2332 3113 2333 3114
rect 2440 3113 2441 3114
rect 2336 3115 2337 3116
rect 2396 3115 2397 3116
rect 2343 3117 2344 3118
rect 2511 3117 2512 3118
rect 2356 3119 2357 3120
rect 2451 3119 2452 3120
rect 2362 3121 2363 3122
rect 2472 3121 2473 3122
rect 2372 3123 2373 3124
rect 2384 3123 2385 3124
rect 2381 3125 2382 3126
rect 2443 3125 2444 3126
rect 2406 3127 2407 3128
rect 2409 3127 2410 3128
rect 2419 3127 2420 3128
rect 2424 3127 2425 3128
rect 2425 3129 2426 3130
rect 2430 3129 2431 3130
rect 2434 3129 2435 3130
rect 2445 3129 2446 3130
rect 2470 3129 2471 3130
rect 2478 3129 2479 3130
rect 2473 3131 2474 3132
rect 2481 3131 2482 3132
rect 2476 3133 2477 3134
rect 2484 3133 2485 3134
rect 2479 3135 2480 3136
rect 2487 3135 2488 3136
rect 2482 3137 2483 3138
rect 2490 3137 2491 3138
rect 2485 3139 2486 3140
rect 2493 3139 2494 3140
rect 2494 3141 2495 3142
rect 2502 3141 2503 3142
rect 2460 3143 2461 3144
rect 2503 3143 2504 3144
rect 2500 3145 2501 3146
rect 2508 3145 2509 3146
rect 2506 3147 2507 3148
rect 2514 3147 2515 3148
rect 2509 3149 2510 3150
rect 2517 3149 2518 3150
rect 2512 3151 2513 3152
rect 2532 3151 2533 3152
rect 2518 3153 2519 3154
rect 2526 3153 2527 3154
rect 2521 3155 2522 3156
rect 2529 3155 2530 3156
rect 2544 3155 2545 3156
rect 2548 3155 2549 3156
rect 2541 3157 2542 3158
rect 2545 3157 2546 3158
rect 2557 3157 2558 3158
rect 2574 3157 2575 3158
rect 2568 3159 2569 3160
rect 2581 3159 2582 3160
rect 2562 3161 2563 3162
rect 2569 3161 2570 3162
rect 2523 3163 2524 3164
rect 2563 3163 2564 3164
rect 2466 3165 2467 3166
rect 2524 3165 2525 3166
rect 2577 3165 2578 3166
rect 2584 3165 2585 3166
rect 2610 3165 2611 3166
rect 2617 3165 2618 3166
rect 2613 3167 2614 3168
rect 2644 3167 2645 3168
rect 2614 3169 2615 3170
rect 2705 3169 2706 3170
rect 2620 3171 2621 3172
rect 2692 3171 2693 3172
rect 2622 3173 2623 3174
rect 2703 3173 2704 3174
rect 2637 3175 2638 3176
rect 2646 3175 2647 3176
rect 2638 3177 2639 3178
rect 2640 3177 2641 3178
rect 2586 3179 2587 3180
rect 2641 3179 2642 3180
rect 2587 3181 2588 3182
rect 2632 3181 2633 3182
rect 2663 3181 2664 3182
rect 2681 3181 2682 3182
rect 2666 3183 2667 3184
rect 2684 3183 2685 3184
rect 2689 3183 2690 3184
rect 2730 3183 2731 3184
rect 2628 3185 2629 3186
rect 2690 3185 2691 3186
rect 2625 3187 2626 3188
rect 2629 3187 2630 3188
rect 2700 3187 2701 3188
rect 2727 3187 2728 3188
rect 2299 3196 2300 3197
rect 2306 3196 2307 3197
rect 2302 3198 2303 3199
rect 2312 3198 2313 3199
rect 2312 3200 2313 3201
rect 2325 3200 2326 3201
rect 2306 3202 2307 3203
rect 2325 3202 2326 3203
rect 2315 3204 2316 3205
rect 2318 3204 2319 3205
rect 2315 3206 2316 3207
rect 2396 3206 2397 3207
rect 2322 3208 2323 3209
rect 2440 3208 2441 3209
rect 2332 3210 2333 3211
rect 2482 3210 2483 3211
rect 2335 3212 2336 3213
rect 2425 3212 2426 3213
rect 2339 3214 2340 3215
rect 2494 3214 2495 3215
rect 2356 3216 2357 3217
rect 2387 3216 2388 3217
rect 2359 3218 2360 3219
rect 2383 3218 2384 3219
rect 2368 3220 2369 3221
rect 2372 3220 2373 3221
rect 2380 3220 2381 3221
rect 2443 3220 2444 3221
rect 2404 3222 2405 3223
rect 2409 3222 2410 3223
rect 2417 3222 2418 3223
rect 2490 3222 2491 3223
rect 2419 3224 2420 3225
rect 2736 3224 2737 3225
rect 2439 3226 2440 3227
rect 2485 3226 2486 3227
rect 2448 3228 2449 3229
rect 2512 3228 2513 3229
rect 2460 3230 2461 3231
rect 2476 3230 2477 3231
rect 2463 3232 2464 3233
rect 2479 3232 2480 3233
rect 2466 3234 2467 3235
rect 2470 3234 2471 3235
rect 2469 3236 2470 3237
rect 2473 3236 2474 3237
rect 2472 3238 2473 3239
rect 2506 3238 2507 3239
rect 2484 3240 2485 3241
rect 2500 3240 2501 3241
rect 2487 3242 2488 3243
rect 2503 3242 2504 3243
rect 2493 3244 2494 3245
rect 2509 3244 2510 3245
rect 2496 3246 2497 3247
rect 2518 3246 2519 3247
rect 2505 3248 2506 3249
rect 2521 3248 2522 3249
rect 2424 3250 2425 3251
rect 2520 3250 2521 3251
rect 2508 3252 2509 3253
rect 2524 3252 2525 3253
rect 2511 3254 2512 3255
rect 2548 3254 2549 3255
rect 2514 3256 2515 3257
rect 2545 3256 2546 3257
rect 2523 3258 2524 3259
rect 2566 3258 2567 3259
rect 2526 3260 2527 3261
rect 2581 3260 2582 3261
rect 2529 3262 2530 3263
rect 2560 3262 2561 3263
rect 2539 3264 2540 3265
rect 2557 3264 2558 3265
rect 2542 3266 2543 3267
rect 2654 3266 2655 3267
rect 2558 3268 2559 3269
rect 2638 3268 2639 3269
rect 2561 3270 2562 3271
rect 2641 3270 2642 3271
rect 2563 3272 2564 3273
rect 2572 3272 2573 3273
rect 2564 3274 2565 3275
rect 2644 3274 2645 3275
rect 2569 3276 2570 3277
rect 2608 3276 2609 3277
rect 2573 3278 2574 3279
rect 2587 3278 2588 3279
rect 2584 3280 2585 3281
rect 2664 3280 2665 3281
rect 2600 3282 2601 3283
rect 2620 3282 2621 3283
rect 2609 3284 2610 3285
rect 2678 3284 2679 3285
rect 2612 3286 2613 3287
rect 2617 3286 2618 3287
rect 2614 3288 2615 3289
rect 2671 3288 2672 3289
rect 2615 3290 2616 3291
rect 2635 3290 2636 3291
rect 2618 3292 2619 3293
rect 2624 3292 2625 3293
rect 2627 3292 2628 3293
rect 2681 3292 2682 3293
rect 2629 3294 2630 3295
rect 2697 3294 2698 3295
rect 2630 3296 2631 3297
rect 2684 3296 2685 3297
rect 2646 3298 2647 3299
rect 2690 3298 2691 3299
rect 2649 3300 2650 3301
rect 2703 3300 2704 3301
rect 2676 3302 2677 3303
rect 2700 3302 2701 3303
rect 2700 3304 2701 3305
rect 2707 3304 2708 3305
rect 2309 3313 2310 3314
rect 2315 3313 2316 3314
rect 2319 3313 2320 3314
rect 2496 3313 2497 3314
rect 2321 3315 2322 3316
rect 2325 3315 2326 3316
rect 2335 3315 2336 3316
rect 2484 3315 2485 3316
rect 2368 3317 2369 3318
rect 2377 3317 2378 3318
rect 2380 3317 2381 3318
rect 2389 3317 2390 3318
rect 2383 3319 2384 3320
rect 2392 3319 2393 3320
rect 2398 3319 2399 3320
rect 2410 3319 2411 3320
rect 2402 3321 2403 3322
rect 2649 3321 2650 3322
rect 2407 3323 2408 3324
rect 2424 3323 2425 3324
rect 2404 3325 2405 3326
rect 2408 3325 2409 3326
rect 2414 3325 2415 3326
rect 2472 3325 2473 3326
rect 2417 3327 2418 3328
rect 2505 3327 2506 3328
rect 2424 3329 2425 3330
rect 2433 3329 2434 3330
rect 2436 3329 2437 3330
rect 2460 3329 2461 3330
rect 2451 3331 2452 3332
rect 2466 3331 2467 3332
rect 2454 3333 2455 3334
rect 2469 3333 2470 3334
rect 2463 3335 2464 3336
rect 2716 3335 2717 3336
rect 2448 3337 2449 3338
rect 2463 3337 2464 3338
rect 2439 3339 2440 3340
rect 2448 3339 2449 3340
rect 2290 3341 2291 3342
rect 2439 3341 2440 3342
rect 2466 3341 2467 3342
rect 2508 3341 2509 3342
rect 2475 3343 2476 3344
rect 2490 3343 2491 3344
rect 2478 3345 2479 3346
rect 2493 3345 2494 3346
rect 2487 3347 2488 3348
rect 2634 3347 2635 3348
rect 2493 3349 2494 3350
rect 2511 3349 2512 3350
rect 2487 3351 2488 3352
rect 2512 3351 2513 3352
rect 2496 3353 2497 3354
rect 2514 3353 2515 3354
rect 2499 3355 2500 3356
rect 2523 3355 2524 3356
rect 2515 3357 2516 3358
rect 2529 3357 2530 3358
rect 2517 3359 2518 3360
rect 2539 3359 2540 3360
rect 2518 3361 2519 3362
rect 2526 3361 2527 3362
rect 2538 3361 2539 3362
rect 2561 3361 2562 3362
rect 2544 3363 2545 3364
rect 2558 3363 2559 3364
rect 2547 3365 2548 3366
rect 2564 3365 2565 3366
rect 2559 3367 2560 3368
rect 2612 3367 2613 3368
rect 2568 3369 2569 3370
rect 2624 3369 2625 3370
rect 2571 3371 2572 3372
rect 2618 3371 2619 3372
rect 2573 3373 2574 3374
rect 2591 3373 2592 3374
rect 2553 3375 2554 3376
rect 2574 3375 2575 3376
rect 2584 3375 2585 3376
rect 2600 3375 2601 3376
rect 2587 3377 2588 3378
rect 2627 3377 2628 3378
rect 2609 3379 2610 3380
rect 2652 3379 2653 3380
rect 2615 3381 2616 3382
rect 2621 3381 2622 3382
rect 2630 3381 2631 3382
rect 2662 3381 2663 3382
rect 2637 3383 2638 3384
rect 2683 3383 2684 3384
rect 2646 3385 2647 3386
rect 2673 3385 2674 3386
rect 2655 3387 2656 3388
rect 2687 3387 2688 3388
rect 2696 3387 2697 3388
rect 2700 3387 2701 3388
rect 2311 3396 2312 3397
rect 2318 3396 2319 3397
rect 2320 3396 2321 3397
rect 2332 3396 2333 3397
rect 2328 3398 2329 3399
rect 2424 3398 2425 3399
rect 2331 3400 2332 3401
rect 2345 3400 2346 3401
rect 2335 3402 2336 3403
rect 2436 3402 2437 3403
rect 2334 3404 2335 3405
rect 2439 3404 2440 3405
rect 2371 3406 2372 3407
rect 2389 3406 2390 3407
rect 2374 3408 2375 3409
rect 2392 3408 2393 3409
rect 2377 3410 2378 3411
rect 2383 3410 2384 3411
rect 2392 3410 2393 3411
rect 2408 3410 2409 3411
rect 2398 3412 2399 3413
rect 2475 3412 2476 3413
rect 2402 3414 2403 3415
rect 2463 3414 2464 3415
rect 2408 3416 2409 3417
rect 2512 3416 2513 3417
rect 2411 3418 2412 3419
rect 2448 3418 2449 3419
rect 2414 3420 2415 3421
rect 2478 3420 2479 3421
rect 2418 3422 2419 3423
rect 2466 3422 2467 3423
rect 2420 3424 2421 3425
rect 2451 3424 2452 3425
rect 2430 3426 2431 3427
rect 2454 3426 2455 3427
rect 2436 3428 2437 3429
rect 2487 3428 2488 3429
rect 2442 3430 2443 3431
rect 2493 3430 2494 3431
rect 2445 3432 2446 3433
rect 2496 3432 2497 3433
rect 2495 3434 2496 3435
rect 2568 3434 2569 3435
rect 2499 3436 2500 3437
rect 2502 3436 2503 3437
rect 2498 3438 2499 3439
rect 2571 3438 2572 3439
rect 2501 3440 2502 3441
rect 2547 3440 2548 3441
rect 2504 3442 2505 3443
rect 2553 3442 2554 3443
rect 2507 3444 2508 3445
rect 2559 3444 2560 3445
rect 2515 3446 2516 3447
rect 2528 3446 2529 3447
rect 2522 3448 2523 3449
rect 2587 3448 2588 3449
rect 2525 3450 2526 3451
rect 2604 3450 2605 3451
rect 2538 3452 2539 3453
rect 2634 3452 2635 3453
rect 2541 3454 2542 3455
rect 2618 3454 2619 3455
rect 2571 3456 2572 3457
rect 2637 3456 2638 3457
rect 2287 3465 2288 3466
rect 2462 3465 2463 3466
rect 2324 3467 2325 3468
rect 2445 3467 2446 3468
rect 2356 3469 2357 3470
rect 2371 3469 2372 3470
rect 2359 3471 2360 3472
rect 2374 3471 2375 3472
rect 2379 3471 2380 3472
rect 2411 3471 2412 3472
rect 2383 3473 2384 3474
rect 2390 3473 2391 3474
rect 2392 3473 2393 3474
rect 2535 3473 2536 3474
rect 2403 3475 2404 3476
rect 2414 3475 2415 3476
rect 2406 3477 2407 3478
rect 2408 3477 2409 3478
rect 2415 3477 2416 3478
rect 2448 3477 2449 3478
rect 2421 3479 2422 3480
rect 2436 3479 2437 3480
rect 2424 3481 2425 3482
rect 2442 3481 2443 3482
rect 2474 3481 2475 3482
rect 2495 3481 2496 3482
rect 2477 3483 2478 3484
rect 2498 3483 2499 3484
rect 2486 3485 2487 3486
rect 2507 3485 2508 3486
rect 2501 3487 2502 3488
rect 2522 3487 2523 3488
rect 2504 3489 2505 3490
rect 2516 3489 2517 3490
rect 2504 3491 2505 3492
rect 2525 3491 2526 3492
rect 2520 3493 2521 3494
rect 2541 3493 2542 3494
rect 2523 3495 2524 3496
rect 2544 3495 2545 3496
rect 2550 3495 2551 3496
rect 2571 3495 2572 3496
rect 2577 3495 2578 3496
rect 2584 3495 2585 3496
rect 2323 3504 2324 3505
rect 2359 3504 2360 3505
rect 2356 3506 2357 3507
rect 2388 3506 2389 3507
rect 2391 3506 2392 3507
rect 2406 3506 2407 3507
rect 2393 3508 2394 3509
rect 2403 3508 2404 3509
rect 2406 3508 2407 3509
rect 2427 3508 2428 3509
rect 2409 3510 2410 3511
rect 2415 3510 2416 3511
rect 2418 3510 2419 3511
rect 2424 3510 2425 3511
rect 2441 3510 2442 3511
rect 2520 3510 2521 3511
rect 2468 3512 2469 3513
rect 2474 3512 2475 3513
rect 2471 3514 2472 3515
rect 2477 3514 2478 3515
rect 2480 3514 2481 3515
rect 2486 3514 2487 3515
rect 2495 3514 2496 3515
rect 2523 3514 2524 3515
rect 2498 3516 2499 3517
rect 2501 3516 2502 3517
rect 2504 3516 2505 3517
rect 2518 3516 2519 3517
rect 2550 3516 2551 3517
rect 2556 3516 2557 3517
rect 2563 3516 2564 3517
rect 2570 3516 2571 3517
rect 2383 3525 2384 3526
rect 2391 3525 2392 3526
rect 2388 3527 2389 3528
rect 2480 3527 2481 3528
rect 2392 3529 2393 3530
rect 2418 3529 2419 3530
rect 2394 3531 2395 3532
rect 2406 3531 2407 3532
rect 2397 3533 2398 3534
rect 2409 3533 2410 3534
rect 2431 3533 2432 3534
rect 2468 3533 2469 3534
rect 2437 3535 2438 3536
rect 2471 3535 2472 3536
rect 2454 3537 2455 3538
rect 2498 3537 2499 3538
rect 2495 3539 2496 3540
rect 2518 3539 2519 3540
rect 2377 3548 2378 3549
rect 2383 3548 2384 3549
rect 2389 3548 2390 3549
rect 2392 3548 2393 3549
rect 2395 3548 2396 3549
rect 2454 3548 2455 3549
rect 2409 3550 2410 3551
rect 2431 3550 2432 3551
rect 2441 3550 2442 3551
rect 2448 3550 2449 3551
<< end >>
