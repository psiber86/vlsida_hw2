magic
tech scmos
timestamp 1395743083
<< m1p >>
use CELL  1
transform -1 0 2078 0 1 2250
box 0 0 6 6
use CELL  2
transform -1 0 2151 0 1 3547
box 0 0 6 6
use CELL  3
transform -1 0 2370 0 1 5273
box 0 0 6 6
use CELL  4
transform 1 0 2128 0 -1 1392
box 0 0 6 6
use CELL  5
transform -1 0 2100 0 1 1138
box 0 0 6 6
use CELL  6
transform -1 0 2156 0 1 5755
box 0 0 6 6
use CELL  7
transform -1 0 2110 0 -1 1059
box 0 0 6 6
use CELL  8
transform -1 0 2792 0 1 2013
box 0 0 6 6
use CELL  9
transform -1 0 2134 0 1 5668
box 0 0 6 6
use CELL  10
transform -1 0 2724 0 -1 3802
box 0 0 6 6
use CELL  11
transform -1 0 2169 0 1 4897
box 0 0 6 6
use CELL  12
transform -1 0 2104 0 1 5273
box 0 0 6 6
use CELL  13
transform -1 0 2183 0 1 2013
box 0 0 6 6
use CELL  14
transform -1 0 2061 0 -1 2517
box 0 0 6 6
use CELL  15
transform -1 0 2066 0 1 1760
box 0 0 6 6
use CELL  16
transform -1 0 2099 0 1 4240
box 0 0 6 6
use CELL  17
transform -1 0 2584 0 -1 1392
box 0 0 6 6
use CELL  18
transform -1 0 2827 0 -1 3553
box 0 0 6 6
use CELL  19
transform -1 0 2720 0 1 2013
box 0 0 6 6
use CELL  20
transform -1 0 2725 0 1 4897
box 0 0 6 6
use CELL  21
transform 1 0 2685 0 1 4704
box 0 0 6 6
use CELL  22
transform -1 0 2742 0 -1 3802
box 0 0 6 6
use CELL  23
transform -1 0 2113 0 1 5668
box 0 0 6 6
use CELL  24
transform 1 0 2408 0 -1 1144
box 0 0 6 6
use CELL  25
transform 1 0 2710 0 1 1573
box 0 0 6 6
use CELL  26
transform -1 0 2134 0 1 2013
box 0 0 6 6
use CELL  27
transform -1 0 2159 0 1 2511
box 0 0 6 6
use CELL  28
transform -1 0 2718 0 1 4021
box 0 0 6 6
use CELL  29
transform -1 0 2552 0 1 4704
box 0 0 6 6
use CELL  30
transform -1 0 2266 0 1 1053
box 0 0 6 6
use CELL  31
transform -1 0 2096 0 1 3796
box 0 0 6 6
use CELL  32
transform -1 0 2813 0 1 2013
box 0 0 6 6
use CELL  33
transform -1 0 2083 0 1 5273
box 0 0 6 6
use CELL  34
transform -1 0 2146 0 1 5668
box 0 0 6 6
use CELL  35
transform -1 0 2162 0 1 4240
box 0 0 6 6
use CELL  36
transform -1 0 2082 0 1 2511
box 0 0 6 6
use CELL  37
transform -1 0 2612 0 -1 1392
box 0 0 6 6
use CELL  38
transform -1 0 2785 0 1 2250
box 0 0 6 6
use CELL  39
transform -1 0 2692 0 1 4897
box 0 0 6 6
use CELL  40
transform -1 0 2145 0 1 1573
box 0 0 6 6
use CELL  41
transform -1 0 2606 0 1 4704
box 0 0 6 6
use CELL  42
transform 1 0 2779 0 1 4240
box 0 0 6 6
use CELL  43
transform -1 0 2241 0 1 1053
box 0 0 6 6
use CELL  44
transform 1 0 2046 0 -1 5424
box 0 0 6 6
use CELL  45
transform -1 0 2260 0 1 2800
box 0 0 6 6
use CELL  46
transform 1 0 2090 0 -1 1766
box 0 0 6 6
use CELL  47
transform -1 0 2119 0 1 3322
box 0 0 6 6
use CELL  48
transform -1 0 2753 0 1 3085
box 0 0 6 6
use CELL  49
transform -1 0 2224 0 1 2250
box 0 0 6 6
use CELL  50
transform -1 0 2059 0 1 1760
box 0 0 6 6
use CELL  51
transform -1 0 2130 0 1 5273
box 0 0 6 6
use CELL  52
transform 1 0 2100 0 -1 4246
box 0 0 6 6
use CELL  53
transform -1 0 2144 0 1 4704
box 0 0 6 6
use CELL  54
transform -1 0 2079 0 1 4704
box 0 0 6 6
use CELL  55
transform -1 0 2502 0 1 5418
box 0 0 6 6
use CELL  56
transform 1 0 2718 0 -1 4710
box 0 0 6 6
use CELL  57
transform -1 0 2112 0 -1 3328
box 0 0 6 6
use CELL  58
transform -1 0 2699 0 -1 4903
box 0 0 6 6
use CELL  59
transform -1 0 2432 0 1 5418
box 0 0 6 6
use CELL  60
transform -1 0 2660 0 1 4897
box 0 0 6 6
use CELL  61
transform -1 0 2751 0 1 4021
box 0 0 6 6
use CELL  62
transform -1 0 2150 0 1 5418
box 0 0 6 6
use CELL  63
transform 1 0 2048 0 1 3796
box 0 0 6 6
use CELL  64
transform -1 0 2144 0 -1 4469
box 0 0 6 6
use CELL  65
transform -1 0 2264 0 1 5755
box 0 0 6 6
use CELL  66
transform 1 0 2065 0 1 4240
box 0 0 6 6
use CELL  67
transform -1 0 2192 0 1 5755
box 0 0 6 6
use CELL  68
transform -1 0 2591 0 1 1386
box 0 0 6 6
use CELL  69
transform -1 0 2926 0 1 2250
box 0 0 6 6
use CELL  70
transform -1 0 2768 0 -1 3328
box 0 0 6 6
use CELL  71
transform -1 0 2172 0 1 5100
box 0 0 6 6
use CELL  72
transform -1 0 2729 0 1 4240
box 0 0 6 6
use CELL  73
transform -1 0 2164 0 1 5668
box 0 0 6 6
use CELL  74
transform 1 0 2065 0 -1 1259
box 0 0 6 6
use CELL  75
transform -1 0 2130 0 1 1760
box 0 0 6 6
use CELL  76
transform -1 0 2768 0 1 4463
box 0 0 6 6
use CELL  77
transform -1 0 2137 0 1 4463
box 0 0 6 6
use CELL  78
transform -1 0 2127 0 1 2250
box 0 0 6 6
use CELL  79
transform -1 0 2176 0 1 3547
box 0 0 6 6
use CELL  80
transform 1 0 2062 0 -1 3802
box 0 0 6 6
use CELL  81
transform 1 0 2041 0 -1 3802
box 0 0 6 6
use CELL  82
transform 1 0 2793 0 -1 3802
box 0 0 6 6
use CELL  83
transform -1 0 2311 0 1 4897
box 0 0 6 6
use CELL  84
transform -1 0 2743 0 1 4240
box 0 0 6 6
use CELL  85
transform -1 0 2080 0 1 2013
box 0 0 6 6
use CELL  86
transform 1 0 2469 0 1 1253
box 0 0 6 6
use CELL  87
transform -1 0 2086 0 1 4897
box 0 0 6 6
use CELL  88
transform 1 0 2355 0 1 1138
box 0 0 6 6
use CELL  89
transform -1 0 2276 0 1 3796
box 0 0 6 6
use CELL  90
transform 1 0 2300 0 -1 5674
box 0 0 6 6
use CELL  91
transform -1 0 2411 0 -1 5674
box 0 0 6 6
use CELL  92
transform 1 0 2631 0 1 5100
box 0 0 6 6
use CELL  93
transform -1 0 2281 0 1 1573
box 0 0 6 6
use CELL  94
transform -1 0 2764 0 1 4240
box 0 0 6 6
use CELL  95
transform -1 0 2872 0 1 2511
box 0 0 6 6
use CELL  96
transform 1 0 2361 0 1 1253
box 0 0 6 6
use CELL  97
transform -1 0 2140 0 1 3085
box 0 0 6 6
use CELL  98
transform -1 0 2662 0 1 3547
box 0 0 6 6
use CELL  99
transform 1 0 2738 0 1 1573
box 0 0 6 6
use CELL  100
transform 1 0 2797 0 1 1760
box 0 0 6 6
use CELL  101
transform -1 0 2810 0 1 2511
box 0 0 6 6
use CELL  102
transform -1 0 2131 0 1 5755
box 0 0 6 6
use CELL  103
transform -1 0 2314 0 1 1760
box 0 0 6 6
use CELL  104
transform -1 0 2113 0 1 1573
box 0 0 6 6
use CELL  105
transform 1 0 2494 0 1 1253
box 0 0 6 6
use CELL  106
transform -1 0 2738 0 -1 4710
box 0 0 6 6
use CELL  107
transform 1 0 2463 0 -1 5279
box 0 0 6 6
use CELL  108
transform -1 0 2077 0 1 5418
box 0 0 6 6
use CELL  109
transform -1 0 2152 0 1 2511
box 0 0 6 6
use CELL  110
transform -1 0 2374 0 1 5668
box 0 0 6 6
use CELL  111
transform -1 0 2101 0 1 5755
box 0 0 6 6
use CELL  112
transform -1 0 2113 0 1 5551
box 0 0 6 6
use CELL  113
transform -1 0 2175 0 1 4463
box 0 0 6 6
use CELL  114
transform 1 0 2592 0 1 1386
box 0 0 6 6
use CELL  115
transform 1 0 2452 0 1 1386
box 0 0 6 6
use CELL  116
transform -1 0 2933 0 1 2800
box 0 0 6 6
use CELL  117
transform 1 0 2834 0 1 3547
box 0 0 6 6
use CELL  118
transform -1 0 2175 0 1 3322
box 0 0 6 6
use CELL  119
transform -1 0 2086 0 1 1138
box 0 0 6 6
use CELL  120
transform -1 0 2093 0 1 4463
box 0 0 6 6
use CELL  121
transform -1 0 2092 0 1 4240
box 0 0 6 6
use CELL  122
transform -1 0 2954 0 1 2511
box 0 0 6 6
use CELL  123
transform -1 0 2682 0 1 3796
box 0 0 6 6
use CELL  124
transform -1 0 2084 0 1 5418
box 0 0 6 6
use CELL  125
transform -1 0 2898 0 1 2250
box 0 0 6 6
use CELL  126
transform -1 0 2516 0 1 5418
box 0 0 6 6
use CELL  127
transform 1 0 2084 0 -1 2256
box 0 0 6 6
use CELL  128
transform -1 0 2171 0 1 5786
box 0 0 6 6
use CELL  129
transform -1 0 2400 0 1 5418
box 0 0 6 6
use CELL  130
transform 1 0 2599 0 1 1386
box 0 0 6 6
use CELL  131
transform -1 0 2365 0 1 1760
box 0 0 6 6
use CELL  132
transform -1 0 2119 0 1 1253
box 0 0 6 6
use CELL  133
transform -1 0 2091 0 1 1573
box 0 0 6 6
use CELL  134
transform 1 0 2752 0 1 4021
box 0 0 6 6
use CELL  135
transform -1 0 2702 0 1 3085
box 0 0 6 6
use CELL  136
transform -1 0 2806 0 -1 2019
box 0 0 6 6
use CELL  137
transform -1 0 2148 0 1 5795
box 0 0 6 6
use CELL  138
transform -1 0 2249 0 1 2013
box 0 0 6 6
use CELL  139
transform 1 0 2707 0 1 4897
box 0 0 6 6
use CELL  140
transform 1 0 2613 0 1 1386
box 0 0 6 6
use CELL  141
transform -1 0 2443 0 1 5551
box 0 0 6 6
use CELL  142
transform -1 0 2104 0 1 5418
box 0 0 6 6
use CELL  143
transform -1 0 2743 0 1 3322
box 0 0 6 6
use CELL  144
transform -1 0 2120 0 1 5668
box 0 0 6 6
use CELL  145
transform -1 0 2462 0 1 5273
box 0 0 6 6
use CELL  146
transform -1 0 2046 0 1 3547
box 0 0 6 6
use CELL  147
transform -1 0 2252 0 1 5418
box 0 0 6 6
use CELL  148
transform -1 0 2799 0 -1 3553
box 0 0 6 6
use CELL  149
transform -1 0 2160 0 1 5100
box 0 0 6 6
use CELL  150
transform 1 0 2235 0 -1 3328
box 0 0 6 6
use CELL  151
transform -1 0 2134 0 1 3796
box 0 0 6 6
use CELL  152
transform -1 0 2064 0 1 3085
box 0 0 6 6
use CELL  153
transform -1 0 2238 0 1 5551
box 0 0 6 6
use CELL  154
transform -1 0 2134 0 1 2800
box 0 0 6 6
use CELL  155
transform -1 0 2813 0 1 3547
box 0 0 6 6
use CELL  156
transform -1 0 2799 0 1 2013
box 0 0 6 6
use CELL  157
transform -1 0 2757 0 1 4240
box 0 0 6 6
use CELL  158
transform -1 0 2499 0 -1 5557
box 0 0 6 6
use CELL  159
transform -1 0 2143 0 1 5418
box 0 0 6 6
use CELL  160
transform -1 0 2187 0 1 1138
box 0 0 6 6
use CELL  161
transform -1 0 2789 0 1 3322
box 0 0 6 6
use CELL  162
transform -1 0 2662 0 1 3322
box 0 0 6 6
use CELL  163
transform -1 0 2139 0 1 1760
box 0 0 6 6
use CELL  164
transform -1 0 2109 0 1 2800
box 0 0 6 6
use CELL  165
transform -1 0 2509 0 1 5100
box 0 0 6 6
use CELL  166
transform -1 0 2140 0 1 1053
box 0 0 6 6
use CELL  167
transform -1 0 2136 0 1 1010
box 0 0 6 6
use CELL  168
transform 1 0 2209 0 -1 5106
box 0 0 6 6
use CELL  169
transform 1 0 2260 0 1 4021
box 0 0 6 6
use CELL  170
transform 1 0 2500 0 1 5273
box 0 0 6 6
use CELL  171
transform -1 0 2047 0 1 2511
box 0 0 6 6
use CELL  172
transform -1 0 2765 0 1 4021
box 0 0 6 6
use CELL  173
transform -1 0 2740 0 1 4463
box 0 0 6 6
use CELL  174
transform 1 0 2658 0 1 4463
box 0 0 6 6
use CELL  175
transform 1 0 2058 0 1 4240
box 0 0 6 6
use CELL  176
transform -1 0 2096 0 -1 1059
box 0 0 6 6
use CELL  177
transform 1 0 2346 0 1 1253
box 0 0 6 6
use CELL  178
transform -1 0 2139 0 1 5551
box 0 0 6 6
use CELL  179
transform -1 0 2593 0 1 1573
box 0 0 6 6
use CELL  180
transform 1 0 2776 0 1 1760
box 0 0 6 6
use CELL  181
transform -1 0 2561 0 1 5100
box 0 0 6 6
use CELL  182
transform -1 0 2792 0 1 3547
box 0 0 6 6
use CELL  183
transform 1 0 2343 0 -1 5674
box 0 0 6 6
use CELL  184
transform -1 0 2834 0 1 3547
box 0 0 6 6
use CELL  185
transform -1 0 2761 0 1 4463
box 0 0 6 6
use CELL  186
transform -1 0 2233 0 1 4021
box 0 0 6 6
use CELL  187
transform -1 0 2233 0 1 5755
box 0 0 6 6
use CELL  188
transform -1 0 2819 0 1 3322
box 0 0 6 6
use CELL  189
transform -1 0 2813 0 1 3796
box 0 0 6 6
use CELL  190
transform -1 0 2098 0 1 4021
box 0 0 6 6
use CELL  191
transform 1 0 2084 0 -1 5279
box 0 0 6 6
use CELL  192
transform 1 0 2696 0 1 1573
box 0 0 6 6
use CELL  193
transform 1 0 2438 0 1 5418
box 0 0 6 6
use CELL  194
transform -1 0 2827 0 1 2013
box 0 0 6 6
use CELL  195
transform -1 0 2087 0 1 2013
box 0 0 6 6
use CELL  196
transform -1 0 2415 0 1 5273
box 0 0 6 6
use CELL  197
transform -1 0 2117 0 1 3085
box 0 0 6 6
use CELL  198
transform 1 0 2955 0 1 2511
box 0 0 6 6
use CELL  199
transform -1 0 2136 0 -1 4903
box 0 0 6 6
use CELL  200
transform -1 0 2417 0 1 2511
box 0 0 6 6
use CELL  201
transform 1 0 2121 0 1 1573
box 0 0 6 6
use CELL  202
transform -1 0 2542 0 -1 1392
box 0 0 6 6
use CELL  203
transform -1 0 2694 0 1 3796
box 0 0 6 6
use CELL  204
transform -1 0 2794 0 -1 4469
box 0 0 6 6
use CELL  205
transform -1 0 2076 0 1 5273
box 0 0 6 6
use CELL  206
transform -1 0 2367 0 1 5668
box 0 0 6 6
use CELL  207
transform -1 0 2091 0 1 4021
box 0 0 6 6
use CELL  208
transform 1 0 2136 0 1 1138
box 0 0 6 6
use CELL  209
transform -1 0 2098 0 1 1386
box 0 0 6 6
use CELL  210
transform 1 0 2814 0 1 2013
box 0 0 6 6
use CELL  211
transform -1 0 2675 0 1 3796
box 0 0 6 6
use CELL  212
transform -1 0 2787 0 1 4463
box 0 0 6 6
use CELL  213
transform 1 0 2100 0 1 5551
box 0 0 6 6
use CELL  214
transform -1 0 2225 0 1 3085
box 0 0 6 6
use CELL  215
transform 1 0 2790 0 1 3322
box 0 0 6 6
use CELL  216
transform -1 0 2626 0 1 1386
box 0 0 6 6
use CELL  217
transform -1 0 2058 0 1 4463
box 0 0 6 6
use CELL  218
transform 1 0 2120 0 -1 1144
box 0 0 6 6
use CELL  219
transform -1 0 2646 0 1 4463
box 0 0 6 6
use CELL  220
transform -1 0 2782 0 1 3322
box 0 0 6 6
use CELL  221
transform 1 0 2476 0 1 1253
box 0 0 6 6
use CELL  222
transform 1 0 2052 0 -1 4710
box 0 0 6 6
use CELL  223
transform -1 0 2107 0 1 3547
box 0 0 6 6
use CELL  224
transform -1 0 2534 0 1 5273
box 0 0 6 6
use CELL  225
transform -1 0 2393 0 1 5418
box 0 0 6 6
use CELL  226
transform -1 0 2110 0 1 4897
box 0 0 6 6
use CELL  227
transform -1 0 2617 0 1 4897
box 0 0 6 6
use CELL  228
transform 1 0 2791 0 1 3085
box 0 0 6 6
use CELL  229
transform -1 0 2072 0 1 4463
box 0 0 6 6
use CELL  230
transform -1 0 2118 0 1 5418
box 0 0 6 6
use CELL  231
transform -1 0 2243 0 1 4240
box 0 0 6 6
use CELL  232
transform -1 0 2248 0 1 1053
box 0 0 6 6
use CELL  233
transform -1 0 2141 0 1 2800
box 0 0 6 6
use CELL  234
transform -1 0 2095 0 1 2800
box 0 0 6 6
use CELL  235
transform 1 0 2259 0 1 1138
box 0 0 6 6
use CELL  236
transform -1 0 2079 0 1 4463
box 0 0 6 6
use CELL  237
transform 1 0 2508 0 1 1253
box 0 0 6 6
use CELL  238
transform -1 0 2648 0 1 4897
box 0 0 6 6
use CELL  239
transform 1 0 2069 0 -1 2517
box 0 0 6 6
use CELL  240
transform -1 0 2127 0 1 5668
box 0 0 6 6
use CELL  241
transform -1 0 2155 0 1 1053
box 0 0 6 6
use CELL  242
transform -1 0 2046 0 -1 4469
box 0 0 6 6
use CELL  243
transform -1 0 2103 0 1 3322
box 0 0 6 6
use CELL  244
transform -1 0 2016 0 1 3322
box 0 0 6 6
use CELL  245
transform -1 0 2442 0 -1 1144
box 0 0 6 6
use CELL  246
transform -1 0 2124 0 1 3085
box 0 0 6 6
use CELL  247
transform 1 0 2144 0 1 4897
box 0 0 6 6
use CELL  248
transform -1 0 2143 0 1 3322
box 0 0 6 6
use CELL  249
transform -1 0 2150 0 1 2800
box 0 0 6 6
use CELL  250
transform -1 0 2520 0 1 5273
box 0 0 6 6
use CELL  251
transform -1 0 2688 0 1 1573
box 0 0 6 6
use CELL  252
transform 1 0 2731 0 -1 1579
box 0 0 6 6
use CELL  253
transform 1 0 2531 0 1 1253
box 0 0 6 6
use CELL  254
transform -1 0 2150 0 1 4240
box 0 0 6 6
use CELL  255
transform -1 0 2229 0 1 2800
box 0 0 6 6
use CELL  256
transform -1 0 2124 0 1 5755
box 0 0 6 6
use CELL  257
transform -1 0 2786 0 -1 4027
box 0 0 6 6
use CELL  258
transform -1 0 2040 0 1 3796
box 0 0 6 6
use CELL  259
transform -1 0 2141 0 1 3796
box 0 0 6 6
use CELL  260
transform -1 0 2768 0 1 1760
box 0 0 6 6
use CELL  261
transform -1 0 2165 0 1 5755
box 0 0 6 6
use CELL  262
transform -1 0 2169 0 1 1138
box 0 0 6 6
use CELL  263
transform -1 0 2155 0 1 5786
box 0 0 6 6
use CELL  264
transform -1 0 2232 0 1 1053
box 0 0 6 6
use CELL  265
transform -1 0 2725 0 1 3322
box 0 0 6 6
use CELL  266
transform -1 0 2820 0 1 3547
box 0 0 6 6
use CELL  267
transform -1 0 2112 0 1 2511
box 0 0 6 6
use CELL  268
transform -1 0 2676 0 1 3547
box 0 0 6 6
use CELL  269
transform -1 0 2127 0 1 2800
box 0 0 6 6
use CELL  270
transform -1 0 2077 0 1 4021
box 0 0 6 6
use CELL  271
transform -1 0 2398 0 1 1138
box 0 0 6 6
use CELL  272
transform -1 0 2233 0 1 1386
box 0 0 6 6
use CELL  273
transform -1 0 2308 0 -1 1392
box 0 0 6 6
use CELL  274
transform -1 0 2642 0 1 4240
box 0 0 6 6
use CELL  275
transform -1 0 2082 0 1 1053
box 0 0 6 6
use CELL  276
transform 1 0 2538 0 1 1253
box 0 0 6 6
use CELL  277
transform 1 0 2559 0 -1 1259
box 0 0 6 6
use CELL  278
transform -1 0 2209 0 1 1053
box 0 0 6 6
use CELL  279
transform -1 0 2933 0 1 2511
box 0 0 6 6
use CELL  280
transform 1 0 2088 0 1 5551
box 0 0 6 6
use CELL  281
transform -1 0 2052 0 1 5273
box 0 0 6 6
use CELL  282
transform 1 0 2695 0 1 3322
box 0 0 6 6
use CELL  283
transform 1 0 2806 0 1 3322
box 0 0 6 6
use CELL  284
transform 1 0 2058 0 1 5100
box 0 0 6 6
use CELL  285
transform -1 0 2170 0 1 1053
box 0 0 6 6
use CELL  286
transform -1 0 2615 0 1 4021
box 0 0 6 6
use CELL  287
transform -1 0 2220 0 1 5551
box 0 0 6 6
use CELL  288
transform -1 0 2116 0 1 5100
box 0 0 6 6
use CELL  289
transform -1 0 2679 0 1 1573
box 0 0 6 6
use CELL  290
transform -1 0 2120 0 1 1386
box 0 0 6 6
use CELL  291
transform 1 0 2769 0 1 1760
box 0 0 6 6
use CELL  292
transform -1 0 2064 0 1 2013
box 0 0 6 6
use CELL  293
transform -1 0 2195 0 1 2013
box 0 0 6 6
use CELL  294
transform -1 0 2131 0 1 3322
box 0 0 6 6
use CELL  295
transform -1 0 2499 0 1 5273
box 0 0 6 6
use CELL  296
transform 1 0 2085 0 1 1386
box 0 0 6 6
use CELL  297
transform -1 0 2117 0 1 5755
box 0 0 6 6
use CELL  298
transform -1 0 2219 0 1 3796
box 0 0 6 6
use CELL  299
transform 1 0 2064 0 1 5755
box 0 0 6 6
use CELL  300
transform 1 0 2091 0 1 5418
box 0 0 6 6
use CELL  301
transform -1 0 2079 0 1 4897
box 0 0 6 6
use CELL  302
transform -1 0 2905 0 -1 2256
box 0 0 6 6
use CELL  303
transform -1 0 2771 0 1 4240
box 0 0 6 6
use CELL  304
transform -1 0 2678 0 1 4897
box 0 0 6 6
use CELL  305
transform -1 0 2811 0 1 3085
box 0 0 6 6
use CELL  306
transform -1 0 2149 0 1 5755
box 0 0 6 6
use CELL  307
transform -1 0 2110 0 1 5100
box 0 0 6 6
use CELL  308
transform -1 0 2212 0 1 1760
box 0 0 6 6
use CELL  309
transform -1 0 2070 0 1 1138
box 0 0 6 6
use CELL  310
transform 1 0 2364 0 1 1138
box 0 0 6 6
use CELL  311
transform -1 0 2096 0 1 3322
box 0 0 6 6
use CELL  312
transform -1 0 2168 0 1 2511
box 0 0 6 6
use CELL  313
transform -1 0 2736 0 1 4240
box 0 0 6 6
use CELL  314
transform -1 0 2106 0 1 5668
box 0 0 6 6
use CELL  315
transform 1 0 2142 0 -1 5792
box 0 0 6 6
use CELL  316
transform -1 0 2127 0 1 2013
box 0 0 6 6
use CELL  317
transform -1 0 2611 0 1 5100
box 0 0 6 6
use CELL  318
transform -1 0 2132 0 1 5551
box 0 0 6 6
use CELL  319
transform -1 0 2655 0 1 3322
box 0 0 6 6
use CELL  320
transform 1 0 2641 0 -1 1392
box 0 0 6 6
use CELL  321
transform -1 0 2485 0 -1 5557
box 0 0 6 6
use CELL  322
transform 1 0 2074 0 1 1760
box 0 0 6 6
use CELL  323
transform -1 0 2812 0 1 2800
box 0 0 6 6
use CELL  324
transform 1 0 2059 0 -1 4469
box 0 0 6 6
use CELL  325
transform 1 0 2106 0 1 1138
box 0 0 6 6
use CELL  326
transform -1 0 2125 0 1 3547
box 0 0 6 6
use CELL  327
transform -1 0 2212 0 1 3547
box 0 0 6 6
use CELL  328
transform -1 0 2084 0 1 1386
box 0 0 6 6
use CELL  329
transform 1 0 2112 0 1 5273
box 0 0 6 6
use CELL  330
transform 1 0 2700 0 1 4897
box 0 0 6 6
use CELL  331
transform 1 0 2552 0 1 1253
box 0 0 6 6
use CELL  332
transform -1 0 2854 0 1 2250
box 0 0 6 6
use CELL  333
transform -1 0 2622 0 1 4021
box 0 0 6 6
use CELL  334
transform -1 0 2425 0 1 5418
box 0 0 6 6
use CELL  335
transform -1 0 2086 0 1 4463
box 0 0 6 6
use CELL  336
transform 1 0 2801 0 -1 4469
box 0 0 6 6
use CELL  337
transform -1 0 2780 0 1 2013
box 0 0 6 6
use CELL  338
transform -1 0 2145 0 1 1010
box 0 0 6 6
use CELL  339
transform 1 0 2202 0 1 5100
box 0 0 6 6
use CELL  340
transform -1 0 2168 0 1 4463
box 0 0 6 6
use CELL  341
transform -1 0 2603 0 1 4021
box 0 0 6 6
use CELL  342
transform -1 0 2290 0 -1 2256
box 0 0 6 6
use CELL  343
transform -1 0 2780 0 1 3796
box 0 0 6 6
use CELL  344
transform 1 0 2717 0 -1 1579
box 0 0 6 6
use CELL  345
transform -1 0 2194 0 1 4021
box 0 0 6 6
use CELL  346
transform 1 0 2133 0 -1 3553
box 0 0 6 6
use CELL  347
transform -1 0 2153 0 1 2013
box 0 0 6 6
use CELL  348
transform -1 0 2243 0 1 3085
box 0 0 6 6
use CELL  349
transform -1 0 2778 0 1 4240
box 0 0 6 6
use CELL  350
transform -1 0 2152 0 1 1573
box 0 0 6 6
use CELL  351
transform -1 0 2158 0 1 3547
box 0 0 6 6
use CELL  352
transform -1 0 2947 0 1 2511
box 0 0 6 6
use CELL  353
transform 1 0 2099 0 1 1386
box 0 0 6 6
use CELL  354
transform -1 0 2164 0 1 1760
box 0 0 6 6
use CELL  355
transform 1 0 2167 0 1 4021
box 0 0 6 6
use CELL  356
transform -1 0 2068 0 1 2511
box 0 0 6 6
use CELL  357
transform -1 0 2071 0 1 2250
box 0 0 6 6
use CELL  358
transform -1 0 2478 0 1 5551
box 0 0 6 6
use CELL  359
transform -1 0 2246 0 1 5668
box 0 0 6 6
use CELL  360
transform -1 0 2391 0 1 1138
box 0 0 6 6
use CELL  361
transform -1 0 2182 0 -1 1579
box 0 0 6 6
use CELL  362
transform 1 0 2606 0 -1 4246
box 0 0 6 6
use CELL  363
transform -1 0 2252 0 1 2511
box 0 0 6 6
use CELL  364
transform 1 0 2109 0 -1 3802
box 0 0 6 6
use CELL  365
transform -1 0 2257 0 1 5755
box 0 0 6 6
use CELL  366
transform -1 0 2092 0 1 3085
box 0 0 6 6
use CELL  367
transform -1 0 2127 0 1 1386
box 0 0 6 6
use CELL  368
transform -1 0 2261 0 1 4240
box 0 0 6 6
use CELL  369
transform -1 0 2084 0 1 4021
box 0 0 6 6
use CELL  370
transform 1 0 2726 0 -1 4903
box 0 0 6 6
use CELL  371
transform -1 0 2070 0 -1 1579
box 0 0 6 6
use CELL  372
transform -1 0 2984 0 1 2511
box 0 0 6 6
use CELL  373
transform -1 0 2236 0 1 2800
box 0 0 6 6
use CELL  374
transform 1 0 2503 0 -1 5424
box 0 0 6 6
use CELL  375
transform -1 0 2124 0 1 4240
box 0 0 6 6
use CELL  376
transform -1 0 2177 0 1 3796
box 0 0 6 6
use CELL  377
transform 1 0 2121 0 -1 5424
box 0 0 6 6
use CELL  378
transform -1 0 2590 0 1 3547
box 0 0 6 6
use CELL  379
transform -1 0 2153 0 1 5551
box 0 0 6 6
use CELL  380
transform 1 0 2259 0 -1 5557
box 0 0 6 6
use CELL  381
transform 1 0 2283 0 1 1138
box 0 0 6 6
use CELL  382
transform -1 0 2231 0 1 1253
box 0 0 6 6
use CELL  383
transform -1 0 2155 0 1 5795
box 0 0 6 6
use CELL  384
transform 1 0 2292 0 1 1138
box 0 0 6 6
use CELL  385
transform -1 0 2086 0 1 4704
box 0 0 6 6
use CELL  386
transform -1 0 2698 0 1 4704
box 0 0 6 6
use CELL  387
transform -1 0 2131 0 1 2511
box 0 0 6 6
use CELL  388
transform -1 0 2164 0 1 2250
box 0 0 6 6
use CELL  389
transform -1 0 2682 0 1 4463
box 0 0 6 6
use CELL  390
transform -1 0 2085 0 1 3085
box 0 0 6 6
use CELL  391
transform -1 0 2082 0 1 3796
box 0 0 6 6
use CELL  392
transform 1 0 2213 0 -1 5761
box 0 0 6 6
use CELL  393
transform -1 0 2094 0 1 2013
box 0 0 6 6
use CELL  394
transform -1 0 2956 0 1 2250
box 0 0 6 6
use CELL  395
transform -1 0 2940 0 1 2511
box 0 0 6 6
use CELL  396
transform -1 0 2903 0 1 2800
box 0 0 6 6
use CELL  397
transform -1 0 2840 0 -1 2517
box 0 0 6 6
use CELL  398
transform -1 0 2747 0 1 4463
box 0 0 6 6
use CELL  399
transform -1 0 2100 0 1 2511
box 0 0 6 6
use CELL  400
transform -1 0 2098 0 1 1573
box 0 0 6 6
use CELL  401
transform -1 0 2263 0 1 1573
box 0 0 6 6
use CELL  402
transform 1 0 2304 0 1 1138
box 0 0 6 6
use CELL  403
transform -1 0 2089 0 1 3547
box 0 0 6 6
use CELL  404
transform -1 0 2912 0 1 2250
box 0 0 6 6
use CELL  405
transform 1 0 2091 0 1 5273
box 0 0 6 6
use CELL  406
transform -1 0 2548 0 1 5273
box 0 0 6 6
use CELL  407
transform -1 0 2065 0 1 4897
box 0 0 6 6
use CELL  408
transform -1 0 2085 0 1 1253
box 0 0 6 6
use CELL  409
transform -1 0 2783 0 1 3085
box 0 0 6 6
use CELL  410
transform 1 0 2458 0 1 5551
box 0 0 6 6
use CELL  411
transform 1 0 2129 0 1 1138
box 0 0 6 6
use CELL  412
transform 1 0 2465 0 1 5551
box 0 0 6 6
use CELL  413
transform -1 0 2157 0 1 4897
box 0 0 6 6
use CELL  414
transform -1 0 2720 0 1 3085
box 0 0 6 6
use CELL  415
transform -1 0 2597 0 1 5100
box 0 0 6 6
use CELL  416
transform -1 0 2861 0 1 2250
box 0 0 6 6
use CELL  417
transform -1 0 2450 0 1 5551
box 0 0 6 6
use CELL  418
transform -1 0 2106 0 1 2013
box 0 0 6 6
use CELL  419
transform -1 0 2078 0 1 5100
box 0 0 6 6
use CELL  420
transform -1 0 2738 0 -1 1766
box 0 0 6 6
use CELL  421
transform -1 0 2889 0 1 2800
box 0 0 6 6
use CELL  422
transform -1 0 2750 0 1 4240
box 0 0 6 6
use CELL  423
transform -1 0 2848 0 1 2013
box 0 0 6 6
use CELL  424
transform -1 0 2072 0 1 4704
box 0 0 6 6
use CELL  425
transform -1 0 2917 0 1 2800
box 0 0 6 6
use CELL  426
transform -1 0 2093 0 1 4704
box 0 0 6 6
use CELL  427
transform -1 0 2146 0 1 5273
box 0 0 6 6
use CELL  428
transform -1 0 2818 0 1 2250
box 0 0 6 6
use CELL  429
transform -1 0 2058 0 1 4897
box 0 0 6 6
use CELL  430
transform -1 0 2654 0 1 4240
box 0 0 6 6
use CELL  431
transform -1 0 2226 0 1 5755
box 0 0 6 6
use CELL  432
transform -1 0 2398 0 1 5668
box 0 0 6 6
use CELL  433
transform -1 0 2140 0 1 1253
box 0 0 6 6
use CELL  434
transform -1 0 2773 0 1 3796
box 0 0 6 6
use CELL  435
transform -1 0 2125 0 1 4704
box 0 0 6 6
use CELL  436
transform -1 0 2040 0 1 2511
box 0 0 6 6
use CELL  437
transform -1 0 2865 0 1 2511
box 0 0 6 6
use CELL  438
transform -1 0 2540 0 1 3796
box 0 0 6 6
use CELL  439
transform 1 0 2399 0 1 1138
box 0 0 6 6
use CELL  440
transform -1 0 2070 0 1 1386
box 0 0 6 6
use CELL  441
transform 1 0 2798 0 1 3085
box 0 0 6 6
use CELL  442
transform -1 0 2108 0 1 3796
box 0 0 6 6
use CELL  443
transform 1 0 2590 0 1 4021
box 0 0 6 6
use CELL  444
transform -1 0 2858 0 1 2511
box 0 0 6 6
use CELL  445
transform -1 0 2484 0 1 5418
box 0 0 6 6
use CELL  446
transform -1 0 2754 0 1 3796
box 0 0 6 6
use CELL  447
transform -1 0 2118 0 1 4463
box 0 0 6 6
use CELL  448
transform -1 0 2720 0 1 4240
box 0 0 6 6
use CELL  449
transform 1 0 2741 0 1 1760
box 0 0 6 6
use CELL  450
transform 1 0 2103 0 -1 2256
box 0 0 6 6
use CELL  451
transform -1 0 2138 0 1 2511
box 0 0 6 6
use CELL  452
transform -1 0 2052 0 -1 1766
box 0 0 6 6
use CELL  453
transform -1 0 2147 0 1 3085
box 0 0 6 6
use CELL  454
transform -1 0 2146 0 1 5100
box 0 0 6 6
use CELL  455
transform -1 0 2134 0 1 2250
box 0 0 6 6
use CELL  456
transform -1 0 2150 0 -1 3328
box 0 0 6 6
use CELL  457
transform -1 0 2157 0 1 2250
box 0 0 6 6
use CELL  458
transform -1 0 2132 0 1 3547
box 0 0 6 6
use CELL  459
transform -1 0 2143 0 1 4897
box 0 0 6 6
use CELL  460
transform 1 0 2071 0 -1 1144
box 0 0 6 6
use CELL  461
transform -1 0 2796 0 1 1760
box 0 0 6 6
use CELL  462
transform -1 0 2073 0 1 1760
box 0 0 6 6
use CELL  463
transform -1 0 2629 0 1 4897
box 0 0 6 6
use CELL  464
transform -1 0 2436 0 1 5551
box 0 0 6 6
use CELL  465
transform -1 0 2761 0 1 3322
box 0 0 6 6
use CELL  466
transform -1 0 2103 0 1 1760
box 0 0 6 6
use CELL  467
transform 1 0 2804 0 -1 1766
box 0 0 6 6
use CELL  468
transform -1 0 2121 0 1 1760
box 0 0 6 6
use CELL  469
transform -1 0 2119 0 1 1053
box 0 0 6 6
use CELL  470
transform -1 0 2224 0 1 1386
box 0 0 6 6
use CELL  471
transform -1 0 2896 0 1 2800
box 0 0 6 6
use CELL  472
transform 1 0 2677 0 -1 2806
box 0 0 6 6
use CELL  473
transform -1 0 2119 0 1 2511
box 0 0 6 6
use CELL  474
transform 1 0 2627 0 1 1386
box 0 0 6 6
use CELL  475
transform -1 0 2133 0 1 3085
box 0 0 6 6
use CELL  476
transform -1 0 2541 0 1 5273
box 0 0 6 6
use CELL  477
transform -1 0 2674 0 1 1760
box 0 0 6 6
use CELL  478
transform -1 0 2070 0 1 3547
box 0 0 6 6
use CELL  479
transform -1 0 2077 0 1 1573
box 0 0 6 6
use CELL  480
transform -1 0 2145 0 -1 2517
box 0 0 6 6
use CELL  481
transform -1 0 2825 0 1 3085
box 0 0 6 6
use CELL  482
transform -1 0 2084 0 1 3322
box 0 0 6 6
use CELL  483
transform -1 0 2091 0 1 5418
box 0 0 6 6
use CELL  484
transform -1 0 2103 0 1 1053
box 0 0 6 6
use CELL  485
transform -1 0 2840 0 1 2800
box 0 0 6 6
use CELL  486
transform -1 0 2492 0 1 5551
box 0 0 6 6
use CELL  487
transform -1 0 2058 0 1 4021
box 0 0 6 6
use CELL  488
transform 1 0 2147 0 -1 5279
box 0 0 6 6
use CELL  489
transform -1 0 2118 0 1 4704
box 0 0 6 6
use CELL  490
transform -1 0 2094 0 1 5668
box 0 0 6 6
use CELL  491
transform -1 0 2429 0 1 5273
box 0 0 6 6
use CELL  492
transform -1 0 2896 0 1 2511
box 0 0 6 6
use CELL  493
transform -1 0 2891 0 1 2250
box 0 0 6 6
use CELL  494
transform -1 0 2557 0 1 1386
box 0 0 6 6
use CELL  495
transform -1 0 2064 0 1 1253
box 0 0 6 6
use CELL  496
transform 1 0 2920 0 1 2800
box 0 0 6 6
use CELL  497
transform 1 0 2071 0 1 1386
box 0 0 6 6
use CELL  498
transform -1 0 2126 0 1 1253
box 0 0 6 6
use CELL  499
transform 1 0 2200 0 1 4897
box 0 0 6 6
use CELL  500
transform -1 0 2801 0 1 4463
box 0 0 6 6
use CELL  501
transform -1 0 2582 0 1 4704
box 0 0 6 6
use CELL  502
transform -1 0 2089 0 1 1053
box 0 0 6 6
use CELL  503
transform -1 0 2604 0 1 5100
box 0 0 6 6
use CELL  504
transform -1 0 2222 0 1 5418
box 0 0 6 6
use CELL  505
transform -1 0 2192 0 1 4704
box 0 0 6 6
use CELL  506
transform -1 0 2146 0 1 5551
box 0 0 6 6
use CELL  507
transform 1 0 2703 0 1 1573
box 0 0 6 6
use CELL  508
transform -1 0 2150 0 1 2250
box 0 0 6 6
use CELL  509
transform 1 0 2069 0 -1 3802
box 0 0 6 6
use CELL  510
transform -1 0 2164 0 1 5786
box 0 0 6 6
use CELL  511
transform 1 0 2105 0 1 5273
box 0 0 6 6
use CELL  512
transform -1 0 2848 0 1 3085
box 0 0 6 6
use CELL  513
transform -1 0 2695 0 1 1573
box 0 0 6 6
use CELL  514
transform -1 0 2153 0 1 5100
box 0 0 6 6
use CELL  515
transform 1 0 2097 0 -1 5106
box 0 0 6 6
use CELL  516
transform -1 0 2078 0 1 4240
box 0 0 6 6
use CELL  517
transform 1 0 2450 0 1 5418
box 0 0 6 6
use CELL  518
transform -1 0 2199 0 -1 4903
box 0 0 6 6
use CELL  519
transform -1 0 2231 0 1 4240
box 0 0 6 6
use CELL  520
transform 1 0 2065 0 1 3085
box 0 0 6 6
use CELL  521
transform 1 0 2750 0 1 2013
box 0 0 6 6
use CELL  522
transform -1 0 2790 0 1 3085
box 0 0 6 6
use CELL  523
transform -1 0 2789 0 1 1760
box 0 0 6 6
use CELL  524
transform 1 0 2088 0 1 5755
box 0 0 6 6
use CELL  525
transform 1 0 2188 0 1 3547
box 0 0 6 6
use CELL  526
transform -1 0 2238 0 1 1253
box 0 0 6 6
use CELL  527
transform -1 0 2223 0 1 1053
box 0 0 6 6
use CELL  528
transform -1 0 2908 0 1 2511
box 0 0 6 6
use CELL  529
transform -1 0 2085 0 1 4240
box 0 0 6 6
use CELL  530
transform -1 0 2139 0 1 5273
box 0 0 6 6
use CELL  531
transform -1 0 2672 0 1 1573
box 0 0 6 6
use CELL  532
transform -1 0 2407 0 1 5418
box 0 0 6 6
use CELL  533
transform -1 0 2078 0 1 1253
box 0 0 6 6
use CELL  534
transform -1 0 2244 0 1 4463
box 0 0 6 6
use CELL  535
transform -1 0 2554 0 1 5100
box 0 0 6 6
use CELL  536
transform -1 0 2253 0 1 4463
box 0 0 6 6
use CELL  537
transform -1 0 2332 0 1 4021
box 0 0 6 6
use CELL  538
transform -1 0 2143 0 1 4021
box 0 0 6 6
use CELL  539
transform -1 0 2670 0 1 4704
box 0 0 6 6
use CELL  540
transform -1 0 2101 0 1 1253
box 0 0 6 6
use CELL  541
transform -1 0 2761 0 -1 1766
box 0 0 6 6
use CELL  542
transform -1 0 2124 0 1 4897
box 0 0 6 6
use CELL  543
transform -1 0 2239 0 1 5668
box 0 0 6 6
use CELL  544
transform -1 0 2573 0 1 5100
box 0 0 6 6
use CELL  545
transform -1 0 2674 0 1 3322
box 0 0 6 6
use CELL  546
transform -1 0 2146 0 1 1760
box 0 0 6 6
use CELL  547
transform -1 0 2122 0 1 3796
box 0 0 6 6
use CELL  548
transform -1 0 2061 0 1 3796
box 0 0 6 6
use CELL  549
transform -1 0 2070 0 1 5418
box 0 0 6 6
use CELL  550
transform 1 0 2569 0 -1 1392
box 0 0 6 6
use CELL  551
transform -1 0 2806 0 1 3796
box 0 0 6 6
use CELL  552
transform -1 0 2739 0 1 4021
box 0 0 6 6
use CELL  553
transform -1 0 2289 0 1 5551
box 0 0 6 6
use CELL  554
transform 1 0 2920 0 1 2511
box 0 0 6 6
use CELL  555
transform -1 0 2234 0 1 5418
box 0 0 6 6
use CELL  556
transform -1 0 2731 0 1 4704
box 0 0 6 6
use CELL  557
transform -1 0 2657 0 1 3796
box 0 0 6 6
use CELL  558
transform -1 0 2947 0 -1 2806
box 0 0 6 6
use CELL  559
transform 1 0 2391 0 1 1253
box 0 0 6 6
use CELL  560
transform -1 0 2168 0 1 3322
box 0 0 6 6
use CELL  561
transform -1 0 2111 0 1 5418
box 0 0 6 6
use CELL  562
transform -1 0 2160 0 1 5273
box 0 0 6 6
use CELL  563
transform -1 0 2405 0 1 5668
box 0 0 6 6
use CELL  564
transform -1 0 2059 0 1 5273
box 0 0 6 6
use CELL  565
transform 1 0 2071 0 -1 5761
box 0 0 6 6
use CELL  566
transform -1 0 2910 0 1 2800
box 0 0 6 6
use CELL  567
transform -1 0 2732 0 1 4021
box 0 0 6 6
use CELL  568
transform -1 0 2421 0 1 1138
box 0 0 6 6
use CELL  569
transform -1 0 2065 0 1 4704
box 0 0 6 6
use CELL  570
transform -1 0 2102 0 1 2250
box 0 0 6 6
use CELL  571
transform -1 0 2216 0 1 4704
box 0 0 6 6
use CELL  572
transform -1 0 2266 0 1 2250
box 0 0 6 6
use CELL  573
transform 1 0 2786 0 -1 4246
box 0 0 6 6
use CELL  574
transform 1 0 2678 0 -1 4710
box 0 0 6 6
use CELL  575
transform -1 0 2120 0 1 5551
box 0 0 6 6
use CELL  576
transform -1 0 2385 0 -1 1259
box 0 0 6 6
use CELL  577
transform 1 0 2064 0 -1 4027
box 0 0 6 6
use CELL  578
transform -1 0 2120 0 1 1573
box 0 0 6 6
use CELL  579
transform -1 0 2730 0 1 1573
box 0 0 6 6
use CELL  580
transform -1 0 2416 0 1 1386
box 0 0 6 6
use CELL  581
transform -1 0 2016 0 1 2250
box 0 0 6 6
use CELL  582
transform -1 0 2070 0 1 3322
box 0 0 6 6
use CELL  583
transform -1 0 2054 0 -1 2517
box 0 0 6 6
use CELL  584
transform 1 0 2607 0 -1 4710
box 0 0 6 6
use CELL  585
transform -1 0 2131 0 1 4240
box 0 0 6 6
use CELL  586
transform -1 0 2064 0 1 2250
box 0 0 6 6
use CELL  587
transform 1 0 2679 0 1 4897
box 0 0 6 6
use CELL  588
transform 1 0 2957 0 -1 2256
box 0 0 6 6
use CELL  589
transform -1 0 2448 0 1 1138
box 0 0 6 6
use CELL  590
transform -1 0 2210 0 1 5755
box 0 0 6 6
use CELL  591
transform 1 0 2774 0 1 4463
box 0 0 6 6
use CELL  592
transform -1 0 2665 0 1 1573
box 0 0 6 6
use CELL  593
transform -1 0 2102 0 1 2800
box 0 0 6 6
use CELL  594
transform 1 0 2471 0 -1 5424
box 0 0 6 6
use CELL  595
transform -1 0 2625 0 1 5100
box 0 0 6 6
use CELL  596
transform -1 0 2785 0 1 3547
box 0 0 6 6
use CELL  597
transform -1 0 2435 0 1 1138
box 0 0 6 6
use CELL  598
transform -1 0 2117 0 1 4897
box 0 0 6 6
use CELL  599
transform -1 0 2817 0 1 1760
box 0 0 6 6
use CELL  600
transform -1 0 2855 0 1 2013
box 0 0 6 6
use CELL  601
transform -1 0 2156 0 1 4704
box 0 0 6 6
use CELL  602
transform -1 0 2176 0 1 1760
box 0 0 6 6
use CELL  603
transform -1 0 2818 0 -1 3091
box 0 0 6 6
use CELL  604
transform 1 0 2457 0 1 5418
box 0 0 6 6
use CELL  605
transform -1 0 2077 0 1 2800
box 0 0 6 6
use CELL  606
transform -1 0 2764 0 1 2800
box 0 0 6 6
use CELL  607
transform -1 0 2422 0 1 5273
box 0 0 6 6
use CELL  608
transform -1 0 2947 0 1 2250
box 0 0 6 6
use CELL  609
transform -1 0 2070 0 1 2800
box 0 0 6 6
use CELL  610
transform -1 0 2099 0 1 3085
box 0 0 6 6
use CELL  611
transform -1 0 2754 0 -1 4469
box 0 0 6 6
use CELL  612
transform -1 0 2649 0 1 4704
box 0 0 6 6
use CELL  613
transform -1 0 2775 0 1 3322
box 0 0 6 6
use CELL  614
transform 1 0 2412 0 1 5668
box 0 0 6 6
use CELL  615
transform -1 0 2779 0 -1 4027
box 0 0 6 6
use CELL  616
transform 1 0 2579 0 1 5100
box 0 0 6 6
use CELL  617
transform -1 0 2201 0 1 3085
box 0 0 6 6
use CELL  618
transform -1 0 2136 0 -1 4027
box 0 0 6 6
use CELL  619
transform -1 0 2165 0 1 3085
box 0 0 6 6
use CELL  620
transform 1 0 2545 0 1 1253
box 0 0 6 6
use CELL  621
transform -1 0 2834 0 1 2013
box 0 0 6 6
use CELL  622
transform -1 0 2977 0 1 2511
box 0 0 6 6
use CELL  623
transform -1 0 2731 0 1 1760
box 0 0 6 6
use CELL  624
transform -1 0 2677 0 1 4704
box 0 0 6 6
use CELL  625
transform -1 0 2806 0 1 3547
box 0 0 6 6
use CELL  626
transform -1 0 2342 0 1 5668
box 0 0 6 6
use CELL  627
transform -1 0 2078 0 1 3085
box 0 0 6 6
use CELL  628
transform -1 0 2725 0 -1 4027
box 0 0 6 6
use CELL  629
transform 1 0 2524 0 1 1253
box 0 0 6 6
use CELL  630
transform -1 0 2119 0 1 1138
box 0 0 6 6
use CELL  631
transform -1 0 2111 0 1 4704
box 0 0 6 6
use CELL  632
transform -1 0 2719 0 1 1760
box 0 0 6 6
use CELL  633
transform -1 0 2689 0 1 4463
box 0 0 6 6
use CELL  634
transform 1 0 2152 0 -1 1392
box 0 0 6 6
use CELL  635
transform 1 0 2820 0 1 1760
box 0 0 6 6
use CELL  636
transform -1 0 2165 0 1 4704
box 0 0 6 6
use CELL  637
transform 1 0 2122 0 1 5100
box 0 0 6 6
use CELL  638
transform -1 0 2169 0 1 2800
box 0 0 6 6
use CELL  639
transform -1 0 2108 0 1 5755
box 0 0 6 6
use CELL  640
transform -1 0 2545 0 1 5100
box 0 0 6 6
use CELL  641
transform -1 0 2245 0 1 3547
box 0 0 6 6
use CELL  642
transform -1 0 2136 0 1 5418
box 0 0 6 6
use CELL  643
transform -1 0 2841 0 1 3085
box 0 0 6 6
use CELL  644
transform -1 0 2146 0 1 2013
box 0 0 6 6
use CELL  645
transform 1 0 2079 0 -1 5106
box 0 0 6 6
use CELL  646
transform 1 0 2849 0 1 3085
box 0 0 6 6
use CELL  647
transform -1 0 2138 0 1 4240
box 0 0 6 6
use CELL  648
transform -1 0 2216 0 1 1053
box 0 0 6 6
use CELL  649
transform -1 0 2766 0 1 3796
box 0 0 6 6
use CELL  650
transform -1 0 2092 0 1 1253
box 0 0 6 6
use CELL  651
transform -1 0 2678 0 1 2013
box 0 0 6 6
use CELL  652
transform 1 0 2065 0 -1 5106
box 0 0 6 6
use CELL  653
transform -1 0 2739 0 1 4897
box 0 0 6 6
use CELL  654
transform -1 0 2388 0 1 4463
box 0 0 6 6
use CELL  655
transform -1 0 2919 0 1 2250
box 0 0 6 6
use CELL  656
transform -1 0 2742 0 1 3547
box 0 0 6 6
use CELL  657
transform -1 0 2489 0 1 3085
box 0 0 6 6
use CELL  658
transform -1 0 2940 0 1 2800
box 0 0 6 6
use CELL  659
transform -1 0 2077 0 1 3322
box 0 0 6 6
use CELL  660
transform 1 0 2766 0 -1 4027
box 0 0 6 6
use CELL  661
transform -1 0 2288 0 1 4704
box 0 0 6 6
use CELL  662
transform -1 0 2717 0 1 4704
box 0 0 6 6
use CELL  663
transform 1 0 2927 0 1 2250
box 0 0 6 6
use CELL  664
transform -1 0 2940 0 1 2250
box 0 0 6 6
use CELL  665
transform -1 0 2143 0 1 2250
box 0 0 6 6
use CELL  666
transform -1 0 2189 0 1 3796
box 0 0 6 6
use CELL  667
transform -1 0 2457 0 1 5551
box 0 0 6 6
use CELL  668
transform -1 0 2125 0 1 4463
box 0 0 6 6
use CELL  669
transform -1 0 2084 0 1 1573
box 0 0 6 6
use CELL  670
transform 1 0 2464 0 1 5418
box 0 0 6 6
use CELL  671
transform -1 0 2852 0 -1 2806
box 0 0 6 6
use CELL  672
transform -1 0 2100 0 1 4463
box 0 0 6 6
use CELL  673
transform -1 0 2093 0 1 1138
box 0 0 6 6
use CELL  674
transform -1 0 2768 0 1 2013
box 0 0 6 6
use CELL  675
transform -1 0 2820 0 1 3796
box 0 0 6 6
use CELL  676
transform -1 0 2118 0 1 2013
box 0 0 6 6
use CELL  677
transform -1 0 2968 0 1 2511
box 0 0 6 6
use CELL  678
transform -1 0 2523 0 1 1253
box 0 0 6 6
use CELL  679
transform -1 0 2624 0 1 4240
box 0 0 6 6
use CELL  680
transform -1 0 2805 0 1 3322
box 0 0 6 6
use CELL  681
transform 1 0 2184 0 1 5273
box 0 0 6 6
use CELL  682
transform -1 0 2732 0 1 3085
box 0 0 6 6
use CELL  683
transform 1 0 2835 0 -1 2019
box 0 0 6 6
use CELL  684
transform -1 0 2792 0 1 3796
box 0 0 6 6
use CELL  685
transform -1 0 2292 0 1 3322
box 0 0 6 6
use CELL  686
transform -1 0 2391 0 1 5551
box 0 0 6 6
use CELL  687
transform -1 0 2072 0 1 4897
box 0 0 6 6
use CELL  688
transform -1 0 2132 0 1 4704
box 0 0 6 6
use CELL  689
transform 1 0 2154 0 -1 1016
box 0 0 6 6
use CELL  690
transform -1 0 2778 0 1 3547
box 0 0 6 6
use CELL  691
transform -1 0 2882 0 1 2800
box 0 0 6 6
use CELL  692
transform -1 0 2133 0 1 1253
box 0 0 6 6
use CELL  693
transform -1 0 2071 0 1 2013
box 0 0 6 6
use CELL  694
transform -1 0 2873 0 1 2250
box 0 0 6 6
use CELL  695
transform 1 0 2151 0 1 2800
box 0 0 6 6
use CELL  696
transform -1 0 2710 0 1 4704
box 0 0 6 6
use CELL  697
transform -1 0 2089 0 1 1760
box 0 0 6 6
use CELL  698
transform -1 0 2641 0 1 4897
box 0 0 6 6
use CELL  699
transform -1 0 2618 0 1 5100
box 0 0 6 6
use CELL  700
transform -1 0 2403 0 -1 5557
box 0 0 6 6
use CELL  701
transform 1 0 2713 0 1 4463
box 0 0 6 6
use CELL  702
transform -1 0 2513 0 1 5273
box 0 0 6 6
use CELL  703
transform -1 0 2105 0 1 4021
box 0 0 6 6
use CELL  704
transform -1 0 2644 0 1 5100
box 0 0 6 6
use CELL  705
transform -1 0 2129 0 1 4021
box 0 0 6 6
use CELL  706
transform -1 0 2669 0 1 3547
box 0 0 6 6
use CELL  707
transform -1 0 2507 0 1 1253
box 0 0 6 6
use CELL  708
transform -1 0 2291 0 1 2013
box 0 0 6 6
use CELL  709
transform -1 0 2213 0 1 5551
box 0 0 6 6
use CELL  710
transform -1 0 2089 0 1 3796
box 0 0 6 6
use CELL  711
transform -1 0 2819 0 1 2800
box 0 0 6 6
use CELL  712
transform -1 0 2754 0 1 1760
box 0 0 6 6
use CELL  713
transform -1 0 2147 0 1 1253
box 0 0 6 6
use CELL  714
transform -1 0 2834 0 1 3085
box 0 0 6 6
use CELL  715
transform -1 0 2077 0 -1 3553
box 0 0 6 6
use CELL  716
transform -1 0 2273 0 1 1053
box 0 0 6 6
use CELL  717
transform 1 0 2422 0 1 1138
box 0 0 6 6
use CELL  718
transform -1 0 2527 0 1 5273
box 0 0 6 6
use CELL  719
transform -1 0 2424 0 1 5551
box 0 0 6 6
use CELL  720
transform 1 0 2634 0 1 1386
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 2312 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 2332 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 2497 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 2088 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 2083 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 2375 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 2347 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 2417 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 2298 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 2335 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 2292 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 2371 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 2380 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 2380 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 2399 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 2503 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 2420 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 2530 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 2399 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 2178 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 2107 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 2224 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 2274 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 2237 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 2274 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 2110 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 2780 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 2879 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 2896 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 2840 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 2753 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 2725 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 2742 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 2140 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 2206 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 2152 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 2724 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 2240 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 2322 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 2491 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 2474 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 2536 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 2381 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 2206 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 2198 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 2175 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 2189 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 2488 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 2458 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 2071 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 2380 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 2360 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 2080 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 2387 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 2224 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 2679 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 2738 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 2768 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 2861 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 2884 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 2819 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 2732 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 2707 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 2727 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 2712 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 2706 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 2690 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 2695 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 2619 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 2797 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 2713 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 2698 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 2768 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 2625 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 2745 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 2728 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 2756 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 2173 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 2180 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 2118 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 2405 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 2273 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 2489 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 2398 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 2404 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 2272 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 2152 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 2133 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 2140 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 2468 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 2709 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 2715 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 2652 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 2634 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 2693 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 2542 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 2622 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 2582 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 2540 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 2545 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 2491 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 2254 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 2379 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 2257 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 2382 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 2488 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 2575 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 2299 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-109
transform 1 0 2111 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-110
transform 1 0 2369 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-111
transform 1 0 2401 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-112
transform 1 0 2094 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-113
transform 1 0 2245 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-114
transform 1 0 2195 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-115
transform 1 0 2292 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-116
transform 1 0 2091 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-117
transform 1 0 2092 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-118
transform 1 0 2099 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-119
transform 1 0 2106 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-120
transform 1 0 2230 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-121
transform 1 0 2182 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-122
transform 1 0 2256 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-123
transform 1 0 2264 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-124
transform 1 0 2192 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-125
transform 1 0 2109 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-126
transform 1 0 2109 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-127
transform 1 0 2435 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-128
transform 1 0 2350 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-129
transform 1 0 2514 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-130
transform 1 0 2734 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-131
transform 1 0 2828 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-132
transform 1 0 2524 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-133
transform 1 0 2612 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-134
transform 1 0 2662 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-135
transform 1 0 2584 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-136
transform 1 0 2434 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-137
transform 1 0 2666 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-138
transform 1 0 2658 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-139
transform 1 0 2669 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-140
transform 1 0 2661 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-141
transform 1 0 2725 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-142
transform 1 0 2702 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-143
transform 1 0 2664 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-144
transform 1 0 2730 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-145
transform 1 0 2730 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-146
transform 1 0 2464 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-147
transform 1 0 2507 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-148
transform 1 0 2563 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-149
transform 1 0 2186 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-150
transform 1 0 2182 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-151
transform 1 0 2159 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-152
transform 1 0 2389 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-153
transform 1 0 2286 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-154
transform 1 0 2154 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-155
transform 1 0 2188 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-156
transform 1 0 2198 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-157
transform 1 0 2151 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-158
transform 1 0 2161 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-159
transform 1 0 2578 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-160
transform 1 0 2564 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-161
transform 1 0 2581 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-162
transform 1 0 2515 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-163
transform 1 0 2646 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-164
transform 1 0 2739 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-165
transform 1 0 2780 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-166
transform 1 0 2349 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-167
transform 1 0 2457 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-168
transform 1 0 2518 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-169
transform 1 0 2635 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-170
transform 1 0 2707 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-171
transform 1 0 2696 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-172
transform 1 0 2352 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-173
transform 1 0 2460 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-174
transform 1 0 2521 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-175
transform 1 0 2638 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-176
transform 1 0 2232 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-177
transform 1 0 2316 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-178
transform 1 0 2445 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-179
transform 1 0 2506 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-180
transform 1 0 2599 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-181
transform 1 0 2710 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-182
transform 1 0 2699 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-183
transform 1 0 2785 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-184
transform 1 0 2846 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-185
transform 1 0 2731 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-186
transform 1 0 2702 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-187
transform 1 0 2662 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-188
transform 1 0 2560 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-189
transform 1 0 2474 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-190
transform 1 0 2595 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-191
transform 1 0 2488 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-192
transform 1 0 2645 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-193
transform 1 0 2584 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-194
transform 1 0 2465 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-195
transform 1 0 2616 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-196
transform 1 0 2486 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-197
transform 1 0 2506 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-198
transform 1 0 2485 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-199
transform 1 0 2277 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-200
transform 1 0 2271 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-201
transform 1 0 2260 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-202
transform 1 0 2291 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-203
transform 1 0 2317 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-204
transform 1 0 2312 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-205
transform 1 0 2374 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-206
transform 1 0 2426 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-207
transform 1 0 2735 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-208
transform 1 0 2606 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-209
transform 1 0 2509 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-210
transform 1 0 2354 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-211
transform 1 0 2554 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-212
transform 1 0 2434 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-213
transform 1 0 2395 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-214
transform 1 0 2355 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-215
transform 1 0 2268 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-216
transform 1 0 2222 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-217
transform 1 0 2251 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-218
transform 1 0 2245 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-219
transform 1 0 2254 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-220
transform 1 0 2345 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-221
transform 1 0 2626 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-222
transform 1 0 2121 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-223
transform 1 0 2311 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-224
transform 1 0 2310 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-225
transform 1 0 2175 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-226
transform 1 0 2174 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-227
transform 1 0 2173 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-228
transform 1 0 2177 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-229
transform 1 0 2449 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-230
transform 1 0 2445 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-231
transform 1 0 2438 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-232
transform 1 0 2410 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-233
transform 1 0 2396 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-234
transform 1 0 2374 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-235
transform 1 0 2330 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-236
transform 1 0 2404 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-237
transform 1 0 2392 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-238
transform 1 0 2190 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-239
transform 1 0 2490 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-240
transform 1 0 2493 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-241
transform 1 0 2648 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-242
transform 1 0 2585 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-243
transform 1 0 2406 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-244
transform 1 0 2374 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-245
transform 1 0 2233 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-246
transform 1 0 2481 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-247
transform 1 0 2605 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-248
transform 1 0 2622 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-249
transform 1 0 2608 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-250
transform 1 0 2545 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-251
transform 1 0 2441 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-252
transform 1 0 2694 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-253
transform 1 0 2697 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-254
transform 1 0 2708 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-255
transform 1 0 2719 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-256
transform 1 0 2625 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-257
transform 1 0 2651 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-258
transform 1 0 2588 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-259
transform 1 0 2487 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-260
transform 1 0 2444 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-261
transform 1 0 2427 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-262
transform 1 0 2156 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-263
transform 1 0 2271 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-264
transform 1 0 2461 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-265
transform 1 0 2416 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-266
transform 1 0 2444 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-267
transform 1 0 2580 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-268
transform 1 0 2393 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-269
transform 1 0 2530 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-270
transform 1 0 2630 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-271
transform 1 0 2162 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-272
transform 1 0 2165 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-273
transform 1 0 2221 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-274
transform 1 0 2201 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-275
transform 1 0 2197 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-276
transform 1 0 2207 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-277
transform 1 0 2164 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-278
transform 1 0 2156 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-279
transform 1 0 2177 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-280
transform 1 0 2217 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-281
transform 1 0 2240 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-282
transform 1 0 2245 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-283
transform 1 0 2248 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-284
transform 1 0 2386 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-285
transform 1 0 2389 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-286
transform 1 0 2412 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-287
transform 1 0 2432 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-288
transform 1 0 2469 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-289
transform 1 0 2561 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-290
transform 1 0 2617 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-291
transform 1 0 2205 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-292
transform 1 0 2171 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-293
transform 1 0 2288 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-294
transform 1 0 2530 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-295
transform 1 0 2653 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-296
transform 1 0 2719 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-297
transform 1 0 2783 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-298
transform 1 0 2882 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-299
transform 1 0 2914 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-300
transform 1 0 2870 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-301
transform 1 0 2771 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-302
transform 1 0 2749 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-303
transform 1 0 2760 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-304
transform 1 0 2754 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-305
transform 1 0 2700 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-306
transform 1 0 2720 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-307
transform 1 0 2731 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-308
transform 1 0 2649 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-309
transform 1 0 2873 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-310
transform 1 0 2917 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-311
transform 1 0 2873 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-312
transform 1 0 2774 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-313
transform 1 0 2752 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-314
transform 1 0 2763 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-315
transform 1 0 2738 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-316
transform 1 0 2825 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-317
transform 1 0 2395 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-318
transform 1 0 2398 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-319
transform 1 0 2320 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-320
transform 1 0 2273 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-321
transform 1 0 2367 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-322
transform 1 0 2215 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-323
transform 1 0 2217 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-324
transform 1 0 2672 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-325
transform 1 0 2646 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-326
transform 1 0 2706 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-327
transform 1 0 2675 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-328
transform 1 0 2649 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-329
transform 1 0 2709 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-330
transform 1 0 2712 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-331
transform 1 0 2701 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-332
transform 1 0 2654 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-333
transform 1 0 2664 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-334
transform 1 0 2582 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-335
transform 1 0 2584 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-336
transform 1 0 2521 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-337
transform 1 0 2429 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-338
transform 1 0 2413 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-339
transform 1 0 2183 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-340
transform 1 0 2168 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-341
transform 1 0 2208 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-342
transform 1 0 2198 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-343
transform 1 0 2183 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-344
transform 1 0 2235 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-345
transform 1 0 2464 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-346
transform 1 0 2419 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-347
transform 1 0 2447 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-348
transform 1 0 2583 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-349
transform 1 0 2390 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-350
transform 1 0 2527 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-351
transform 1 0 2627 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-352
transform 1 0 2459 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-353
transform 1 0 2527 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-354
transform 1 0 2216 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-355
transform 1 0 2193 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-356
transform 1 0 2422 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-357
transform 1 0 2410 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-358
transform 1 0 2353 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-359
transform 1 0 2316 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-360
transform 1 0 2158 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-361
transform 1 0 2164 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-362
transform 1 0 2171 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-363
transform 1 0 2142 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-364
transform 1 0 2701 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-365
transform 1 0 2274 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-366
transform 1 0 2183 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-367
transform 1 0 2362 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-368
transform 1 0 2318 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-369
transform 1 0 2372 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-370
transform 1 0 2485 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-371
transform 1 0 2194 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-372
transform 1 0 2210 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-373
transform 1 0 2187 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-374
transform 1 0 2495 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-375
transform 1 0 2367 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-376
transform 1 0 2201 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-377
transform 1 0 2242 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-378
transform 1 0 2288 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-379
transform 1 0 2242 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-380
transform 1 0 2471 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-381
transform 1 0 2239 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-382
transform 1 0 2224 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-383
transform 1 0 2407 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-384
transform 1 0 2269 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-385
transform 1 0 2103 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-386
transform 1 0 2124 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-387
transform 1 0 2125 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-388
transform 1 0 2116 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-389
transform 1 0 2122 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-390
transform 1 0 2156 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-391
transform 1 0 2141 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-392
transform 1 0 2159 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-393
transform 1 0 2134 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-394
transform 1 0 2118 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-395
transform 1 0 2130 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-396
transform 1 0 2104 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-397
transform 1 0 2111 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-398
transform 1 0 2092 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-399
transform 1 0 2077 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-400
transform 1 0 2688 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-401
transform 1 0 2489 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-402
transform 1 0 2619 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-403
transform 1 0 2509 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-404
transform 1 0 2488 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-405
transform 1 0 2705 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-406
transform 1 0 2728 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-407
transform 1 0 2588 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-408
transform 1 0 2593 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-409
transform 1 0 2564 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-410
transform 1 0 2472 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-411
transform 1 0 2170 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-412
transform 1 0 2176 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-413
transform 1 0 2192 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-414
transform 1 0 2164 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-415
transform 1 0 2409 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-416
transform 1 0 2470 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-417
transform 1 0 2593 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-418
transform 1 0 2683 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-419
transform 1 0 2684 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-420
transform 1 0 2132 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-421
transform 1 0 2156 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-422
transform 1 0 2315 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-423
transform 1 0 2293 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-424
transform 1 0 2252 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-425
transform 1 0 2515 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-426
transform 1 0 2324 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-427
transform 1 0 2558 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-428
transform 1 0 2473 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-429
transform 1 0 2475 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-430
transform 1 0 2468 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-431
transform 1 0 2244 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-432
transform 1 0 2318 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-433
transform 1 0 2424 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-434
transform 1 0 2475 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-435
transform 1 0 2659 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-436
transform 1 0 2549 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-437
transform 1 0 2569 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-438
transform 1 0 2789 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-439
transform 1 0 2542 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-440
transform 1 0 2569 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-441
transform 1 0 2333 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-442
transform 1 0 2353 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-443
transform 1 0 2792 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-444
transform 1 0 2791 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-445
transform 1 0 2431 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-446
transform 1 0 2311 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-447
transform 1 0 2656 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-448
transform 1 0 2378 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-449
transform 1 0 2395 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-450
transform 1 0 2750 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-451
transform 1 0 2341 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-452
transform 1 0 2321 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-453
transform 1 0 2598 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-454
transform 1 0 2491 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-455
transform 1 0 2648 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-456
transform 1 0 2587 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-457
transform 1 0 2468 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-458
transform 1 0 2517 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-459
transform 1 0 2207 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-460
transform 1 0 2236 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-461
transform 1 0 2175 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-462
transform 1 0 2213 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-463
transform 1 0 2181 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-464
transform 1 0 2176 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-465
transform 1 0 2372 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-466
transform 1 0 2245 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-467
transform 1 0 2644 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-468
transform 1 0 2639 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-469
transform 1 0 2542 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-470
transform 1 0 2450 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-471
transform 1 0 2529 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-472
transform 1 0 2456 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-473
transform 1 0 2440 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-474
transform 1 0 2443 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-475
transform 1 0 2346 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-476
transform 1 0 2321 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-477
transform 1 0 2247 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-478
transform 1 0 2619 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-479
transform 1 0 2684 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-480
transform 1 0 2620 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-481
transform 1 0 2566 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-482
transform 1 0 2546 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-483
transform 1 0 2641 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-484
transform 1 0 2137 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-485
transform 1 0 2197 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-486
transform 1 0 2203 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-487
transform 1 0 2223 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-488
transform 1 0 2198 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-489
transform 1 0 2190 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-490
transform 1 0 2221 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-491
transform 1 0 2287 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-492
transform 1 0 2228 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-493
transform 1 0 2277 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-494
transform 1 0 2194 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-495
transform 1 0 2206 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-496
transform 1 0 2180 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-497
transform 1 0 2200 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-498
transform 1 0 2233 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-499
transform 1 0 2637 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-500
transform 1 0 2640 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-501
transform 1 0 2707 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-502
transform 1 0 2696 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-503
transform 1 0 2682 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-504
transform 1 0 2742 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-505
transform 1 0 2766 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-506
transform 1 0 2524 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-507
transform 1 0 2587 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-508
transform 1 0 2585 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-509
transform 1 0 2667 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-510
transform 1 0 2612 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-511
transform 1 0 2121 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-512
transform 1 0 2137 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-513
transform 1 0 2124 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-514
transform 1 0 2258 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-515
transform 1 0 2278 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-516
transform 1 0 2249 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-517
transform 1 0 2266 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-518
transform 1 0 2236 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-519
transform 1 0 2233 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-520
transform 1 0 2216 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-521
transform 1 0 2157 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-522
transform 1 0 2264 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-523
transform 1 0 2355 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-524
transform 1 0 2382 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-525
transform 1 0 2379 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-526
transform 1 0 2171 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-527
transform 1 0 2177 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-528
transform 1 0 2170 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-529
transform 1 0 2283 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-530
transform 1 0 2581 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-531
transform 1 0 2665 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-532
transform 1 0 2615 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-533
transform 1 0 2737 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-534
transform 1 0 2831 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-535
transform 1 0 2473 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-536
transform 1 0 2480 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-537
transform 1 0 2481 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-538
transform 1 0 2500 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-539
transform 1 0 2597 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-540
transform 1 0 2858 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-541
transform 1 0 2861 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-542
transform 1 0 2759 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-543
transform 1 0 2731 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-544
transform 1 0 2748 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-545
transform 1 0 2783 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-546
transform 1 0 2742 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-547
transform 1 0 2678 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-548
transform 1 0 2689 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-549
transform 1 0 2613 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-550
transform 1 0 2796 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-551
transform 1 0 2825 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-552
transform 1 0 2917 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-553
transform 1 0 2968 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-554
transform 1 0 2947 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-555
transform 1 0 2855 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-556
transform 1 0 2817 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-557
transform 1 0 2744 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-558
transform 1 0 2647 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-559
transform 1 0 2295 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-560
transform 1 0 2330 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-561
transform 1 0 2302 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-562
transform 1 0 2384 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-563
transform 1 0 2383 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-564
transform 1 0 2345 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-565
transform 1 0 2437 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-566
transform 1 0 2280 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-567
transform 1 0 2281 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-568
transform 1 0 2271 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-569
transform 1 0 2311 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-570
transform 1 0 2350 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-571
transform 1 0 2368 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-572
transform 1 0 2465 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-573
transform 1 0 2275 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-574
transform 1 0 2279 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-575
transform 1 0 2467 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-576
transform 1 0 2153 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-577
transform 1 0 2176 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-578
transform 1 0 2188 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-579
transform 1 0 2218 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-580
transform 1 0 2204 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-581
transform 1 0 2230 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-582
transform 1 0 2126 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-583
transform 1 0 2159 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-584
transform 1 0 2162 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-585
transform 1 0 2316 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-586
transform 1 0 2878 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-587
transform 1 0 2872 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-588
transform 1 0 2828 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-589
transform 1 0 2566 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-590
transform 1 0 2459 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-591
transform 1 0 2649 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-592
transform 1 0 2567 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-593
transform 1 0 2470 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-594
transform 1 0 2518 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-595
transform 1 0 2608 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-596
transform 1 0 2665 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-597
transform 1 0 2705 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-598
transform 1 0 2127 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-599
transform 1 0 2130 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-600
transform 1 0 2840 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-601
transform 1 0 2788 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-602
transform 1 0 2708 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-603
transform 1 0 2228 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-604
transform 1 0 2205 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-605
transform 1 0 2288 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-606
transform 1 0 2180 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-607
transform 1 0 2294 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-608
transform 1 0 2325 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-609
transform 1 0 2378 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-610
transform 1 0 2370 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-611
transform 1 0 2381 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-612
transform 1 0 2593 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-613
transform 1 0 2539 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-614
transform 1 0 2587 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-615
transform 1 0 2473 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-616
transform 1 0 2503 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-617
transform 1 0 2575 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-618
transform 1 0 2359 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-619
transform 1 0 2386 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-620
transform 1 0 2392 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-621
transform 1 0 2228 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-622
transform 1 0 2310 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-623
transform 1 0 2221 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-624
transform 1 0 2203 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-625
transform 1 0 2218 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-626
transform 1 0 2200 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-627
transform 1 0 2642 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-628
transform 1 0 2704 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-629
transform 1 0 2687 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-630
transform 1 0 2566 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-631
transform 1 0 2783 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-632
transform 1 0 2642 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-633
transform 1 0 2622 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-634
transform 1 0 2647 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-635
transform 1 0 2642 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-636
transform 1 0 2738 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-637
transform 1 0 2836 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-638
transform 1 0 2587 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-639
transform 1 0 2747 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-640
transform 1 0 2638 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-641
transform 1 0 2590 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-642
transform 1 0 2527 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-643
transform 1 0 2453 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-644
transform 1 0 2447 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-645
transform 1 0 2490 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-646
transform 1 0 2509 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-647
transform 1 0 2566 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-648
transform 1 0 2628 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-649
transform 1 0 2169 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-650
transform 1 0 2187 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-651
transform 1 0 2251 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-652
transform 1 0 2643 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-653
transform 1 0 2690 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-654
transform 1 0 2843 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-655
transform 1 0 2194 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-656
transform 1 0 2195 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-657
transform 1 0 2366 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-658
transform 1 0 2444 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-659
transform 1 0 2369 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-660
transform 1 0 2385 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-661
transform 1 0 2107 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-662
transform 1 0 2119 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-663
transform 1 0 2153 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-664
transform 1 0 2113 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-665
transform 1 0 2122 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-666
transform 1 0 2264 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-667
transform 1 0 2349 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-668
transform 1 0 2446 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-669
transform 1 0 2676 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-670
transform 1 0 2682 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-671
transform 1 0 2278 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-672
transform 1 0 2284 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-673
transform 1 0 2237 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-674
transform 1 0 2319 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-675
transform 1 0 2261 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-676
transform 1 0 2353 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-677
transform 1 0 2492 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-678
transform 1 0 2263 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-679
transform 1 0 2384 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-680
transform 1 0 2389 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-681
transform 1 0 2744 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-682
transform 1 0 2356 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-683
transform 1 0 2540 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-684
transform 1 0 2485 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-685
transform 1 0 2294 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-686
transform 1 0 2460 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-687
transform 1 0 2348 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-688
transform 1 0 2329 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-689
transform 1 0 2260 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-690
transform 1 0 2220 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-691
transform 1 0 2257 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-692
transform 1 0 2405 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-693
transform 1 0 2271 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-694
transform 1 0 2240 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-695
transform 1 0 2431 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-696
transform 1 0 2433 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-697
transform 1 0 2233 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-698
transform 1 0 2223 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-699
transform 1 0 2354 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-700
transform 1 0 2596 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-701
transform 1 0 2444 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-702
transform 1 0 2545 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-703
transform 1 0 2291 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-704
transform 1 0 2278 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-705
transform 1 0 2243 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-706
transform 1 0 2217 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-707
transform 1 0 2706 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-708
transform 1 0 2689 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-709
transform 1 0 2700 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-710
transform 1 0 2683 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-711
transform 1 0 2645 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-712
transform 1 0 2622 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-713
transform 1 0 2657 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-714
transform 1 0 2225 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-715
transform 1 0 2226 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-716
transform 1 0 2215 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-717
transform 1 0 2193 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-718
transform 1 0 2205 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-719
transform 1 0 2262 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-720
transform 1 0 2314 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-721
transform 1 0 2359 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-722
transform 1 0 2194 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-723
transform 1 0 2674 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-724
transform 1 0 2694 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-725
transform 1 0 2757 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-726
transform 1 0 2703 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-727
transform 1 0 2514 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-728
transform 1 0 2636 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-729
transform 1 0 2577 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-730
transform 1 0 2573 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-731
transform 1 0 2272 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-732
transform 1 0 2263 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-733
transform 1 0 2269 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-734
transform 1 0 2255 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-735
transform 1 0 2323 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-736
transform 1 0 2327 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-737
transform 1 0 2290 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-738
transform 1 0 2261 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-739
transform 1 0 2278 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-740
transform 1 0 2302 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-741
transform 1 0 2279 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-742
transform 1 0 2494 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-743
transform 1 0 2296 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-744
transform 1 0 2158 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-745
transform 1 0 2197 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-746
transform 1 0 2211 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-747
transform 1 0 2295 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-748
transform 1 0 2362 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-749
transform 1 0 2413 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-750
transform 1 0 2173 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-751
transform 1 0 2217 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-752
transform 1 0 2334 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-753
transform 1 0 2380 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-754
transform 1 0 2431 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-755
transform 1 0 2551 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-756
transform 1 0 2351 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-757
transform 1 0 2407 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-758
transform 1 0 2603 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-759
transform 1 0 2365 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-760
transform 1 0 2136 0 1 1010
box 0 0 3 6
use FEEDTHRU  F-761
transform 1 0 2182 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-762
transform 1 0 2244 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-763
transform 1 0 2280 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-764
transform 1 0 2240 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-765
transform 1 0 2479 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-766
transform 1 0 2522 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-767
transform 1 0 2329 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-768
transform 1 0 2346 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-769
transform 1 0 2363 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-770
transform 1 0 2419 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-771
transform 1 0 2714 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-772
transform 1 0 2435 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-773
transform 1 0 2415 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-774
transform 1 0 2349 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-775
transform 1 0 2604 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-776
transform 1 0 2549 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-777
transform 1 0 2572 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-778
transform 1 0 2603 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-779
transform 1 0 2638 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-780
transform 1 0 2592 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-781
transform 1 0 2504 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-782
transform 1 0 2512 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-783
transform 1 0 2131 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-784
transform 1 0 2169 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-785
transform 1 0 2210 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-786
transform 1 0 2239 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-787
transform 1 0 2220 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-788
transform 1 0 2195 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-789
transform 1 0 2545 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-790
transform 1 0 2389 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-791
transform 1 0 2458 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-792
transform 1 0 2462 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-793
transform 1 0 2538 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-794
transform 1 0 2453 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-795
transform 1 0 2533 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-796
transform 1 0 2585 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-797
transform 1 0 2733 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-798
transform 1 0 2733 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-799
transform 1 0 2609 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-800
transform 1 0 2667 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-801
transform 1 0 2561 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-802
transform 1 0 2598 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-803
transform 1 0 2522 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-804
transform 1 0 2528 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-805
transform 1 0 2711 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-806
transform 1 0 2356 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-807
transform 1 0 2450 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-808
transform 1 0 2303 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-809
transform 1 0 2340 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-810
transform 1 0 2258 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-811
transform 1 0 2453 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-812
transform 1 0 2278 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-813
transform 1 0 2292 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-814
transform 1 0 2327 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-815
transform 1 0 2210 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-816
transform 1 0 2358 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-817
transform 1 0 2373 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-818
transform 1 0 2416 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-819
transform 1 0 2432 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-820
transform 1 0 2407 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-821
transform 1 0 2476 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-822
transform 1 0 2468 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-823
transform 1 0 2550 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-824
transform 1 0 2543 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-825
transform 1 0 2536 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-826
transform 1 0 2570 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-827
transform 1 0 2590 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-828
transform 1 0 2601 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-829
transform 1 0 2324 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-830
transform 1 0 2340 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-831
transform 1 0 2680 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-832
transform 1 0 2769 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-833
transform 1 0 2745 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-834
transform 1 0 2603 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-835
transform 1 0 2681 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-836
transform 1 0 2692 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-837
transform 1 0 2616 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-838
transform 1 0 2572 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-839
transform 1 0 2221 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-840
transform 1 0 2605 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-841
transform 1 0 2524 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-842
transform 1 0 2463 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-843
transform 1 0 2361 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-844
transform 1 0 2756 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-845
transform 1 0 2266 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-846
transform 1 0 2270 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-847
transform 1 0 2260 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-848
transform 1 0 2260 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-849
transform 1 0 2251 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-850
transform 1 0 2234 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-851
transform 1 0 2272 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-852
transform 1 0 2276 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-853
transform 1 0 2266 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-854
transform 1 0 2231 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-855
transform 1 0 2361 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-856
transform 1 0 2389 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-857
transform 1 0 2259 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-858
transform 1 0 2326 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-859
transform 1 0 2443 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-860
transform 1 0 2459 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-861
transform 1 0 2393 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-862
transform 1 0 2296 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-863
transform 1 0 2321 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-864
transform 1 0 2391 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-865
transform 1 0 2206 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-866
transform 1 0 2660 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-867
transform 1 0 2443 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-868
transform 1 0 2483 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-869
transform 1 0 2557 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-870
transform 1 0 2491 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-871
transform 1 0 2428 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-872
transform 1 0 2369 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-873
transform 1 0 2340 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-874
transform 1 0 2323 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-875
transform 1 0 2621 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-876
transform 1 0 2434 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-877
transform 1 0 2365 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-878
transform 1 0 2371 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-879
transform 1 0 2321 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-880
transform 1 0 2365 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-881
transform 1 0 2588 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-882
transform 1 0 2545 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-883
transform 1 0 2574 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-884
transform 1 0 2633 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-885
transform 1 0 2656 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-886
transform 1 0 2759 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-887
transform 1 0 2794 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-888
transform 1 0 2633 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-889
transform 1 0 2623 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-890
transform 1 0 2542 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-891
transform 1 0 2571 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-892
transform 1 0 2630 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-893
transform 1 0 2653 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-894
transform 1 0 2534 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-895
transform 1 0 2554 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-896
transform 1 0 2134 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-897
transform 1 0 2157 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-898
transform 1 0 2168 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-899
transform 1 0 2304 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-900
transform 1 0 2357 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-901
transform 1 0 2269 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-902
transform 1 0 2264 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-903
transform 1 0 2407 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-904
transform 1 0 2192 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-905
transform 1 0 2334 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-906
transform 1 0 2333 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-907
transform 1 0 2307 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-908
transform 1 0 2215 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-909
transform 1 0 2219 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-910
transform 1 0 2214 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-911
transform 1 0 2219 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-912
transform 1 0 2263 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-913
transform 1 0 2283 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-914
transform 1 0 2251 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-915
transform 1 0 2219 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-916
transform 1 0 2175 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-917
transform 1 0 2128 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-918
transform 1 0 2257 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-919
transform 1 0 2281 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-920
transform 1 0 2290 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-921
transform 1 0 2267 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-922
transform 1 0 2311 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-923
transform 1 0 2303 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-924
transform 1 0 2317 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-925
transform 1 0 2270 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-926
transform 1 0 2263 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-927
transform 1 0 2287 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-928
transform 1 0 2296 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-929
transform 1 0 2273 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-930
transform 1 0 2317 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-931
transform 1 0 2315 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-932
transform 1 0 2323 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-933
transform 1 0 2276 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-934
transform 1 0 2720 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-935
transform 1 0 2818 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-936
transform 1 0 2810 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-937
transform 1 0 2794 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-938
transform 1 0 2528 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-939
transform 1 0 2771 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-940
transform 1 0 2204 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-941
transform 1 0 2174 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-942
transform 1 0 2166 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-943
transform 1 0 2178 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-944
transform 1 0 2227 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-945
transform 1 0 2201 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-946
transform 1 0 2337 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-947
transform 1 0 2345 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-948
transform 1 0 2251 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-949
transform 1 0 2222 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-950
transform 1 0 2257 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-951
transform 1 0 2268 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-952
transform 1 0 2309 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-953
transform 1 0 2359 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-954
transform 1 0 2339 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-955
transform 1 0 2341 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-956
transform 1 0 2291 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-957
transform 1 0 2314 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-958
transform 1 0 2405 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-959
transform 1 0 2382 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-960
transform 1 0 2350 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-961
transform 1 0 2456 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-962
transform 1 0 2371 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-963
transform 1 0 2318 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-964
transform 1 0 2358 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-965
transform 1 0 2276 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-966
transform 1 0 2323 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-967
transform 1 0 2563 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-968
transform 1 0 2491 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-969
transform 1 0 2647 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-970
transform 1 0 2695 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-971
transform 1 0 2759 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-972
transform 1 0 2876 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-973
transform 1 0 2822 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-974
transform 1 0 2800 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-975
transform 1 0 2566 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-976
transform 1 0 2650 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-977
transform 1 0 2698 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-978
transform 1 0 2726 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-979
transform 1 0 2824 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-980
transform 1 0 2816 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-981
transform 1 0 2187 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-982
transform 1 0 2180 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-983
transform 1 0 2179 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-984
transform 1 0 2237 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-985
transform 1 0 2371 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-986
transform 1 0 2373 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-987
transform 1 0 2155 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-988
transform 1 0 2625 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-989
transform 1 0 2400 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-990
transform 1 0 2585 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-991
transform 1 0 2413 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-992
transform 1 0 2600 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-993
transform 1 0 2503 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-994
transform 1 0 2421 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-995
transform 1 0 2477 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-996
transform 1 0 2509 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-997
transform 1 0 2708 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-998
transform 1 0 2536 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-999
transform 1 0 2498 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1000
transform 1 0 2626 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1001
transform 1 0 2660 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1002
transform 1 0 2625 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1003
transform 1 0 2631 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1004
transform 1 0 2672 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1005
transform 1 0 2797 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1006
transform 1 0 2813 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1007
transform 1 0 2821 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1008
transform 1 0 2723 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1009
transform 1 0 2677 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1010
transform 1 0 2632 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1011
transform 1 0 2548 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1012
transform 1 0 2219 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1013
transform 1 0 2377 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1014
transform 1 0 2403 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1015
transform 1 0 2478 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1016
transform 1 0 2628 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1017
transform 1 0 2716 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1018
transform 1 0 2701 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1019
transform 1 0 2586 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1020
transform 1 0 2391 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1021
transform 1 0 2473 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1022
transform 1 0 2530 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1023
transform 1 0 2510 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1024
transform 1 0 2467 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1025
transform 1 0 2282 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1026
transform 1 0 2278 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1027
transform 1 0 2232 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1028
transform 1 0 2243 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1029
transform 1 0 2307 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1030
transform 1 0 2258 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-1031
transform 1 0 2156 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-1032
transform 1 0 2543 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1033
transform 1 0 2394 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1034
transform 1 0 2330 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1035
transform 1 0 2416 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1036
transform 1 0 2504 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1037
transform 1 0 2362 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1038
transform 1 0 2436 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1039
transform 1 0 2423 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1040
transform 1 0 2488 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1041
transform 1 0 2684 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1042
transform 1 0 2470 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1043
transform 1 0 2426 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1044
transform 1 0 2202 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1045
transform 1 0 2156 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1046
transform 1 0 2198 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1047
transform 1 0 2194 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1048
transform 1 0 2370 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1049
transform 1 0 2337 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1050
transform 1 0 2340 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1051
transform 1 0 2427 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1052
transform 1 0 2488 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1053
transform 1 0 2575 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1054
transform 1 0 2626 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1055
transform 1 0 2223 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-1056
transform 1 0 2322 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1057
transform 1 0 2430 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1058
transform 1 0 2491 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1059
transform 1 0 2578 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1060
transform 1 0 2599 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1061
transform 1 0 2636 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1062
transform 1 0 2665 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1063
transform 1 0 2762 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1064
transform 1 0 2383 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1065
transform 1 0 2375 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1066
transform 1 0 2335 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1067
transform 1 0 2285 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1068
transform 1 0 2262 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1069
transform 1 0 2220 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1070
transform 1 0 2207 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1071
transform 1 0 2203 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1072
transform 1 0 2189 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1073
transform 1 0 2227 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1074
transform 1 0 2409 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1075
transform 1 0 2282 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1076
transform 1 0 2329 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1077
transform 1 0 2309 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1078
transform 1 0 2305 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1079
transform 1 0 2261 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1080
transform 1 0 2284 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1081
transform 1 0 2356 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1082
transform 1 0 2347 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1083
transform 1 0 2277 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1084
transform 1 0 2160 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1085
transform 1 0 2119 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-1086
transform 1 0 2226 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1087
transform 1 0 2213 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1088
transform 1 0 2209 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1089
transform 1 0 2198 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1090
transform 1 0 2232 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1091
transform 1 0 2165 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1092
transform 1 0 2461 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1093
transform 1 0 2485 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1094
transform 1 0 2170 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-1095
transform 1 0 2241 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1096
transform 1 0 2331 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1097
transform 1 0 2374 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1098
transform 1 0 2443 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1099
transform 1 0 2485 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1100
transform 1 0 2189 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1101
transform 1 0 2251 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1102
transform 1 0 2303 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1103
transform 1 0 2353 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1104
transform 1 0 2333 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1105
transform 1 0 2329 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1106
transform 1 0 2337 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1107
transform 1 0 2342 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1108
transform 1 0 2500 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1109
transform 1 0 2354 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1110
transform 1 0 2449 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1111
transform 1 0 2201 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1112
transform 1 0 2230 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1113
transform 1 0 2370 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1114
transform 1 0 2485 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1115
transform 1 0 2545 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1116
transform 1 0 2626 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1117
transform 1 0 2674 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1118
transform 1 0 2702 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1119
transform 1 0 2803 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1120
transform 1 0 2795 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1121
transform 1 0 2782 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1122
transform 1 0 2678 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1123
transform 1 0 2637 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1124
transform 1 0 2632 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1125
transform 1 0 2582 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1126
transform 1 0 2691 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1127
transform 1 0 2579 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1128
transform 1 0 2568 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1129
transform 1 0 2498 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1130
transform 1 0 2518 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1131
transform 1 0 2455 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1132
transform 1 0 2376 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1133
transform 1 0 2371 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1134
transform 1 0 2363 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1135
transform 1 0 2347 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1136
transform 1 0 2297 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1137
transform 1 0 2284 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1138
transform 1 0 2342 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1139
transform 1 0 2272 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1140
transform 1 0 2270 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1141
transform 1 0 2304 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1142
transform 1 0 2290 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1143
transform 1 0 2310 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1144
transform 1 0 2296 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1145
transform 1 0 2294 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1146
transform 1 0 2302 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1147
transform 1 0 2333 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1148
transform 1 0 2328 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1149
transform 1 0 2311 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1150
transform 1 0 2318 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1151
transform 1 0 2320 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1152
transform 1 0 2276 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1153
transform 1 0 2295 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1154
transform 1 0 2401 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1155
transform 1 0 2345 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1156
transform 1 0 2393 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1157
transform 1 0 2371 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1158
transform 1 0 2327 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1159
transform 1 0 2401 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1160
transform 1 0 2389 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1161
transform 1 0 2332 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1162
transform 1 0 2358 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1163
transform 1 0 2431 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1164
transform 1 0 2494 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1165
transform 1 0 2434 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1166
transform 1 0 2497 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1167
transform 1 0 2419 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1168
transform 1 0 2482 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1169
transform 1 0 2474 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1170
transform 1 0 2544 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1171
transform 1 0 2629 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1172
transform 1 0 2339 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1173
transform 1 0 2355 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1174
transform 1 0 2477 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1175
transform 1 0 2401 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1176
transform 1 0 2600 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1177
transform 1 0 2574 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1178
transform 1 0 2224 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1179
transform 1 0 2241 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1180
transform 1 0 2267 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1181
transform 1 0 2314 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1182
transform 1 0 2294 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1183
transform 1 0 2290 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1184
transform 1 0 2240 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1185
transform 1 0 2257 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1186
transform 1 0 2242 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1187
transform 1 0 2224 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1188
transform 1 0 2177 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1189
transform 1 0 2312 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1190
transform 1 0 2302 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1191
transform 1 0 2316 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1192
transform 1 0 2357 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1193
transform 1 0 2407 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1194
transform 1 0 2741 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1195
transform 1 0 2839 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1196
transform 1 0 2666 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1197
transform 1 0 2761 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1198
transform 1 0 2756 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1199
transform 1 0 2635 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1200
transform 1 0 2660 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1201
transform 1 0 2755 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1202
transform 1 0 2638 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1203
transform 1 0 2648 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1204
transform 1 0 2749 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1205
transform 1 0 2261 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-1206
transform 1 0 2238 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1207
transform 1 0 2328 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1208
transform 1 0 2155 0 1 5786
box 0 0 3 6
use FEEDTHRU  F-1209
transform 1 0 2200 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-1210
transform 1 0 2506 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1211
transform 1 0 2510 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1212
transform 1 0 2491 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1213
transform 1 0 2612 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1214
transform 1 0 2822 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1215
transform 1 0 2887 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1216
transform 1 0 2864 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1217
transform 1 0 2635 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1218
transform 1 0 2640 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1219
transform 1 0 2681 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1220
transform 1 0 2785 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1221
transform 1 0 2479 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1222
transform 1 0 2523 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1223
transform 1 0 2567 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1224
transform 1 0 2395 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1225
transform 1 0 2369 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1226
transform 1 0 2359 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1227
transform 1 0 2315 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1228
transform 1 0 2329 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1229
transform 1 0 2329 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1230
transform 1 0 2296 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1231
transform 1 0 2256 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1232
transform 1 0 2235 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1233
transform 1 0 2146 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-1234
transform 1 0 2239 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1235
transform 1 0 2243 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1236
transform 1 0 2253 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1237
transform 1 0 2439 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1238
transform 1 0 2533 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1239
transform 1 0 2656 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1240
transform 1 0 2722 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1241
transform 1 0 2627 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1242
transform 1 0 2683 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1243
transform 1 0 2899 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1244
transform 1 0 2647 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1245
transform 1 0 2579 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1246
transform 1 0 2553 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1247
transform 1 0 2334 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1248
transform 1 0 2442 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1249
transform 1 0 2494 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1250
transform 1 0 2563 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1251
transform 1 0 2392 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1252
transform 1 0 2340 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1253
transform 1 0 2253 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1254
transform 1 0 2494 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1255
transform 1 0 2560 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1256
transform 1 0 2363 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1257
transform 1 0 2413 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1258
transform 1 0 2537 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1259
transform 1 0 2462 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1260
transform 1 0 2569 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1261
transform 1 0 2486 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1262
transform 1 0 2611 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1263
transform 1 0 2496 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1264
transform 1 0 2426 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1265
transform 1 0 2455 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1266
transform 1 0 2489 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1267
transform 1 0 2440 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1268
transform 1 0 2490 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1269
transform 1 0 2432 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1270
transform 1 0 2436 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1271
transform 1 0 2354 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1272
transform 1 0 2377 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1273
transform 1 0 2308 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1274
transform 1 0 2482 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1275
transform 1 0 2542 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1276
transform 1 0 2611 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1277
transform 1 0 2653 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1278
transform 1 0 2678 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1279
transform 1 0 2767 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1280
transform 1 0 2771 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1281
transform 1 0 2776 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1282
transform 1 0 2762 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1283
transform 1 0 2734 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1284
transform 1 0 2751 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1285
transform 1 0 2552 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1286
transform 1 0 2548 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1287
transform 1 0 2594 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1288
transform 1 0 2562 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1289
transform 1 0 2492 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1290
transform 1 0 2575 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1291
transform 1 0 2437 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1292
transform 1 0 2382 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1293
transform 1 0 2384 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1294
transform 1 0 2280 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1295
transform 1 0 2358 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1296
transform 1 0 2416 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1297
transform 1 0 2485 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1298
transform 1 0 2530 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1299
transform 1 0 2369 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1300
transform 1 0 2428 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1301
transform 1 0 2591 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1302
transform 1 0 2191 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-1303
transform 1 0 2118 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1304
transform 1 0 2482 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1305
transform 1 0 2501 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1306
transform 1 0 2163 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1307
transform 1 0 2265 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1308
transform 1 0 2437 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1309
transform 1 0 2462 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1310
transform 1 0 2277 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1311
transform 1 0 2184 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1312
transform 1 0 2248 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1313
transform 1 0 2581 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1314
transform 1 0 2558 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1315
transform 1 0 2554 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1316
transform 1 0 2702 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1317
transform 1 0 2569 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1318
transform 1 0 2301 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1319
transform 1 0 2419 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1320
transform 1 0 2507 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1321
transform 1 0 2322 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1322
transform 1 0 2351 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1323
transform 1 0 2413 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1324
transform 1 0 2399 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1325
transform 1 0 2371 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1326
transform 1 0 2434 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1327
transform 1 0 2432 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1328
transform 1 0 2496 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1329
transform 1 0 2354 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1330
transform 1 0 2181 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1331
transform 1 0 2187 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1332
transform 1 0 2695 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1333
transform 1 0 2675 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1334
transform 1 0 2683 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1335
transform 1 0 2732 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1336
transform 1 0 2728 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1337
transform 1 0 2227 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-1338
transform 1 0 2253 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1339
transform 1 0 2222 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1340
transform 1 0 2214 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1341
transform 1 0 2254 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1342
transform 1 0 2317 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1343
transform 1 0 2264 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1344
transform 1 0 2364 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1345
transform 1 0 2233 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1346
transform 1 0 2247 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1347
transform 1 0 2275 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1348
transform 1 0 2326 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1349
transform 1 0 2244 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1350
transform 1 0 2440 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1351
transform 1 0 2446 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1352
transform 1 0 2447 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1353
transform 1 0 2452 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1354
transform 1 0 2378 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1355
transform 1 0 2364 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1356
transform 1 0 2504 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1357
transform 1 0 2499 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1358
transform 1 0 2435 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1359
transform 1 0 2437 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1360
transform 1 0 2374 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1361
transform 1 0 2484 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1362
transform 1 0 2327 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1363
transform 1 0 2409 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1364
transform 1 0 2377 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1365
transform 1 0 2337 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1366
transform 1 0 2339 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1367
transform 1 0 2210 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1368
transform 1 0 2205 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1369
transform 1 0 2245 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1370
transform 1 0 2302 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1371
transform 1 0 2252 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1372
transform 1 0 2346 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1373
transform 1 0 2336 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1374
transform 1 0 2350 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1375
transform 1 0 2207 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1376
transform 1 0 2202 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1377
transform 1 0 2242 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1378
transform 1 0 2299 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1379
transform 1 0 2249 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1380
transform 1 0 2454 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1381
transform 1 0 2429 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1382
transform 1 0 2515 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1383
transform 1 0 2478 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1384
transform 1 0 2422 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1385
transform 1 0 2402 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1386
transform 1 0 2395 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1387
transform 1 0 2408 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1388
transform 1 0 2388 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1389
transform 1 0 2294 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1390
transform 1 0 2447 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1391
transform 1 0 2521 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1392
transform 1 0 2597 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1393
transform 1 0 2512 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1394
transform 1 0 2474 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1395
transform 1 0 2563 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1396
transform 1 0 2305 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1397
transform 1 0 2495 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1398
transform 1 0 2849 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1399
transform 1 0 2788 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1400
transform 1 0 2510 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1401
transform 1 0 2267 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1402
transform 1 0 2233 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1403
transform 1 0 2195 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1404
transform 1 0 2266 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1405
transform 1 0 2285 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1406
transform 1 0 2278 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1407
transform 1 0 2375 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1408
transform 1 0 2307 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1409
transform 1 0 2308 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1410
transform 1 0 2255 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1411
transform 1 0 2284 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1412
transform 1 0 2366 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1413
transform 1 0 2365 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1414
transform 1 0 2410 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1415
transform 1 0 2360 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1416
transform 1 0 2359 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1417
transform 1 0 2378 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1418
transform 1 0 2448 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1419
transform 1 0 2317 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1420
transform 1 0 2320 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1421
transform 1 0 2309 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1422
transform 1 0 2290 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1423
transform 1 0 2452 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1424
transform 1 0 2477 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1425
transform 1 0 2511 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1426
transform 1 0 2507 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1427
transform 1 0 2516 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1428
transform 1 0 2456 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1429
transform 1 0 2408 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1430
transform 1 0 2346 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1431
transform 1 0 2312 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1432
transform 1 0 2608 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1433
transform 1 0 2654 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1434
transform 1 0 2611 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1435
transform 1 0 2555 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1436
transform 1 0 2710 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1437
transform 1 0 2494 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1438
transform 1 0 2438 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1439
transform 1 0 2771 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1440
transform 1 0 2620 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1441
transform 1 0 2648 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1442
transform 1 0 2629 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1443
transform 1 0 2507 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1444
transform 1 0 2502 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1445
transform 1 0 2579 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1446
transform 1 0 2632 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1447
transform 1 0 2630 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1448
transform 1 0 2179 0 1 1053
box 0 0 3 6
use FEEDTHRU  F-1449
transform 1 0 2277 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1450
transform 1 0 2352 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1451
transform 1 0 2545 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1452
transform 1 0 2629 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1453
transform 1 0 2634 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1454
transform 1 0 2680 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1455
transform 1 0 2384 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1456
transform 1 0 2461 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1457
transform 1 0 2437 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1458
transform 1 0 2402 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1459
transform 1 0 2452 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1460
transform 1 0 2435 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1461
transform 1 0 2584 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1462
transform 1 0 2444 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1463
transform 1 0 2427 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1464
transform 1 0 2395 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1465
transform 1 0 2330 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1466
transform 1 0 2471 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1467
transform 1 0 2557 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1468
transform 1 0 2543 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1469
transform 1 0 2567 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1470
transform 1 0 2509 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1471
transform 1 0 2512 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1472
transform 1 0 2498 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1473
transform 1 0 2602 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1474
transform 1 0 2589 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1475
transform 1 0 2473 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1476
transform 1 0 2392 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1477
transform 1 0 2333 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1478
transform 1 0 2672 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1479
transform 1 0 2710 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1480
transform 1 0 2666 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1481
transform 1 0 2408 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1482
transform 1 0 2443 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1483
transform 1 0 2425 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1484
transform 1 0 2357 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1485
transform 1 0 2377 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1486
transform 1 0 2389 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1487
transform 1 0 2453 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1488
transform 1 0 2501 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1489
transform 1 0 2506 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1490
transform 1 0 2495 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1491
transform 1 0 2236 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-1492
transform 1 0 2377 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-1493
transform 1 0 2358 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1494
transform 1 0 2309 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-1495
transform 1 0 2420 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1496
transform 1 0 2312 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1497
transform 1 0 2289 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1498
transform 1 0 2696 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1499
transform 1 0 2699 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1500
transform 1 0 2551 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1501
transform 1 0 2453 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1502
transform 1 0 2460 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1503
transform 1 0 2434 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1504
transform 1 0 2342 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1505
transform 1 0 2334 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1506
transform 1 0 2314 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1507
transform 1 0 2288 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1508
transform 1 0 2250 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1509
transform 1 0 2464 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1510
transform 1 0 2271 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1511
transform 1 0 2234 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1512
transform 1 0 2404 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1513
transform 1 0 2455 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1514
transform 1 0 2467 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1515
transform 1 0 2438 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1516
transform 1 0 2192 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1517
transform 1 0 2242 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1518
transform 1 0 2482 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1519
transform 1 0 2390 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1520
transform 1 0 2388 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1521
transform 1 0 2476 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1522
transform 1 0 2468 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1523
transform 1 0 2488 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1524
transform 1 0 2471 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1525
transform 1 0 2533 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1526
transform 1 0 2330 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1527
transform 1 0 2371 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1528
transform 1 0 2302 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1529
transform 1 0 2253 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1530
transform 1 0 2285 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1531
transform 1 0 2295 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1532
transform 1 0 2297 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-1533
transform 1 0 2183 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-1534
transform 1 0 2358 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1535
transform 1 0 2344 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1536
transform 1 0 2464 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1537
transform 1 0 2266 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1538
transform 1 0 2228 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1539
transform 1 0 2338 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1540
transform 1 0 2352 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1541
transform 1 0 2375 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1542
transform 1 0 2425 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1543
transform 1 0 2390 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1544
transform 1 0 2476 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1545
transform 1 0 2746 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1546
transform 1 0 2678 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1547
transform 1 0 2597 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1548
transform 1 0 2636 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1549
transform 1 0 2701 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1550
transform 1 0 2384 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1551
transform 1 0 2407 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1552
transform 1 0 2344 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1553
transform 1 0 2301 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1554
transform 1 0 2498 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1555
transform 1 0 2425 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1556
transform 1 0 2420 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1557
transform 1 0 2326 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1558
transform 1 0 2289 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1559
transform 1 0 2479 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1560
transform 1 0 2480 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1561
transform 1 0 2530 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1562
transform 1 0 2489 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1563
transform 1 0 2545 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1564
transform 1 0 2459 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1565
transform 1 0 2466 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1566
transform 1 0 2452 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1567
transform 1 0 2689 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1568
transform 1 0 2615 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1569
transform 1 0 2710 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1570
transform 1 0 2440 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1571
transform 1 0 2464 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1572
transform 1 0 2450 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1573
transform 1 0 2532 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1574
transform 1 0 2573 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1575
transform 1 0 2497 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1576
transform 1 0 2480 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1577
transform 1 0 2239 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1578
transform 1 0 2218 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1579
transform 1 0 2160 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1580
transform 1 0 2268 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1581
transform 1 0 2308 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1582
transform 1 0 2347 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1583
transform 1 0 2353 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1584
transform 1 0 2489 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1585
transform 1 0 2734 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1586
transform 1 0 2519 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1587
transform 1 0 2572 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1588
transform 1 0 2522 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1589
transform 1 0 2545 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1590
transform 1 0 2527 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1591
transform 1 0 2464 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1592
transform 1 0 2403 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1593
transform 1 0 2605 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1594
transform 1 0 2531 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1595
transform 1 0 2578 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1596
transform 1 0 2528 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1597
transform 1 0 2536 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1598
transform 1 0 2521 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1599
transform 1 0 2295 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1600
transform 1 0 2330 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1601
transform 1 0 2321 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-1602
transform 1 0 2324 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1603
transform 1 0 2361 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1604
transform 1 0 2365 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1605
transform 1 0 2428 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1606
transform 1 0 2414 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1607
transform 1 0 2502 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1608
transform 1 0 2537 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1609
transform 1 0 2461 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1610
transform 1 0 2396 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1611
transform 1 0 2464 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1612
transform 1 0 2519 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1613
transform 1 0 2449 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1614
transform 1 0 2525 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1615
transform 1 0 2722 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1616
transform 1 0 2396 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1617
transform 1 0 2681 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1618
transform 1 0 2770 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1619
transform 1 0 2774 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1620
transform 1 0 2737 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1621
transform 1 0 2743 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1622
transform 1 0 2603 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1623
transform 1 0 2204 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1624
transform 1 0 2254 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1625
transform 1 0 2800 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1626
transform 1 0 2543 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1627
transform 1 0 2512 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1628
transform 1 0 2224 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1629
transform 1 0 2541 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1630
transform 1 0 2465 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1631
transform 1 0 2195 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-1632
transform 1 0 2282 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-1633
transform 1 0 2337 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1634
transform 1 0 2276 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1635
transform 1 0 2265 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1636
transform 1 0 2614 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1637
transform 1 0 2552 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1638
transform 1 0 2524 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1639
transform 1 0 2515 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1640
transform 1 0 2458 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1641
transform 1 0 2397 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1642
transform 1 0 2310 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1643
transform 1 0 2323 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1644
transform 1 0 2326 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1645
transform 1 0 2390 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1646
transform 1 0 2458 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1647
transform 1 0 2381 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1648
transform 1 0 2494 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1649
transform 1 0 2374 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1650
transform 1 0 2400 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1651
transform 1 0 2396 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1652
transform 1 0 2527 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1653
transform 1 0 2405 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1654
transform 1 0 2500 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1655
transform 1 0 2617 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1656
transform 1 0 2786 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1657
transform 1 0 2596 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1658
transform 1 0 2540 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1659
transform 1 0 2515 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1660
transform 1 0 2497 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1661
transform 1 0 2602 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1662
transform 1 0 2328 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1663
transform 1 0 2383 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1664
transform 1 0 2557 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1665
transform 1 0 2537 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1666
transform 1 0 2508 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1667
transform 1 0 2570 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1668
transform 1 0 2473 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1669
transform 1 0 2501 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1670
transform 1 0 2605 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1671
transform 1 0 2592 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1672
transform 1 0 2609 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1673
transform 1 0 2749 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1674
transform 1 0 2627 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1675
transform 1 0 2707 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1676
transform 1 0 2639 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1677
transform 1 0 2428 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1678
transform 1 0 2501 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1679
transform 1 0 2454 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1680
transform 1 0 2366 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1681
transform 1 0 2401 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1682
transform 1 0 2423 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1683
transform 1 0 2527 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1684
transform 1 0 2520 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1685
transform 1 0 2711 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1686
transform 1 0 2791 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1687
transform 1 0 2843 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1688
transform 1 0 2638 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1689
transform 1 0 2576 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1690
transform 1 0 2542 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1691
transform 1 0 2608 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1692
transform 1 0 2527 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1693
transform 1 0 2466 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1694
transform 1 0 2524 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1695
transform 1 0 2372 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1696
transform 1 0 2308 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1697
transform 1 0 2276 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1698
transform 1 0 2698 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1699
transform 1 0 2342 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1700
transform 1 0 2483 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1701
transform 1 0 2418 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1702
transform 1 0 2423 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1703
transform 1 0 2518 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1704
transform 1 0 2444 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1705
transform 1 0 2419 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1706
transform 1 0 2407 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1707
transform 1 0 2338 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1708
transform 1 0 2313 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1709
transform 1 0 2441 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1710
transform 1 0 2575 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1711
transform 1 0 2459 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1712
transform 1 0 2581 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1713
transform 1 0 2465 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1714
transform 1 0 2233 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1715
transform 1 0 2524 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1716
transform 1 0 2456 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1717
transform 1 0 2413 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1718
transform 1 0 2395 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1719
transform 1 0 2350 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1720
transform 1 0 2492 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1721
transform 1 0 2431 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1722
transform 1 0 2440 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1723
transform 1 0 2386 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1724
transform 1 0 2274 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1725
transform 1 0 2320 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1726
transform 1 0 2335 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1727
transform 1 0 2335 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1728
transform 1 0 2414 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1729
transform 1 0 2705 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1730
transform 1 0 2420 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1731
transform 1 0 2482 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1732
transform 1 0 2359 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1733
transform 1 0 2272 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1734
transform 1 0 2352 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1735
transform 1 0 2513 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1736
transform 1 0 2389 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1737
transform 1 0 2383 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1738
transform 1 0 2383 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1739
transform 1 0 2371 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1740
transform 1 0 2356 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1741
transform 1 0 2307 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1742
transform 1 0 2232 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1743
transform 1 0 2250 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1744
transform 1 0 2325 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1745
transform 1 0 2398 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1746
transform 1 0 2549 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1747
transform 1 0 2535 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1748
transform 1 0 2679 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1749
transform 1 0 2689 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1750
transform 1 0 2618 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1751
transform 1 0 2692 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1752
transform 1 0 2707 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1753
transform 1 0 2552 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1754
transform 1 0 2417 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1755
transform 1 0 2430 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1756
transform 1 0 2428 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1757
transform 1 0 2455 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1758
transform 1 0 2397 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1759
transform 1 0 2341 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1760
transform 1 0 2341 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1761
transform 1 0 2432 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1762
transform 1 0 2494 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1763
transform 1 0 2386 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1764
transform 1 0 2249 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1765
transform 1 0 2671 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1766
transform 1 0 2525 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1767
transform 1 0 2403 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1768
transform 1 0 2351 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1769
transform 1 0 2343 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1770
transform 1 0 2386 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1771
transform 1 0 2188 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-1772
transform 1 0 2108 0 1 5755
box 0 0 3 6
use FEEDTHRU  F-1773
transform 1 0 2392 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1774
transform 1 0 2446 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1775
transform 1 0 2461 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1776
transform 1 0 2280 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1777
transform 1 0 2490 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1778
transform 1 0 2408 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1779
transform 1 0 2300 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1780
transform 1 0 2353 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1781
transform 1 0 2229 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1782
transform 1 0 2314 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1783
transform 1 0 2283 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1784
transform 1 0 2270 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1785
transform 1 0 2311 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1786
transform 1 0 2591 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1787
transform 1 0 2594 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1788
transform 1 0 2199 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1789
transform 1 0 2196 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1790
transform 1 0 2260 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1791
transform 1 0 2216 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1792
transform 1 0 2313 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1793
transform 1 0 2366 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1794
transform 1 0 2296 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1795
transform 1 0 2267 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1796
transform 1 0 2398 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1797
transform 1 0 2412 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1798
transform 1 0 2402 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1799
transform 1 0 2354 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1800
transform 1 0 2301 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1801
transform 1 0 2306 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1802
transform 1 0 2289 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1803
transform 1 0 2320 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1804
transform 1 0 2389 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1805
transform 1 0 2360 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1806
transform 1 0 2448 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1807
transform 1 0 2513 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1808
transform 1 0 2431 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1809
transform 1 0 2685 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1810
transform 1 0 2554 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1811
transform 1 0 2538 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1812
transform 1 0 2531 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1813
transform 1 0 2695 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1814
transform 1 0 2555 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1815
transform 1 0 2641 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1816
transform 1 0 2585 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1817
transform 1 0 2509 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1818
transform 1 0 2500 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1819
transform 1 0 2518 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1820
transform 1 0 2600 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1821
transform 1 0 2659 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1822
transform 1 0 2579 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1823
transform 1 0 2713 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1824
transform 1 0 2352 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1825
transform 1 0 2289 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1826
transform 1 0 2373 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1827
transform 1 0 2437 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1828
transform 1 0 2626 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1829
transform 1 0 2570 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1830
transform 1 0 2290 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1831
transform 1 0 2467 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1832
transform 1 0 2440 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1833
transform 1 0 2385 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1834
transform 1 0 2298 0 1 1138
box 0 0 3 6
use FEEDTHRU  F-1835
transform 1 0 2270 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1836
transform 1 0 2328 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1837
transform 1 0 2285 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-1838
transform 1 0 2344 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1839
transform 1 0 2353 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1840
transform 1 0 2347 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1841
transform 1 0 2341 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1842
transform 1 0 2306 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1843
transform 1 0 2348 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1844
transform 1 0 2476 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1845
transform 1 0 2344 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1846
transform 1 0 2300 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1847
transform 1 0 2338 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1848
transform 1 0 2424 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1849
transform 1 0 2489 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1850
transform 1 0 2401 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1851
transform 1 0 2378 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1852
transform 1 0 2368 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1853
transform 1 0 2377 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1854
transform 1 0 2377 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1855
transform 1 0 2234 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1856
transform 1 0 2368 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1857
transform 1 0 2370 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1858
transform 1 0 2375 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1859
transform 1 0 2316 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1860
transform 1 0 2322 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1861
transform 1 0 2304 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1862
transform 1 0 2246 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-1863
transform 1 0 2384 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1864
transform 1 0 2518 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1865
transform 1 0 2198 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1866
transform 1 0 2236 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1867
transform 1 0 2584 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1868
transform 1 0 2483 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1869
transform 1 0 2635 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1870
transform 1 0 2465 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1871
transform 1 0 2472 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1872
transform 1 0 2470 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1873
transform 1 0 2336 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1874
transform 1 0 2213 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1875
transform 1 0 2199 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1876
transform 1 0 2230 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1877
transform 1 0 2296 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1878
transform 1 0 2255 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1879
transform 1 0 2376 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-1880
transform 1 0 2425 0 1 1386
box 0 0 3 6
use FEEDTHRU  F-1881
transform 1 0 2449 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1882
transform 1 0 2449 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1883
transform 1 0 2401 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1884
transform 1 0 2395 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1885
transform 1 0 2486 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1886
transform 1 0 2542 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1887
transform 1 0 2441 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1888
transform 1 0 2593 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1889
transform 1 0 2509 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1890
transform 1 0 2503 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1891
transform 1 0 2588 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1892
transform 1 0 2647 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1893
transform 1 0 2549 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1894
transform 1 0 2701 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1895
transform 1 0 2543 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1896
transform 1 0 2541 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1897
transform 1 0 2548 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1898
transform 1 0 2446 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1899
transform 1 0 2351 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1900
transform 1 0 2497 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1901
transform 1 0 2339 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1902
transform 1 0 2334 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1903
transform 1 0 2335 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1904
transform 1 0 2204 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1905
transform 1 0 2236 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1906
transform 1 0 2300 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1907
transform 1 0 2244 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1908
transform 1 0 2394 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1909
transform 1 0 2402 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1910
transform 1 0 2530 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1911
transform 1 0 2618 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1912
transform 1 0 2256 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1913
transform 1 0 2573 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1914
transform 1 0 2725 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1915
transform 1 0 2671 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1916
transform 1 0 2567 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1917
transform 1 0 2719 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1918
transform 1 0 2561 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1919
transform 1 0 2559 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1920
transform 1 0 2566 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1921
transform 1 0 2324 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1922
transform 1 0 2412 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1923
transform 1 0 2477 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1924
transform 1 0 2389 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1925
transform 1 0 2536 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1926
transform 1 0 2396 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1927
transform 1 0 2525 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1928
transform 1 0 2306 0 1 5668
box 0 0 3 6
use FEEDTHRU  F-1929
transform 1 0 2364 0 1 5551
box 0 0 3 6
use FEEDTHRU  F-1930
transform 1 0 2623 0 1 2800
box 0 0 3 6
use FEEDTHRU  F-1931
transform 1 0 2234 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1932
transform 1 0 2325 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1933
transform 1 0 2384 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1934
transform 1 0 2312 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1935
transform 1 0 2347 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1936
transform 1 0 2284 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1937
transform 1 0 2373 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1938
transform 1 0 2258 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1939
transform 1 0 2425 0 1 1573
box 0 0 3 6
use FEEDTHRU  F-1940
transform 1 0 2407 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1941
transform 1 0 2504 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1942
transform 1 0 2560 0 1 2250
box 0 0 3 6
use FEEDTHRU  F-1943
transform 1 0 2453 0 1 2511
box 0 0 3 6
use FEEDTHRU  F-1944
transform 1 0 2414 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1945
transform 1 0 2332 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1946
transform 1 0 2306 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1947
transform 1 0 2446 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1948
transform 1 0 2442 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1949
transform 1 0 2435 0 1 3085
box 0 0 3 6
use FEEDTHRU  F-1950
transform 1 0 2288 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1951
transform 1 0 2376 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1952
transform 1 0 2444 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1953
transform 1 0 2406 0 1 3322
box 0 0 3 6
use FEEDTHRU  F-1954
transform 1 0 2404 0 1 3547
box 0 0 3 6
use FEEDTHRU  F-1955
transform 1 0 2261 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1956
transform 1 0 2365 0 1 1760
box 0 0 3 6
use FEEDTHRU  F-1957
transform 1 0 2462 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1958
transform 1 0 2426 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1959
transform 1 0 2685 0 1 4021
box 0 0 3 6
use FEEDTHRU  F-1960
transform 1 0 2699 0 1 4240
box 0 0 3 6
use FEEDTHRU  F-1961
transform 1 0 2710 0 1 4463
box 0 0 3 6
use FEEDTHRU  F-1962
transform 1 0 2378 0 1 4704
box 0 0 3 6
use FEEDTHRU  F-1963
transform 1 0 2413 0 1 4897
box 0 0 3 6
use FEEDTHRU  F-1964
transform 1 0 2350 0 1 5100
box 0 0 3 6
use FEEDTHRU  F-1965
transform 1 0 2313 0 1 5273
box 0 0 3 6
use FEEDTHRU  F-1966
transform 1 0 2450 0 1 2013
box 0 0 3 6
use FEEDTHRU  F-1967
transform 1 0 2288 0 1 5418
box 0 0 3 6
use FEEDTHRU  F-1968
transform 1 0 2282 0 1 3796
box 0 0 3 6
<< metal1 >>
rect 2134 1007 2138 1008
rect 2077 1017 2148 1018
rect 2087 1019 2121 1020
rect 2101 1021 2130 1022
rect 2108 1023 2112 1024
rect 2131 1023 2175 1024
rect 2091 1025 2133 1026
rect 2134 1025 2199 1026
rect 2135 1027 2208 1028
rect 2137 1029 2184 1030
rect 2138 1031 2160 1032
rect 2140 1033 2212 1034
rect 2143 1035 2181 1036
rect 2150 1037 2172 1038
rect 2155 1039 2202 1040
rect 2156 1041 2228 1042
rect 2162 1043 2215 1044
rect 2195 1045 2222 1046
rect 2224 1045 2244 1046
rect 2233 1047 2237 1048
rect 2246 1047 2275 1048
rect 2255 1049 2265 1050
rect 2258 1051 2262 1052
rect 2084 1060 2231 1061
rect 2084 1062 2144 1063
rect 2087 1064 2160 1065
rect 2077 1066 2159 1067
rect 2078 1068 2390 1069
rect 2098 1070 2312 1071
rect 2114 1072 2252 1073
rect 2124 1074 2157 1075
rect 2129 1076 2177 1077
rect 2138 1078 2156 1079
rect 2152 1080 2163 1081
rect 2120 1082 2162 1083
rect 2111 1084 2122 1085
rect 2165 1084 2219 1085
rect 2168 1086 2267 1087
rect 2174 1088 2219 1089
rect 2180 1090 2279 1091
rect 2095 1092 2180 1093
rect 2201 1092 2228 1093
rect 2207 1094 2282 1095
rect 2185 1096 2207 1097
rect 2221 1096 2291 1097
rect 2224 1098 2324 1099
rect 2233 1100 2318 1101
rect 2091 1102 2234 1103
rect 2236 1102 2354 1103
rect 2147 1104 2237 1105
rect 2239 1104 2351 1105
rect 2167 1106 2240 1107
rect 2243 1106 2342 1107
rect 2171 1108 2243 1109
rect 2132 1110 2171 1111
rect 2246 1110 2339 1111
rect 2183 1112 2246 1113
rect 2182 1114 2196 1115
rect 2080 1116 2195 1117
rect 2081 1118 2128 1119
rect 2255 1118 2381 1119
rect 2211 1120 2255 1121
rect 2198 1122 2213 1123
rect 2258 1122 2384 1123
rect 2268 1124 2363 1125
rect 2088 1126 2270 1127
rect 2271 1126 2387 1127
rect 2274 1128 2407 1129
rect 2299 1130 2431 1131
rect 2335 1132 2394 1133
rect 2371 1134 2441 1135
rect 2409 1136 2417 1137
rect 2068 1145 2249 1146
rect 2072 1147 2276 1148
rect 2078 1149 2094 1150
rect 2084 1151 2273 1152
rect 2087 1153 2303 1154
rect 2098 1155 2294 1156
rect 2099 1157 2231 1158
rect 2108 1159 2180 1160
rect 2117 1161 2146 1162
rect 2121 1163 2405 1164
rect 2124 1165 2279 1166
rect 2135 1167 2267 1168
rect 2137 1169 2285 1170
rect 2143 1171 2173 1172
rect 2152 1173 2200 1174
rect 2155 1175 2288 1176
rect 2081 1177 2155 1178
rect 2161 1177 2279 1178
rect 2127 1179 2161 1180
rect 2128 1181 2315 1182
rect 2167 1183 2246 1184
rect 2065 1185 2246 1186
rect 2062 1187 2067 1188
rect 2176 1187 2221 1188
rect 2178 1189 2390 1190
rect 2182 1191 2195 1192
rect 2206 1191 2264 1192
rect 2212 1193 2297 1194
rect 2170 1195 2212 1196
rect 2233 1195 2309 1196
rect 2236 1197 2258 1198
rect 2239 1199 2330 1200
rect 2242 1201 2333 1202
rect 2251 1203 2327 1204
rect 2269 1205 2357 1206
rect 2080 1207 2270 1208
rect 2281 1207 2360 1208
rect 2281 1209 2444 1210
rect 2290 1211 2375 1212
rect 2114 1213 2291 1214
rect 2114 1215 2182 1216
rect 2299 1215 2387 1216
rect 2311 1217 2399 1218
rect 2117 1219 2312 1220
rect 2317 1219 2447 1220
rect 2131 1221 2318 1222
rect 2335 1221 2444 1222
rect 2218 1223 2336 1224
rect 2158 1225 2218 1226
rect 2338 1225 2519 1226
rect 2341 1227 2429 1228
rect 2254 1229 2342 1230
rect 2350 1229 2459 1230
rect 2353 1231 2462 1232
rect 2142 1233 2354 1234
rect 2362 1233 2465 1234
rect 2371 1235 2487 1236
rect 2380 1237 2503 1238
rect 2383 1239 2490 1240
rect 2377 1241 2384 1242
rect 2396 1241 2441 1242
rect 2406 1243 2410 1244
rect 2410 1245 2471 1246
rect 2430 1247 2493 1248
rect 2323 1249 2432 1250
rect 2433 1249 2468 1250
rect 2483 1249 2564 1250
rect 2515 1251 2522 1252
rect 2059 1260 2282 1261
rect 2068 1262 2109 1263
rect 2073 1264 2346 1265
rect 2072 1266 2246 1267
rect 2080 1268 2205 1269
rect 2086 1270 2202 1271
rect 2093 1272 2113 1273
rect 2096 1274 2370 1275
rect 2118 1276 2303 1277
rect 2124 1278 2409 1279
rect 2125 1280 2312 1281
rect 2128 1282 2352 1283
rect 2142 1284 2327 1285
rect 2131 1286 2142 1287
rect 2160 1286 2232 1287
rect 2165 1288 2173 1289
rect 2181 1288 2208 1289
rect 2189 1290 2200 1291
rect 2211 1290 2241 1291
rect 2220 1292 2253 1293
rect 2226 1294 2330 1295
rect 2178 1296 2226 1297
rect 2154 1298 2178 1299
rect 2233 1298 2354 1299
rect 2217 1300 2235 1301
rect 2272 1300 2313 1301
rect 2138 1302 2274 1303
rect 2275 1302 2322 1303
rect 2248 1304 2277 1305
rect 2278 1304 2349 1305
rect 2284 1306 2393 1307
rect 2287 1308 2391 1309
rect 2290 1310 2328 1311
rect 2079 1312 2292 1313
rect 2293 1312 2373 1313
rect 2296 1314 2364 1315
rect 2257 1316 2298 1317
rect 2096 1318 2259 1319
rect 2314 1318 2340 1319
rect 2263 1320 2316 1321
rect 2093 1322 2265 1323
rect 2317 1322 2355 1323
rect 2335 1324 2382 1325
rect 2236 1326 2337 1327
rect 2341 1326 2394 1327
rect 2356 1328 2397 1329
rect 2308 1330 2358 1331
rect 2269 1332 2310 1333
rect 2100 1334 2271 1335
rect 2359 1334 2418 1335
rect 2114 1336 2361 1337
rect 2374 1336 2439 1337
rect 2332 1338 2376 1339
rect 2121 1340 2334 1341
rect 2377 1340 2427 1341
rect 2410 1342 2472 1343
rect 2435 1344 2590 1345
rect 2440 1346 2535 1347
rect 2386 1348 2442 1349
rect 2090 1350 2388 1351
rect 2443 1350 2496 1351
rect 2446 1352 2508 1353
rect 2447 1354 2556 1355
rect 2458 1356 2520 1357
rect 2398 1358 2460 1359
rect 2145 1360 2400 1361
rect 2461 1360 2523 1361
rect 2464 1362 2526 1363
rect 2404 1364 2466 1365
rect 2229 1366 2406 1367
rect 2467 1366 2529 1367
rect 2483 1368 2544 1369
rect 2486 1370 2547 1371
rect 2489 1372 2577 1373
rect 2428 1374 2490 1375
rect 2492 1374 2565 1375
rect 2431 1376 2493 1377
rect 2365 1378 2433 1379
rect 2502 1378 2550 1379
rect 2515 1380 2608 1381
rect 2531 1382 2587 1383
rect 2567 1384 2622 1385
rect 2645 1384 2649 1385
rect 2065 1393 2325 1394
rect 2072 1395 2343 1396
rect 2082 1397 2319 1398
rect 2086 1399 2202 1400
rect 2093 1401 2328 1402
rect 2096 1403 2253 1404
rect 2096 1405 2241 1406
rect 2105 1407 2113 1408
rect 2108 1409 2148 1410
rect 2111 1411 2202 1412
rect 2115 1413 2253 1414
rect 2115 1415 2403 1416
rect 2118 1417 2505 1418
rect 2118 1419 2385 1420
rect 2122 1421 2367 1422
rect 2132 1423 2337 1424
rect 2134 1425 2142 1426
rect 2140 1427 2190 1428
rect 2143 1429 2391 1430
rect 2159 1431 2166 1432
rect 2177 1431 2190 1432
rect 2177 1433 2475 1434
rect 2195 1435 2208 1436
rect 2204 1437 2223 1438
rect 2219 1439 2400 1440
rect 2089 1441 2220 1442
rect 2225 1441 2244 1442
rect 2225 1443 2409 1444
rect 2228 1445 2394 1446
rect 2231 1447 2247 1448
rect 2234 1449 2238 1450
rect 2258 1449 2283 1450
rect 2068 1451 2259 1452
rect 2068 1453 2292 1454
rect 2264 1455 2289 1456
rect 2264 1457 2271 1458
rect 2276 1457 2328 1458
rect 2279 1459 2394 1460
rect 2297 1461 2331 1462
rect 2321 1463 2337 1464
rect 2333 1465 2391 1466
rect 2339 1467 2409 1468
rect 2354 1469 2412 1470
rect 2345 1471 2355 1472
rect 2369 1471 2379 1472
rect 2375 1473 2445 1474
rect 2405 1475 2457 1476
rect 2273 1477 2406 1478
rect 2414 1477 2499 1478
rect 2363 1479 2415 1480
rect 2417 1479 2487 1480
rect 2426 1481 2451 1482
rect 2156 1483 2427 1484
rect 2435 1483 2586 1484
rect 2396 1485 2436 1486
rect 2351 1487 2397 1488
rect 2312 1489 2352 1490
rect 2312 1491 2433 1492
rect 2381 1493 2433 1494
rect 2372 1495 2382 1496
rect 2357 1497 2373 1498
rect 2348 1499 2358 1500
rect 2309 1501 2349 1502
rect 2438 1501 2668 1502
rect 2125 1503 2439 1504
rect 2441 1503 2469 1504
rect 2387 1505 2442 1506
rect 2360 1507 2388 1508
rect 2315 1509 2361 1510
rect 2447 1509 2463 1510
rect 2453 1511 2583 1512
rect 2459 1513 2517 1514
rect 2459 1515 2553 1516
rect 2471 1517 2595 1518
rect 2501 1519 2574 1520
rect 2507 1521 2601 1522
rect 2510 1523 2729 1524
rect 2519 1525 2637 1526
rect 2522 1527 2640 1528
rect 2522 1529 2726 1530
rect 2525 1531 2607 1532
rect 2528 1533 2610 1534
rect 2465 1535 2529 1536
rect 2531 1535 2655 1536
rect 2534 1537 2658 1538
rect 2537 1539 2661 1540
rect 2540 1541 2592 1542
rect 2543 1543 2613 1544
rect 2276 1545 2544 1546
rect 2546 1545 2628 1546
rect 2546 1547 2664 1548
rect 2549 1549 2634 1550
rect 2564 1551 2625 1552
rect 2495 1553 2565 1554
rect 2306 1555 2496 1556
rect 2306 1557 2691 1558
rect 2567 1559 2652 1560
rect 2576 1561 2675 1562
rect 2489 1563 2577 1564
rect 2579 1563 2681 1564
rect 2492 1565 2580 1566
rect 2261 1567 2493 1568
rect 2630 1567 2736 1568
rect 2648 1569 2746 1570
rect 2621 1571 2649 1572
rect 2057 1580 2123 1581
rect 2072 1582 2095 1583
rect 2075 1584 2097 1585
rect 2075 1586 2307 1587
rect 2089 1588 2223 1589
rect 2101 1590 2220 1591
rect 2105 1592 2132 1593
rect 2111 1594 2196 1595
rect 2116 1596 2328 1597
rect 2119 1598 2361 1599
rect 2128 1600 2160 1601
rect 2134 1602 2154 1603
rect 2134 1604 2304 1605
rect 2140 1606 2184 1607
rect 2143 1608 2466 1609
rect 2171 1610 2565 1611
rect 2189 1612 2220 1613
rect 2201 1614 2235 1615
rect 2225 1616 2241 1617
rect 2231 1618 2684 1619
rect 2237 1620 2268 1621
rect 2258 1622 2415 1623
rect 2243 1624 2259 1625
rect 2261 1624 2481 1625
rect 2252 1626 2262 1627
rect 2246 1628 2253 1629
rect 2264 1628 2274 1629
rect 2276 1628 2640 1629
rect 2282 1630 2292 1631
rect 2285 1632 2358 1633
rect 2288 1634 2298 1635
rect 2315 1634 2705 1635
rect 2318 1636 2322 1637
rect 2324 1636 2328 1637
rect 2351 1636 2370 1637
rect 2098 1638 2352 1639
rect 2363 1638 2505 1639
rect 2396 1640 2415 1641
rect 2396 1642 2403 1643
rect 2390 1644 2403 1645
rect 2384 1646 2391 1647
rect 2372 1648 2385 1649
rect 2366 1650 2373 1651
rect 2082 1652 2367 1653
rect 2068 1654 2082 1655
rect 2068 1656 2166 1657
rect 2399 1656 2406 1657
rect 2393 1658 2406 1659
rect 2387 1660 2394 1661
rect 2408 1660 2421 1661
rect 2408 1662 2427 1663
rect 2411 1664 2424 1665
rect 2432 1664 2553 1665
rect 2432 1666 2442 1667
rect 2435 1668 2556 1669
rect 2459 1670 2490 1671
rect 2462 1672 2727 1673
rect 2438 1674 2463 1675
rect 2438 1676 2671 1677
rect 2468 1678 2668 1679
rect 2456 1680 2469 1681
rect 2456 1682 2670 1683
rect 2474 1684 2589 1685
rect 2150 1686 2475 1687
rect 2486 1686 2532 1687
rect 2444 1688 2487 1689
rect 2162 1690 2445 1691
rect 2492 1690 2559 1691
rect 2495 1692 2562 1693
rect 2504 1694 2511 1695
rect 2501 1696 2511 1697
rect 2516 1696 2526 1697
rect 2498 1698 2517 1699
rect 2519 1698 2785 1699
rect 2522 1700 2538 1701
rect 2543 1700 2571 1701
rect 2543 1702 2610 1703
rect 2546 1704 2592 1705
rect 2528 1706 2547 1707
rect 2564 1706 2792 1707
rect 2582 1708 2667 1709
rect 2582 1710 2675 1711
rect 2585 1712 2664 1713
rect 2594 1714 2685 1715
rect 2540 1716 2595 1717
rect 2600 1716 2712 1717
rect 2579 1718 2601 1719
rect 2606 1718 2698 1719
rect 2624 1720 2795 1721
rect 2627 1722 2676 1723
rect 2576 1724 2628 1725
rect 2360 1726 2577 1727
rect 2630 1726 2788 1727
rect 2633 1728 2679 1729
rect 2636 1730 2709 1731
rect 2636 1732 2767 1733
rect 2639 1734 2764 1735
rect 2642 1736 2757 1737
rect 2648 1738 2697 1739
rect 2651 1740 2700 1741
rect 2654 1742 2721 1743
rect 2612 1744 2655 1745
rect 2657 1744 2724 1745
rect 2312 1746 2658 1747
rect 2159 1748 2313 1749
rect 2660 1748 2715 1749
rect 2279 1750 2661 1751
rect 2137 1752 2280 1753
rect 2680 1752 2740 1753
rect 2681 1754 2719 1755
rect 2513 1756 2718 1757
rect 2745 1756 2819 1757
rect 2808 1758 2813 1759
rect 2047 1767 2123 1768
rect 2054 1769 2076 1770
rect 2059 1771 2076 1772
rect 2061 1773 2082 1774
rect 2071 1775 2455 1776
rect 2064 1777 2073 1778
rect 2078 1777 2166 1778
rect 2087 1779 2349 1780
rect 2089 1781 2235 1782
rect 2082 1783 2236 1784
rect 2092 1785 2377 1786
rect 2113 1787 2355 1788
rect 2116 1789 2385 1790
rect 2119 1791 2391 1792
rect 2119 1793 2132 1794
rect 2125 1795 2424 1796
rect 2128 1797 2461 1798
rect 2129 1799 2154 1800
rect 2134 1801 2257 1802
rect 2137 1803 2274 1804
rect 2144 1805 2445 1806
rect 2125 1807 2145 1808
rect 2148 1807 2500 1808
rect 2171 1809 2379 1810
rect 2174 1811 2280 1812
rect 2181 1813 2490 1814
rect 2202 1815 2232 1816
rect 2205 1817 2220 1818
rect 2207 1819 2487 1820
rect 2210 1821 2674 1822
rect 2223 1823 2253 1824
rect 2229 1825 2394 1826
rect 2240 1827 2473 1828
rect 2241 1829 2259 1830
rect 2244 1831 2310 1832
rect 2250 1833 2268 1834
rect 2268 1835 2292 1836
rect 2274 1837 2298 1838
rect 2280 1839 2304 1840
rect 2289 1841 2628 1842
rect 2292 1843 2316 1844
rect 2310 1845 2322 1846
rect 2312 1847 2716 1848
rect 2316 1849 2331 1850
rect 2322 1851 2373 1852
rect 2327 1853 2392 1854
rect 2328 1855 2403 1856
rect 2151 1857 2404 1858
rect 2331 1859 2406 1860
rect 2334 1861 2571 1862
rect 2346 1863 2439 1864
rect 2351 1865 2437 1866
rect 2352 1867 2553 1868
rect 2355 1869 2556 1870
rect 2360 1871 2589 1872
rect 2363 1873 2595 1874
rect 2364 1875 2562 1876
rect 2379 1877 2658 1878
rect 2385 1879 2463 1880
rect 2366 1881 2464 1882
rect 2396 1883 2488 1884
rect 2101 1885 2398 1886
rect 2399 1885 2491 1886
rect 2381 1887 2401 1888
rect 2420 1887 2446 1888
rect 2068 1889 2422 1890
rect 2069 1891 2320 1892
rect 2427 1891 2809 1892
rect 2432 1893 2494 1894
rect 2342 1895 2434 1896
rect 2439 1895 2469 1896
rect 2098 1897 2470 1898
rect 2465 1899 2509 1900
rect 2369 1901 2467 1902
rect 2370 1903 2532 1904
rect 2474 1905 2734 1906
rect 2475 1907 2565 1908
rect 2484 1909 2559 1910
rect 2504 1911 2590 1912
rect 2408 1913 2506 1914
rect 2159 1915 2410 1916
rect 2160 1917 2184 1918
rect 2510 1917 2587 1918
rect 2511 1919 2730 1920
rect 2516 1921 2542 1922
rect 2141 1923 2518 1924
rect 2141 1925 2299 1926
rect 2523 1925 2547 1926
rect 2525 1927 2554 1928
rect 2529 1929 2538 1930
rect 2547 1929 2643 1930
rect 2550 1931 2661 1932
rect 2559 1933 2583 1934
rect 2571 1935 2750 1936
rect 2580 1937 2776 1938
rect 2613 1939 2664 1940
rect 2616 1941 2667 1942
rect 2619 1943 2851 1944
rect 2624 1945 2635 1946
rect 2628 1947 2724 1948
rect 2636 1949 2662 1950
rect 2600 1951 2638 1952
rect 2519 1953 2602 1954
rect 2639 1953 2650 1954
rect 2640 1955 2840 1956
rect 2667 1957 2764 1958
rect 2576 1959 2764 1960
rect 2543 1961 2578 1962
rect 2513 1963 2545 1964
rect 2675 1963 2704 1964
rect 2678 1965 2725 1966
rect 2654 1967 2680 1968
rect 2681 1967 2753 1968
rect 2682 1969 2844 1970
rect 2696 1971 2761 1972
rect 2697 1973 2709 1974
rect 2699 1975 2728 1976
rect 2700 1977 2712 1978
rect 2706 1979 2792 1980
rect 2720 1981 2785 1982
rect 2736 1983 2743 1984
rect 2739 1985 2770 1986
rect 2739 1987 2802 1988
rect 2742 1989 2767 1990
rect 2450 1991 2767 1992
rect 2084 1993 2452 1994
rect 2085 1995 2262 1996
rect 2262 1997 2286 1998
rect 2286 1999 2457 2000
rect 2414 2001 2458 2002
rect 2336 2003 2416 2004
rect 2757 2003 2830 2004
rect 2772 2005 2779 2006
rect 2781 2005 2791 2006
rect 2797 2005 2809 2006
rect 2812 2005 2822 2006
rect 2811 2007 2826 2008
rect 2818 2009 2857 2010
rect 2721 2011 2819 2012
rect 2822 2011 2847 2012
rect 2011 2020 2448 2021
rect 2066 2022 2464 2023
rect 2069 2024 2452 2025
rect 2072 2026 2382 2027
rect 2078 2028 2172 2029
rect 2092 2030 2123 2031
rect 2104 2032 2161 2033
rect 2110 2034 2437 2035
rect 2113 2036 2410 2037
rect 2119 2038 2136 2039
rect 2129 2040 2491 2041
rect 2141 2042 2502 2043
rect 2141 2044 2416 2045
rect 2144 2046 2440 2047
rect 2148 2048 2386 2049
rect 2148 2050 2230 2051
rect 2152 2052 2311 2053
rect 2155 2054 2494 2055
rect 2159 2056 2490 2057
rect 2178 2058 2208 2059
rect 2075 2060 2178 2061
rect 2181 2060 2493 2061
rect 2190 2062 2716 2063
rect 2202 2064 2451 2065
rect 2205 2066 2232 2067
rect 2243 2068 2473 2069
rect 2256 2070 2325 2071
rect 2219 2072 2256 2073
rect 2262 2072 2307 2073
rect 2264 2074 2604 2075
rect 2268 2076 2313 2077
rect 2082 2078 2268 2079
rect 2276 2078 2467 2079
rect 2280 2080 2850 2081
rect 2250 2082 2280 2083
rect 2289 2082 2698 2083
rect 2292 2084 2343 2085
rect 2241 2086 2292 2087
rect 2298 2086 2349 2087
rect 2316 2088 2361 2089
rect 2322 2090 2367 2091
rect 2328 2092 2373 2093
rect 2346 2094 2385 2095
rect 2352 2096 2409 2097
rect 2364 2098 2415 2099
rect 2319 2100 2364 2101
rect 2274 2102 2319 2103
rect 2235 2104 2274 2105
rect 2370 2104 2430 2105
rect 2397 2106 2466 2107
rect 2379 2108 2397 2109
rect 2059 2110 2379 2111
rect 2427 2110 2472 2111
rect 2376 2112 2427 2113
rect 2331 2114 2376 2115
rect 2125 2116 2331 2117
rect 2125 2118 2196 2119
rect 2433 2118 2496 2119
rect 2445 2120 2520 2121
rect 2444 2122 2485 2123
rect 2421 2124 2484 2125
rect 2193 2126 2421 2127
rect 2457 2126 2526 2127
rect 2469 2128 2478 2129
rect 2475 2130 2514 2131
rect 2481 2132 2532 2133
rect 2499 2134 2538 2135
rect 2076 2136 2499 2137
rect 2505 2136 2562 2137
rect 2400 2138 2505 2139
rect 2508 2138 2565 2139
rect 2116 2140 2508 2141
rect 2511 2140 2790 2141
rect 2355 2142 2511 2143
rect 2334 2144 2355 2145
rect 2517 2144 2853 2145
rect 2523 2146 2574 2147
rect 2541 2148 2598 2149
rect 2544 2150 2802 2151
rect 2487 2152 2544 2153
rect 2069 2154 2487 2155
rect 2547 2154 2568 2155
rect 2286 2156 2547 2157
rect 2555 2156 2560 2157
rect 2586 2156 2643 2157
rect 2261 2158 2586 2159
rect 2609 2158 2776 2159
rect 2619 2160 2833 2161
rect 2621 2162 2773 2163
rect 2640 2164 2709 2165
rect 2577 2166 2640 2167
rect 2649 2166 2751 2167
rect 2589 2168 2649 2169
rect 2247 2170 2589 2171
rect 2667 2170 2763 2171
rect 2637 2172 2667 2173
rect 2673 2172 2866 2173
rect 2672 2174 2943 2175
rect 2676 2176 2707 2177
rect 2682 2178 2772 2179
rect 2685 2180 2860 2181
rect 2628 2182 2685 2183
rect 2571 2184 2628 2185
rect 2550 2186 2571 2187
rect 2690 2186 2908 2187
rect 2693 2188 2890 2189
rect 2696 2190 2901 2191
rect 2703 2192 2805 2193
rect 2711 2194 2755 2195
rect 2718 2196 2799 2197
rect 2721 2198 2820 2199
rect 2724 2200 2823 2201
rect 2729 2202 2936 2203
rect 2739 2204 2838 2205
rect 2616 2206 2739 2207
rect 2553 2208 2616 2209
rect 2742 2208 2841 2209
rect 2747 2210 2955 2211
rect 2757 2212 2826 2213
rect 2661 2214 2757 2215
rect 2601 2216 2661 2217
rect 2727 2216 2826 2217
rect 2760 2218 2878 2219
rect 2766 2220 2897 2221
rect 2769 2222 2863 2223
rect 2679 2224 2769 2225
rect 2781 2224 2881 2225
rect 2613 2226 2781 2227
rect 2784 2226 2884 2227
rect 2735 2228 2784 2229
rect 2787 2228 2795 2229
rect 2634 2230 2796 2231
rect 2580 2232 2634 2233
rect 2529 2234 2580 2235
rect 2460 2236 2529 2237
rect 2391 2238 2460 2239
rect 2390 2240 2455 2241
rect 2403 2242 2454 2243
rect 2145 2244 2403 2245
rect 2700 2244 2787 2245
rect 2792 2244 2869 2245
rect 2856 2246 2949 2247
rect 2702 2248 2857 2249
rect 2874 2248 2922 2249
rect 2045 2257 2050 2258
rect 2062 2257 2484 2258
rect 2066 2259 2391 2260
rect 2070 2261 2487 2262
rect 2080 2263 2111 2264
rect 2088 2265 2230 2266
rect 2089 2267 2499 2268
rect 2097 2269 2401 2270
rect 2098 2271 2323 2272
rect 2107 2273 2172 2274
rect 2107 2275 2232 2276
rect 2117 2277 2419 2278
rect 2125 2279 2364 2280
rect 2126 2281 2367 2282
rect 2129 2283 2526 2284
rect 2138 2285 2155 2286
rect 2141 2287 2466 2288
rect 2143 2289 2496 2290
rect 2157 2291 2470 2292
rect 2159 2293 2289 2294
rect 2135 2295 2161 2296
rect 2162 2295 2478 2296
rect 2152 2297 2164 2298
rect 2177 2297 2194 2298
rect 2187 2299 2565 2300
rect 2195 2301 2212 2302
rect 2199 2303 2208 2304
rect 2217 2303 2529 2304
rect 2219 2305 2511 2306
rect 2222 2307 2608 2308
rect 2243 2309 2290 2310
rect 2250 2311 2497 2312
rect 2255 2313 2347 2314
rect 2259 2315 2280 2316
rect 2267 2317 2272 2318
rect 2276 2317 2281 2318
rect 2273 2319 2278 2320
rect 2291 2319 2296 2320
rect 2304 2319 2313 2320
rect 2076 2321 2314 2322
rect 2306 2323 2311 2324
rect 2316 2323 2319 2324
rect 2324 2323 2329 2324
rect 2330 2323 2335 2324
rect 2340 2323 2343 2324
rect 2348 2323 2365 2324
rect 2352 2325 2448 2326
rect 2166 2327 2449 2328
rect 2358 2329 2379 2330
rect 2360 2331 2371 2332
rect 2361 2333 2382 2334
rect 2372 2335 2395 2336
rect 2122 2337 2374 2338
rect 2382 2337 2460 2338
rect 2148 2339 2461 2340
rect 2147 2341 2266 2342
rect 2391 2341 2427 2342
rect 2247 2343 2428 2344
rect 2402 2345 2479 2346
rect 2406 2347 2502 2348
rect 2412 2349 2746 2350
rect 2424 2351 2520 2352
rect 2429 2353 2593 2354
rect 2436 2355 2454 2356
rect 2442 2357 2544 2358
rect 2136 2359 2545 2360
rect 2454 2361 2562 2362
rect 2466 2363 2872 2364
rect 2475 2365 2493 2366
rect 2484 2367 2586 2368
rect 2502 2369 2508 2370
rect 2420 2371 2509 2372
rect 2421 2373 2505 2374
rect 2520 2373 2574 2374
rect 2526 2375 2890 2376
rect 2550 2377 2649 2378
rect 2574 2379 2946 2380
rect 2609 2381 2656 2382
rect 2619 2383 2694 2384
rect 2621 2385 2650 2386
rect 2627 2387 2904 2388
rect 2628 2389 2709 2390
rect 2537 2391 2710 2392
rect 2414 2393 2539 2394
rect 2415 2395 2623 2396
rect 2631 2395 2634 2396
rect 2637 2395 2703 2396
rect 2555 2397 2704 2398
rect 2556 2399 2643 2400
rect 2639 2401 2845 2402
rect 2679 2403 2748 2404
rect 2588 2405 2749 2406
rect 2684 2407 2901 2408
rect 2471 2409 2686 2410
rect 2472 2411 2490 2412
rect 2490 2413 2532 2414
rect 2532 2415 2580 2416
rect 2580 2417 2661 2418
rect 2444 2419 2662 2420
rect 2445 2421 2547 2422
rect 2696 2421 2936 2422
rect 2697 2423 2959 2424
rect 2241 2425 2960 2426
rect 2700 2427 2967 2428
rect 2715 2429 2915 2430
rect 2729 2431 2734 2432
rect 2735 2431 2830 2432
rect 2738 2433 2833 2434
rect 2750 2435 2932 2436
rect 2396 2437 2752 2438
rect 2375 2439 2398 2440
rect 2100 2441 2377 2442
rect 2756 2441 2939 2442
rect 2757 2443 2763 2444
rect 2666 2445 2764 2446
rect 2667 2447 2946 2448
rect 2760 2449 2796 2450
rect 2771 2451 2776 2452
rect 2768 2453 2773 2454
rect 2784 2453 2814 2454
rect 2786 2455 2848 2456
rect 2597 2457 2788 2458
rect 2513 2459 2599 2460
rect 2789 2459 2851 2460
rect 2570 2461 2791 2462
rect 2796 2461 2805 2462
rect 2567 2463 2806 2464
rect 2568 2465 2673 2466
rect 2673 2467 2712 2468
rect 2798 2467 2871 2468
rect 2801 2469 2817 2470
rect 2811 2471 2820 2472
rect 2814 2473 2823 2474
rect 2817 2475 2826 2476
rect 2823 2477 2878 2478
rect 2837 2479 2892 2480
rect 2840 2481 2869 2482
rect 2792 2483 2868 2484
rect 2354 2485 2794 2486
rect 2355 2487 2451 2488
rect 2841 2487 2894 2488
rect 2852 2489 2857 2490
rect 2603 2491 2857 2492
rect 2408 2493 2605 2494
rect 2865 2493 2889 2494
rect 2874 2495 2919 2496
rect 2873 2497 2953 2498
rect 2880 2499 2898 2500
rect 2879 2501 2939 2502
rect 2883 2503 2887 2504
rect 2862 2505 2886 2506
rect 2615 2507 2864 2508
rect 2616 2509 2691 2510
rect 2915 2509 2922 2510
rect 2948 2509 2970 2510
rect 2035 2518 2362 2519
rect 2038 2520 2043 2521
rect 2049 2520 2057 2521
rect 2063 2520 2359 2521
rect 2080 2522 2105 2523
rect 2084 2524 2090 2525
rect 2093 2524 2337 2525
rect 2095 2526 2539 2527
rect 2098 2528 2794 2529
rect 2100 2530 2419 2531
rect 2110 2532 2481 2533
rect 2077 2534 2111 2535
rect 2114 2534 2188 2535
rect 2129 2536 2509 2537
rect 2133 2538 2425 2539
rect 2139 2540 2238 2541
rect 2142 2542 2161 2543
rect 2145 2544 2395 2545
rect 2147 2546 2260 2547
rect 2148 2548 2403 2549
rect 2176 2550 2200 2551
rect 2188 2552 2212 2553
rect 2206 2554 2230 2555
rect 2224 2556 2479 2557
rect 2227 2558 2266 2559
rect 2231 2560 2553 2561
rect 2243 2562 2290 2563
rect 2247 2564 2503 2565
rect 2255 2566 2562 2567
rect 2261 2568 2272 2569
rect 2267 2570 2278 2571
rect 2291 2570 2329 2571
rect 2297 2572 2323 2573
rect 2304 2574 2319 2575
rect 2303 2576 2386 2577
rect 2310 2578 2331 2579
rect 2316 2580 2325 2581
rect 2295 2582 2316 2583
rect 2340 2582 2361 2583
rect 2342 2584 2752 2585
rect 2352 2586 2499 2587
rect 2355 2588 2502 2589
rect 2334 2590 2355 2591
rect 2313 2592 2334 2593
rect 2366 2592 2605 2593
rect 2373 2594 2487 2595
rect 2364 2596 2373 2597
rect 2376 2596 2385 2597
rect 2375 2598 2428 2599
rect 2066 2600 2427 2601
rect 2391 2602 2478 2603
rect 2390 2604 2746 2605
rect 2406 2606 2529 2607
rect 2408 2608 2861 2609
rect 2412 2610 2430 2611
rect 2397 2612 2412 2613
rect 2370 2614 2397 2615
rect 2415 2614 2662 2615
rect 2400 2616 2415 2617
rect 2436 2616 2586 2617
rect 2435 2618 2623 2619
rect 2442 2620 2595 2621
rect 2166 2622 2442 2623
rect 2167 2624 2455 2625
rect 2448 2626 2454 2627
rect 2163 2628 2448 2629
rect 2164 2630 2625 2631
rect 2460 2632 2577 2633
rect 2466 2634 2583 2635
rect 2097 2636 2466 2637
rect 2472 2636 2535 2637
rect 2475 2638 2538 2639
rect 2474 2640 2833 2641
rect 2490 2642 2547 2643
rect 2489 2644 2686 2645
rect 2496 2646 2936 2647
rect 2382 2648 2496 2649
rect 2510 2648 2710 2649
rect 2516 2650 2836 2651
rect 2520 2652 2736 2653
rect 2522 2654 2599 2655
rect 2445 2656 2598 2657
rect 2544 2658 2559 2659
rect 2568 2658 2721 2659
rect 2567 2660 2785 2661
rect 2570 2662 2704 2663
rect 2550 2664 2703 2665
rect 2574 2666 2727 2667
rect 2592 2668 2878 2669
rect 2607 2670 2806 2671
rect 2532 2672 2607 2673
rect 2421 2674 2532 2675
rect 2420 2676 2716 2677
rect 2580 2678 2715 2679
rect 2612 2680 2656 2681
rect 2616 2682 2712 2683
rect 2619 2684 2691 2685
rect 2618 2686 2857 2687
rect 2628 2688 2751 2689
rect 2346 2690 2628 2691
rect 2639 2690 2749 2691
rect 2654 2692 2892 2693
rect 2657 2694 2761 2695
rect 2621 2696 2760 2697
rect 2667 2698 2907 2699
rect 2673 2700 2946 2701
rect 2526 2702 2673 2703
rect 2525 2704 2830 2705
rect 2679 2706 2939 2707
rect 2469 2708 2679 2709
rect 2280 2710 2469 2711
rect 2129 2712 2280 2713
rect 2684 2712 2734 2713
rect 2697 2714 2983 2715
rect 2556 2716 2697 2717
rect 2700 2716 2980 2717
rect 2708 2718 2892 2719
rect 2732 2720 2848 2721
rect 2738 2722 2973 2723
rect 2744 2724 2913 2725
rect 2757 2726 2864 2727
rect 2763 2728 2895 2729
rect 2631 2730 2895 2731
rect 2630 2732 2650 2733
rect 2648 2734 2901 2735
rect 2637 2736 2902 2737
rect 2484 2738 2637 2739
rect 2126 2740 2484 2741
rect 2125 2742 2194 2743
rect 2194 2744 2218 2745
rect 2218 2746 2242 2747
rect 2772 2746 2778 2747
rect 2783 2746 2797 2747
rect 2787 2748 2854 2749
rect 2786 2750 2967 2751
rect 2792 2752 2845 2753
rect 2122 2754 2845 2755
rect 2795 2756 2812 2757
rect 2154 2758 2811 2759
rect 2798 2760 2815 2761
rect 2790 2762 2815 2763
rect 2789 2764 2842 2765
rect 2801 2766 2824 2767
rect 2808 2768 2839 2769
rect 2807 2770 2851 2771
rect 2817 2772 2964 2773
rect 2820 2774 2886 2775
rect 2823 2776 2889 2777
rect 2826 2778 2909 2779
rect 2829 2780 2874 2781
rect 2841 2782 2898 2783
rect 2859 2784 2943 2785
rect 2862 2786 2929 2787
rect 2871 2788 2916 2789
rect 2775 2790 2916 2791
rect 2874 2792 2919 2793
rect 2879 2794 2950 2795
rect 2918 2796 2970 2797
rect 2935 2798 2943 2799
rect 2059 2807 2155 2808
rect 2065 2809 2481 2810
rect 2068 2811 2085 2812
rect 2069 2813 2111 2814
rect 2075 2815 2262 2816
rect 2076 2817 2496 2818
rect 2083 2819 2466 2820
rect 2087 2821 2427 2822
rect 2093 2823 2628 2824
rect 2094 2825 2189 2826
rect 2097 2827 2478 2828
rect 2104 2829 2526 2830
rect 2119 2831 2373 2832
rect 2122 2833 2334 2834
rect 2125 2835 2397 2836
rect 2080 2837 2126 2838
rect 2129 2837 2469 2838
rect 2112 2839 2470 2840
rect 2131 2841 2448 2842
rect 2136 2843 2385 2844
rect 2135 2845 2215 2846
rect 2142 2847 2158 2848
rect 2142 2849 2535 2850
rect 2145 2851 2335 2852
rect 2145 2853 2583 2854
rect 2160 2855 2487 2856
rect 2163 2857 2195 2858
rect 2167 2859 2595 2860
rect 2176 2861 2191 2862
rect 2178 2863 2219 2864
rect 2196 2865 2367 2866
rect 2199 2867 2625 2868
rect 2202 2869 2244 2870
rect 2206 2871 2290 2872
rect 2208 2873 2238 2874
rect 2220 2875 2407 2876
rect 2224 2877 2707 2878
rect 2223 2879 2640 2880
rect 2227 2881 2329 2882
rect 2231 2883 2436 2884
rect 2152 2885 2437 2886
rect 2232 2887 2268 2888
rect 2244 2889 2280 2890
rect 2262 2891 2292 2892
rect 2268 2893 2316 2894
rect 2271 2895 2319 2896
rect 2277 2897 2325 2898
rect 2283 2899 2331 2900
rect 2286 2901 2337 2902
rect 2297 2903 2395 2904
rect 2303 2905 2332 2906
rect 2304 2907 2355 2908
rect 2310 2909 2361 2910
rect 2313 2911 2376 2912
rect 2072 2913 2377 2914
rect 2322 2915 2343 2916
rect 2340 2917 2499 2918
rect 2343 2919 2502 2920
rect 2346 2921 2403 2922
rect 2352 2923 2415 2924
rect 2355 2925 2598 2926
rect 2358 2927 2409 2928
rect 2364 2929 2421 2930
rect 2370 2931 2430 2932
rect 2379 2933 2454 2934
rect 2382 2935 2538 2936
rect 2385 2937 2391 2938
rect 2391 2939 2484 2940
rect 2397 2941 2529 2942
rect 2400 2943 2532 2944
rect 2403 2945 2763 2946
rect 2411 2947 2440 2948
rect 2424 2949 2490 2950
rect 2430 2951 2517 2952
rect 2441 2953 2485 2954
rect 2442 2955 2577 2956
rect 2445 2957 2586 2958
rect 2448 2959 2523 2960
rect 2454 2961 2553 2962
rect 2460 2963 2547 2964
rect 2466 2965 2637 2966
rect 2472 2967 2559 2968
rect 2474 2969 2482 2970
rect 2475 2971 2562 2972
rect 2478 2973 2511 2974
rect 2490 2975 2736 2976
rect 2496 2977 2811 2978
rect 2508 2979 2631 2980
rect 2514 2981 2731 2982
rect 2526 2983 2878 2984
rect 2532 2985 2697 2986
rect 2544 2987 2703 2988
rect 2550 2989 2895 2990
rect 2553 2991 2709 2992
rect 2556 2993 2613 2994
rect 2562 2995 2721 2996
rect 2567 2997 2689 2998
rect 2241 2999 2569 3000
rect 2570 2999 2760 3000
rect 2574 3001 2839 3002
rect 2580 3003 2649 3004
rect 2592 3005 2854 3006
rect 2595 3007 2847 3008
rect 2598 3009 2902 3010
rect 2604 3011 2745 3012
rect 2606 3013 2719 3014
rect 2610 3015 2751 3016
rect 2613 3017 2824 3018
rect 2618 3019 2818 3020
rect 2631 3021 2655 3022
rect 2634 3023 2658 3024
rect 2637 3025 2851 3026
rect 2643 3027 2698 3028
rect 2672 3029 2836 3030
rect 2673 3031 2799 3032
rect 2676 3033 2685 3034
rect 2621 3035 2686 3036
rect 2678 3037 2758 3038
rect 2679 3039 2784 3040
rect 2682 3041 2787 3042
rect 2502 3043 2786 3044
rect 2690 3045 2892 3046
rect 2691 3047 2845 3048
rect 2703 3049 2733 3050
rect 2709 3051 2790 3052
rect 2711 3053 2789 3054
rect 2712 3055 2793 3056
rect 2733 3057 2821 3058
rect 2736 3059 2749 3060
rect 2738 3061 2913 3062
rect 2739 3063 2827 3064
rect 2754 3065 2842 3066
rect 2760 3067 2863 3068
rect 2763 3069 2778 3070
rect 2772 3071 2872 3072
rect 2775 3073 2875 3074
rect 2781 3075 2796 3076
rect 2801 3075 2885 3076
rect 2826 3077 2919 3078
rect 2829 3079 2939 3080
rect 2726 3081 2830 3082
rect 2714 3083 2728 3084
rect 2859 3083 2932 3084
rect 2062 3092 2191 3093
rect 2065 3094 2375 3095
rect 2087 3096 2278 3097
rect 2097 3098 2290 3099
rect 2079 3100 2099 3101
rect 2101 3100 2305 3101
rect 2104 3102 2126 3103
rect 2110 3104 2401 3105
rect 2115 3106 2395 3107
rect 2073 3108 2396 3109
rect 2114 3110 2314 3111
rect 2120 3112 2155 3113
rect 2123 3114 2158 3115
rect 2126 3116 2347 3117
rect 2135 3118 2177 3119
rect 2138 3120 2209 3121
rect 2142 3122 2263 3123
rect 2141 3124 2306 3125
rect 2145 3126 2443 3127
rect 2157 3128 2179 3129
rect 2173 3130 2282 3131
rect 2182 3132 2215 3133
rect 2202 3134 2369 3135
rect 2218 3136 2245 3137
rect 2224 3138 2356 3139
rect 2232 3140 2363 3141
rect 2236 3142 2386 3143
rect 2238 3144 2383 3145
rect 2241 3146 2473 3147
rect 2242 3148 2269 3149
rect 2263 3150 2287 3151
rect 2269 3152 2311 3153
rect 2138 3154 2312 3155
rect 2283 3156 2411 3157
rect 2293 3158 2329 3159
rect 2296 3160 2332 3161
rect 2317 3162 2359 3163
rect 2083 3164 2360 3165
rect 2329 3166 2335 3167
rect 2335 3168 2341 3169
rect 2338 3170 2344 3171
rect 2341 3172 2371 3173
rect 2347 3174 2365 3175
rect 2365 3176 2380 3177
rect 2371 3178 2377 3179
rect 2383 3178 2407 3179
rect 2072 3180 2408 3181
rect 2389 3182 2392 3183
rect 2112 3184 2393 3185
rect 2397 3184 2402 3185
rect 2076 3186 2399 3187
rect 2075 3188 2272 3189
rect 2403 3188 2414 3189
rect 2094 3190 2405 3191
rect 2094 3192 2273 3193
rect 2422 3192 2479 3193
rect 2428 3194 2446 3195
rect 2436 3196 2444 3197
rect 2424 3198 2438 3199
rect 2439 3198 2447 3199
rect 2448 3198 2651 3199
rect 2160 3200 2450 3201
rect 2466 3200 2474 3201
rect 2460 3202 2468 3203
rect 2454 3204 2462 3205
rect 2430 3206 2456 3207
rect 2131 3208 2432 3209
rect 2479 3208 2654 3209
rect 2490 3210 2719 3211
rect 2287 3212 2492 3213
rect 2496 3212 2731 3213
rect 2484 3214 2498 3215
rect 2502 3214 2697 3215
rect 2503 3216 2509 3217
rect 2521 3216 2713 3217
rect 2524 3218 2569 3219
rect 2532 3220 2540 3221
rect 2536 3222 2551 3223
rect 2542 3224 2545 3225
rect 2553 3224 2821 3225
rect 2554 3226 2581 3227
rect 2556 3228 2712 3229
rect 2560 3230 2563 3231
rect 2572 3230 2632 3231
rect 2574 3232 2661 3233
rect 2575 3234 2635 3235
rect 2578 3236 2670 3237
rect 2590 3238 2801 3239
rect 2592 3240 2847 3241
rect 2593 3242 2611 3243
rect 2595 3244 2840 3245
rect 2475 3246 2597 3247
rect 2469 3248 2477 3249
rect 2598 3248 2837 3249
rect 2322 3250 2600 3251
rect 2323 3252 2353 3253
rect 2128 3254 2354 3255
rect 2129 3256 2435 3257
rect 2602 3256 2833 3257
rect 2604 3258 2804 3259
rect 2613 3260 2721 3261
rect 2620 3262 2686 3263
rect 2623 3264 2644 3265
rect 2632 3266 2807 3267
rect 2635 3268 2824 3269
rect 2641 3270 2683 3271
rect 2644 3272 2742 3273
rect 2663 3274 2704 3275
rect 2666 3276 2707 3277
rect 2673 3278 2778 3279
rect 2676 3280 2810 3281
rect 2675 3282 2788 3283
rect 2681 3284 2818 3285
rect 2684 3286 2814 3287
rect 2688 3288 2701 3289
rect 2702 3288 2792 3289
rect 2709 3290 2785 3291
rect 2708 3292 2734 3293
rect 2723 3294 2749 3295
rect 2726 3296 2755 3297
rect 2729 3298 2758 3299
rect 2732 3300 2761 3301
rect 2514 3302 2760 3303
rect 2515 3304 2638 3305
rect 2638 3306 2680 3307
rect 2736 3306 2752 3307
rect 2735 3308 2764 3309
rect 2739 3310 2767 3311
rect 2691 3312 2739 3313
rect 2690 3314 2781 3315
rect 2750 3316 2773 3317
rect 2526 3318 2774 3319
rect 2753 3320 2776 3321
rect 2797 3320 2827 3321
rect 2011 3329 2339 3330
rect 2065 3331 2396 3332
rect 2068 3333 2268 3334
rect 2068 3335 2399 3336
rect 2072 3337 2139 3338
rect 2079 3339 2390 3340
rect 2082 3341 2388 3342
rect 2094 3343 2264 3344
rect 2098 3345 2253 3346
rect 2108 3347 2121 3348
rect 2114 3349 2262 3350
rect 2041 3351 2115 3352
rect 2117 3351 2273 3352
rect 2117 3353 2124 3354
rect 2120 3355 2310 3356
rect 2126 3357 2324 3358
rect 2127 3359 2219 3360
rect 2129 3361 2149 3362
rect 2141 3363 2286 3364
rect 2166 3365 2393 3366
rect 2153 3367 2394 3368
rect 2157 3369 2166 3370
rect 2156 3371 2586 3372
rect 2171 3373 2369 3374
rect 2173 3375 2297 3376
rect 2174 3377 2664 3378
rect 2176 3379 2288 3380
rect 2177 3381 2183 3382
rect 2207 3381 2450 3382
rect 2224 3383 2235 3384
rect 2225 3385 2243 3386
rect 2228 3387 2411 3388
rect 2210 3389 2412 3390
rect 2239 3391 2358 3392
rect 2243 3393 2366 3394
rect 2258 3395 2270 3396
rect 2104 3397 2271 3398
rect 2279 3397 2294 3398
rect 2291 3399 2306 3400
rect 2297 3401 2312 3402
rect 2303 3403 2318 3404
rect 2312 3405 2330 3406
rect 2324 3407 2342 3408
rect 2330 3409 2348 3410
rect 2339 3411 2354 3412
rect 2345 3413 2360 3414
rect 2351 3415 2384 3416
rect 2362 3417 2391 3418
rect 2363 3419 2438 3420
rect 2369 3421 2372 3422
rect 2372 3423 2375 3424
rect 2375 3425 2402 3426
rect 2087 3427 2403 3428
rect 2378 3429 2405 3430
rect 2396 3431 2429 3432
rect 2399 3433 2414 3434
rect 2405 3435 2408 3436
rect 2075 3437 2409 3438
rect 2429 3437 2432 3438
rect 2432 3439 2435 3440
rect 2435 3441 2462 3442
rect 2441 3443 2492 3444
rect 2446 3445 2451 3446
rect 2443 3447 2448 3448
rect 2453 3447 2468 3448
rect 2455 3449 2651 3450
rect 2465 3451 2670 3452
rect 2471 3453 2474 3454
rect 2474 3455 2477 3456
rect 2240 3457 2478 3458
rect 2482 3457 2502 3458
rect 2483 3459 2697 3460
rect 2489 3461 2597 3462
rect 2492 3463 2600 3464
rect 2495 3465 2712 3466
rect 2497 3467 2613 3468
rect 2507 3469 2724 3470
rect 2515 3471 2661 3472
rect 2521 3473 2529 3474
rect 2542 3473 2550 3474
rect 2543 3475 2573 3476
rect 2546 3477 2576 3478
rect 2554 3479 2738 3480
rect 2539 3481 2556 3482
rect 2560 3481 2568 3482
rect 2578 3481 2658 3482
rect 2593 3483 2607 3484
rect 2609 3483 2667 3484
rect 2503 3485 2668 3486
rect 2422 3487 2505 3488
rect 2423 3489 2480 3490
rect 2620 3489 2658 3490
rect 2623 3491 2649 3492
rect 2627 3493 2781 3494
rect 2519 3495 2781 3496
rect 2630 3497 2636 3498
rect 2632 3499 2778 3500
rect 2633 3501 2639 3502
rect 2636 3503 2642 3504
rect 2639 3505 2741 3506
rect 2644 3507 2833 3508
rect 2645 3509 2661 3510
rect 2675 3509 2696 3510
rect 2702 3509 2714 3510
rect 2701 3511 2812 3512
rect 2720 3513 2805 3514
rect 2726 3515 2744 3516
rect 2725 3517 2760 3518
rect 2729 3519 2747 3520
rect 2708 3521 2729 3522
rect 2690 3523 2708 3524
rect 2750 3523 2762 3524
rect 2732 3525 2750 3526
rect 2753 3525 2765 3526
rect 2735 3527 2753 3528
rect 2734 3529 2788 3530
rect 2767 3531 2808 3532
rect 2684 3533 2809 3534
rect 2773 3535 2785 3536
rect 2264 3537 2774 3538
rect 2674 3539 2784 3540
rect 2797 3539 2839 3540
rect 2677 3541 2798 3542
rect 2817 3541 2826 3542
rect 2814 3543 2819 3544
rect 2731 3545 2816 3546
rect 2038 3554 2226 3555
rect 2044 3556 2109 3557
rect 2052 3558 2060 3559
rect 2056 3560 2346 3561
rect 2066 3562 2271 3563
rect 2072 3564 2430 3565
rect 2068 3566 2074 3567
rect 2084 3566 2391 3567
rect 2084 3568 2200 3569
rect 2094 3570 2403 3571
rect 2102 3572 2379 3573
rect 2105 3574 2221 3575
rect 2106 3576 2376 3577
rect 2110 3578 2253 3579
rect 2114 3580 2124 3581
rect 2117 3582 2127 3583
rect 2117 3584 2278 3585
rect 2130 3586 2290 3587
rect 2129 3588 2656 3589
rect 2132 3590 2235 3591
rect 2134 3592 2254 3593
rect 2137 3594 2484 3595
rect 2139 3596 2292 3597
rect 2146 3598 2377 3599
rect 2184 3600 2283 3601
rect 2087 3602 2284 3603
rect 2190 3604 2229 3605
rect 2192 3606 2436 3607
rect 2196 3608 2268 3609
rect 2205 3610 2337 3611
rect 2207 3612 2368 3613
rect 2165 3614 2209 3615
rect 2217 3614 2356 3615
rect 2223 3616 2259 3617
rect 2229 3618 2340 3619
rect 2235 3620 2370 3621
rect 2238 3622 2373 3623
rect 2177 3624 2374 3625
rect 2178 3626 2451 3627
rect 2241 3628 2433 3629
rect 2243 3630 2454 3631
rect 2250 3632 2388 3633
rect 2256 3634 2310 3635
rect 2261 3636 2293 3637
rect 2262 3638 2406 3639
rect 2268 3640 2400 3641
rect 2279 3642 2455 3643
rect 2285 3644 2344 3645
rect 2120 3646 2287 3647
rect 2120 3648 2302 3649
rect 2295 3650 2298 3651
rect 2307 3650 2448 3651
rect 2312 3652 2320 3653
rect 2303 3654 2314 3655
rect 2324 3654 2536 3655
rect 2330 3656 2524 3657
rect 2331 3658 2397 3659
rect 2334 3660 2394 3661
rect 2337 3662 2472 3663
rect 2349 3664 2478 3665
rect 2351 3666 2458 3667
rect 2357 3668 2542 3669
rect 2361 3670 2412 3671
rect 2379 3672 2668 3673
rect 2385 3674 2520 3675
rect 2397 3676 2538 3677
rect 2403 3678 2424 3679
rect 2424 3680 2529 3681
rect 2439 3682 2496 3683
rect 2174 3684 2497 3685
rect 2175 3686 2452 3687
rect 2463 3686 2738 3687
rect 2465 3688 2586 3689
rect 2474 3690 2560 3691
rect 2487 3692 2613 3693
rect 2499 3694 2604 3695
rect 2501 3696 2599 3697
rect 2502 3698 2607 3699
rect 2504 3700 2602 3701
rect 2363 3702 2506 3703
rect 2507 3702 2512 3703
rect 2529 3702 2671 3703
rect 2543 3704 2690 3705
rect 2546 3706 2590 3707
rect 2549 3708 2777 3709
rect 2553 3710 2753 3711
rect 2555 3712 2687 3713
rect 2571 3714 2592 3715
rect 2583 3716 2634 3717
rect 2586 3718 2693 3719
rect 2604 3720 2640 3721
rect 2627 3722 2662 3723
rect 2628 3724 2665 3725
rect 2630 3726 2779 3727
rect 2631 3728 2658 3729
rect 2636 3730 2819 3731
rect 2427 3732 2819 3733
rect 2640 3734 2646 3735
rect 2489 3736 2647 3737
rect 2441 3738 2491 3739
rect 2643 3738 2649 3739
rect 2492 3740 2650 3741
rect 2264 3742 2494 3743
rect 2265 3744 2409 3745
rect 2409 3746 2753 3747
rect 2658 3748 2809 3749
rect 2673 3750 2717 3751
rect 2677 3752 2684 3753
rect 2609 3754 2678 3755
rect 2610 3756 2735 3757
rect 2680 3758 2802 3759
rect 2695 3760 2759 3761
rect 2701 3762 2816 3763
rect 2707 3764 2812 3765
rect 2707 3766 2774 3767
rect 2710 3768 2714 3769
rect 2713 3770 2729 3771
rect 2722 3772 2726 3773
rect 2734 3772 2791 3773
rect 2737 3774 2747 3775
rect 2743 3776 2788 3777
rect 2421 3778 2788 3779
rect 2743 3780 2768 3781
rect 2481 3782 2769 3783
rect 2746 3784 2771 3785
rect 2755 3786 2762 3787
rect 2567 3788 2762 3789
rect 2764 3788 2784 3789
rect 2680 3790 2765 3791
rect 2749 3792 2785 3793
rect 2525 3794 2750 3795
rect 2781 3794 2812 3795
rect 2815 3794 2833 3795
rect 2038 3803 2124 3804
rect 2042 3805 2127 3806
rect 2059 3807 2236 3808
rect 2068 3809 2226 3810
rect 2077 3811 2230 3812
rect 2087 3813 2251 3814
rect 2089 3815 2217 3816
rect 2091 3817 2113 3818
rect 2100 3819 2284 3820
rect 2124 3821 2340 3822
rect 2129 3823 2242 3824
rect 2072 3825 2241 3826
rect 2132 3827 2259 3828
rect 2139 3829 2314 3830
rect 2120 3831 2313 3832
rect 2141 3833 2356 3834
rect 2172 3835 2599 3836
rect 2175 3837 2335 3838
rect 2174 3839 2179 3840
rect 2180 3839 2239 3840
rect 2184 3841 2338 3842
rect 2187 3843 2263 3844
rect 2192 3845 2497 3846
rect 2196 3847 2235 3848
rect 2075 3849 2196 3850
rect 2199 3849 2211 3850
rect 2198 3851 2209 3852
rect 2205 3853 2238 3854
rect 2190 3855 2205 3856
rect 2214 3855 2530 3856
rect 2228 3857 2455 3858
rect 2246 3859 2374 3860
rect 2268 3861 2298 3862
rect 2080 3863 2268 3864
rect 2079 3865 2221 3866
rect 2271 3865 2560 3866
rect 2265 3867 2271 3868
rect 2274 3867 2517 3868
rect 2273 3869 2344 3870
rect 2277 3871 2310 3872
rect 2279 3873 2287 3874
rect 2256 3875 2286 3876
rect 2289 3875 2316 3876
rect 2295 3877 2304 3878
rect 2253 3879 2295 3880
rect 2223 3881 2253 3882
rect 2301 3881 2346 3882
rect 2094 3883 2301 3884
rect 2093 3885 2223 3886
rect 2307 3885 2334 3886
rect 2319 3887 2322 3888
rect 2292 3889 2319 3890
rect 2117 3891 2292 3892
rect 2327 3891 2350 3892
rect 2348 3893 2377 3894
rect 2351 3895 2536 3896
rect 2354 3897 2494 3898
rect 2357 3899 2452 3900
rect 2372 3901 2458 3902
rect 2385 3903 2728 3904
rect 2390 3905 2765 3906
rect 2397 3907 2816 3908
rect 2396 3909 2404 3910
rect 2379 3911 2403 3912
rect 2409 3911 2618 3912
rect 2414 3913 2602 3914
rect 2417 3915 2506 3916
rect 2424 3917 2750 3918
rect 2429 3919 2753 3920
rect 2432 3921 2687 3922
rect 2427 3923 2687 3924
rect 2421 3925 2427 3926
rect 2439 3925 2772 3926
rect 2438 3927 2464 3928
rect 2456 3929 2491 3930
rect 2462 3931 2656 3932
rect 2474 3933 2503 3934
rect 2492 3935 2512 3936
rect 2499 3937 2514 3938
rect 2481 3939 2499 3940
rect 2480 3941 2524 3942
rect 2510 3943 2802 3944
rect 2528 3945 2629 3946
rect 2531 3947 2632 3948
rect 2534 3949 2587 3950
rect 2537 3951 2572 3952
rect 2487 3953 2571 3954
rect 2486 3955 2542 3956
rect 2543 3955 2641 3956
rect 2546 3957 2602 3958
rect 2549 3959 2554 3960
rect 2567 3959 2678 3960
rect 2573 3961 2605 3962
rect 2583 3963 2693 3964
rect 2585 3965 2647 3966
rect 2589 3967 2690 3968
rect 2588 3969 2650 3970
rect 2604 3971 2812 3972
rect 2610 3973 2669 3974
rect 2610 3975 2735 3976
rect 2331 3977 2735 3978
rect 2623 3979 2659 3980
rect 2626 3981 2662 3982
rect 2643 3983 2674 3984
rect 2647 3985 2708 3986
rect 2650 3987 2711 3988
rect 2653 3989 2721 3990
rect 2665 3991 2732 3992
rect 2450 3993 2731 3994
rect 2683 3995 2809 3996
rect 2683 3997 2744 3998
rect 2689 3999 2795 4000
rect 2695 4001 2776 4002
rect 2701 4003 2756 4004
rect 2704 4005 2759 4006
rect 2707 4007 2714 4008
rect 2710 4009 2717 4010
rect 2635 4011 2717 4012
rect 2737 4011 2764 4012
rect 2740 4013 2782 4014
rect 2743 4015 2785 4016
rect 2746 4017 2788 4018
rect 2698 4019 2747 4020
rect 2056 4028 2268 4029
rect 2082 4030 2286 4031
rect 2083 4032 2292 4033
rect 2087 4034 2164 4035
rect 2089 4036 2301 4037
rect 2097 4038 2128 4039
rect 2100 4040 2386 4041
rect 2103 4042 2319 4043
rect 2104 4044 2313 4045
rect 2079 4046 2314 4047
rect 2080 4048 2095 4049
rect 2112 4048 2371 4049
rect 2119 4050 2316 4051
rect 2122 4052 2344 4053
rect 2129 4054 2223 4055
rect 2131 4056 2304 4057
rect 2133 4058 2247 4059
rect 2138 4060 2340 4061
rect 2141 4062 2346 4063
rect 2148 4064 2341 4065
rect 2157 4066 2194 4067
rect 2189 4068 2266 4069
rect 2068 4070 2191 4071
rect 2198 4070 2203 4071
rect 2195 4072 2200 4073
rect 2204 4072 2209 4073
rect 2210 4072 2215 4073
rect 2216 4072 2221 4073
rect 2225 4072 2389 4073
rect 2226 4074 2547 4075
rect 2228 4076 2305 4077
rect 2231 4078 2358 4079
rect 2234 4080 2269 4081
rect 2237 4082 2302 4083
rect 2240 4084 2245 4085
rect 2252 4084 2347 4085
rect 2256 4086 2422 4087
rect 2258 4088 2407 4089
rect 2261 4090 2481 4091
rect 2262 4092 2355 4093
rect 2076 4094 2356 4095
rect 2270 4096 2359 4097
rect 2271 4098 2274 4099
rect 2277 4098 2322 4099
rect 2279 4100 2377 4101
rect 2294 4102 2317 4103
rect 2295 4104 2487 4105
rect 2319 4106 2373 4107
rect 2309 4108 2374 4109
rect 2325 4110 2517 4111
rect 2330 4112 2584 4113
rect 2331 4114 2418 4115
rect 2337 4116 2352 4117
rect 2348 4118 2419 4119
rect 2360 4120 2380 4121
rect 2366 4122 2595 4123
rect 2297 4124 2368 4125
rect 2390 4124 2479 4125
rect 2391 4126 2529 4127
rect 2394 4128 2532 4129
rect 2396 4130 2410 4131
rect 2402 4132 2491 4133
rect 2126 4134 2404 4135
rect 2429 4134 2503 4135
rect 2438 4136 2611 4137
rect 2450 4138 2521 4139
rect 2451 4140 2544 4141
rect 2454 4142 2535 4143
rect 2460 4144 2568 4145
rect 2466 4146 2586 4147
rect 2414 4148 2587 4149
rect 2333 4150 2416 4151
rect 2469 4150 2589 4151
rect 2492 4152 2719 4153
rect 2508 4154 2731 4155
rect 2505 4156 2732 4157
rect 2510 4158 2569 4159
rect 2513 4160 2774 4161
rect 2432 4162 2515 4163
rect 2433 4164 2638 4165
rect 2537 4166 2545 4167
rect 2462 4168 2539 4169
rect 2463 4170 2571 4171
rect 2474 4172 2572 4173
rect 2549 4174 2596 4175
rect 2550 4176 2574 4177
rect 2498 4178 2575 4179
rect 2426 4180 2500 4181
rect 2427 4182 2457 4183
rect 2457 4184 2618 4185
rect 2562 4186 2669 4187
rect 2580 4188 2693 4189
rect 2598 4190 2614 4191
rect 2238 4192 2614 4193
rect 2601 4194 2782 4195
rect 2623 4196 2756 4197
rect 2445 4198 2623 4199
rect 2643 4198 2754 4199
rect 2647 4200 2674 4201
rect 2646 4202 2768 4203
rect 2650 4204 2728 4205
rect 2653 4206 2714 4207
rect 2652 4208 2677 4209
rect 2655 4210 2725 4211
rect 2679 4212 2744 4213
rect 2689 4214 2761 4215
rect 2691 4216 2708 4217
rect 2695 4218 2750 4219
rect 2526 4220 2749 4221
rect 2635 4222 2695 4223
rect 2701 4222 2722 4223
rect 2686 4224 2701 4225
rect 2704 4224 2778 4225
rect 2665 4226 2704 4227
rect 2710 4226 2717 4227
rect 2484 4228 2716 4229
rect 2698 4230 2710 4231
rect 2683 4232 2698 4233
rect 2604 4234 2683 4235
rect 2712 4234 2735 4235
rect 2626 4236 2735 4237
rect 2740 4236 2781 4237
rect 2706 4238 2742 4239
rect 2044 4247 2191 4248
rect 2059 4249 2088 4250
rect 2063 4251 2269 4252
rect 2067 4253 2200 4254
rect 2069 4255 2207 4256
rect 2074 4257 2234 4258
rect 2076 4259 2084 4260
rect 2084 4261 2294 4262
rect 2095 4263 2366 4264
rect 2097 4265 2389 4266
rect 2098 4267 2404 4268
rect 2104 4269 2312 4270
rect 2107 4271 2117 4272
rect 2113 4273 2374 4274
rect 2129 4275 2354 4276
rect 2133 4277 2416 4278
rect 2135 4279 2276 4280
rect 2142 4281 2203 4282
rect 2070 4283 2204 4284
rect 2148 4285 2272 4286
rect 2157 4287 2317 4288
rect 2160 4289 2266 4290
rect 2163 4291 2318 4292
rect 2166 4293 2285 4294
rect 2181 4295 2189 4296
rect 2193 4295 2227 4296
rect 2214 4297 2228 4298
rect 2215 4299 2221 4300
rect 2208 4301 2222 4302
rect 2238 4301 2326 4302
rect 2244 4303 2255 4304
rect 2245 4305 2302 4306
rect 2248 4307 2627 4308
rect 2256 4309 2371 4310
rect 2241 4311 2372 4312
rect 2119 4313 2243 4314
rect 2272 4313 2407 4314
rect 2290 4315 2314 4316
rect 2299 4317 2419 4318
rect 2302 4319 2356 4320
rect 2308 4321 2377 4322
rect 2314 4323 2368 4324
rect 2326 4325 2386 4326
rect 2323 4327 2387 4328
rect 2335 4329 2344 4330
rect 2340 4331 2357 4332
rect 2304 4333 2342 4334
rect 2305 4335 2359 4336
rect 2319 4337 2360 4338
rect 2262 4339 2321 4340
rect 2368 4339 2719 4340
rect 2377 4341 2446 4342
rect 2389 4343 2410 4344
rect 2401 4345 2587 4346
rect 2413 4347 2479 4348
rect 2419 4349 2485 4350
rect 2425 4351 2491 4352
rect 2427 4353 2638 4354
rect 2433 4355 2438 4356
rect 2449 4355 2515 4356
rect 2451 4357 2531 4358
rect 2457 4359 2620 4360
rect 2229 4361 2621 4362
rect 2463 4363 2641 4364
rect 2466 4365 2618 4366
rect 2469 4367 2519 4368
rect 2491 4369 2797 4370
rect 2497 4371 2685 4372
rect 2508 4373 2513 4374
rect 2509 4375 2572 4376
rect 2520 4377 2746 4378
rect 2421 4379 2746 4380
rect 2533 4381 2575 4382
rect 2542 4383 2653 4384
rect 2550 4385 2606 4386
rect 2544 4387 2552 4388
rect 2545 4389 2650 4390
rect 2460 4391 2651 4392
rect 2295 4393 2462 4394
rect 2277 4395 2297 4396
rect 2562 4395 2600 4396
rect 2563 4397 2596 4398
rect 2568 4399 2774 4400
rect 2569 4401 2581 4402
rect 2394 4403 2582 4404
rect 2331 4405 2396 4406
rect 2575 4405 2602 4406
rect 2587 4407 2688 4408
rect 2593 4409 2739 4410
rect 2610 4411 2623 4412
rect 2583 4413 2624 4414
rect 2391 4415 2585 4416
rect 2613 4415 2669 4416
rect 2646 4417 2756 4418
rect 2647 4419 2735 4420
rect 2655 4421 2666 4422
rect 2673 4421 2728 4422
rect 2676 4423 2725 4424
rect 2526 4425 2724 4426
rect 2694 4427 2742 4428
rect 2499 4429 2743 4430
rect 2500 4431 2506 4432
rect 2682 4431 2694 4432
rect 2703 4431 2727 4432
rect 2702 4433 2786 4434
rect 2706 4435 2730 4436
rect 2643 4437 2706 4438
rect 2712 4437 2757 4438
rect 2700 4439 2712 4440
rect 2699 4441 2716 4442
rect 2278 4443 2715 4444
rect 2762 4443 2767 4444
rect 2731 4445 2764 4446
rect 2721 4447 2733 4448
rect 2709 4449 2721 4450
rect 2697 4451 2709 4452
rect 2691 4453 2697 4454
rect 2679 4455 2691 4456
rect 2379 4457 2681 4458
rect 2769 4457 2788 4458
rect 2769 4459 2777 4460
rect 2772 4461 2783 4462
rect 2053 4470 2061 4471
rect 2056 4472 2189 4473
rect 2063 4474 2200 4475
rect 2070 4476 2207 4477
rect 2074 4478 2228 4479
rect 2074 4480 2300 4481
rect 2077 4482 2222 4483
rect 2081 4484 2194 4485
rect 2084 4486 2273 4487
rect 2088 4488 2312 4489
rect 2088 4490 2206 4491
rect 2091 4492 2336 4493
rect 2095 4494 2303 4495
rect 2098 4496 2255 4497
rect 2100 4498 2108 4499
rect 2113 4498 2136 4499
rect 2113 4500 2318 4501
rect 2116 4502 2297 4503
rect 2120 4504 2309 4505
rect 2123 4506 2257 4507
rect 2123 4508 2291 4509
rect 2133 4510 2158 4511
rect 2142 4512 2177 4513
rect 2151 4514 2357 4515
rect 2157 4516 2204 4517
rect 2160 4518 2246 4519
rect 2163 4520 2354 4521
rect 2166 4522 2252 4523
rect 2166 4524 2234 4525
rect 2169 4526 2306 4527
rect 2173 4528 2285 4529
rect 2184 4530 2276 4531
rect 2187 4532 2372 4533
rect 2190 4534 2272 4535
rect 2196 4536 2294 4537
rect 2202 4538 2339 4539
rect 2211 4540 2284 4541
rect 2215 4542 2221 4543
rect 2217 4544 2315 4545
rect 2229 4546 2279 4547
rect 2235 4548 2327 4549
rect 2238 4550 2321 4551
rect 2242 4552 2630 4553
rect 2241 4554 2324 4555
rect 2250 4556 2685 4557
rect 2253 4558 2348 4559
rect 2259 4560 2342 4561
rect 2265 4562 2366 4563
rect 2274 4564 2369 4565
rect 2277 4566 2360 4567
rect 2289 4568 2387 4569
rect 2295 4570 2390 4571
rect 2307 4572 2750 4573
rect 2313 4574 2688 4575
rect 2325 4576 2414 4577
rect 2331 4578 2681 4579
rect 2343 4580 2700 4581
rect 2349 4582 2462 4583
rect 2355 4584 2438 4585
rect 2361 4586 2450 4587
rect 2367 4588 2456 4589
rect 2377 4590 2384 4591
rect 2379 4592 2712 4593
rect 2385 4594 2746 4595
rect 2397 4596 2724 4597
rect 2401 4598 2642 4599
rect 2409 4600 2492 4601
rect 2415 4602 2504 4603
rect 2419 4604 2609 4605
rect 2433 4606 2498 4607
rect 2436 4608 2501 4609
rect 2445 4610 2582 4611
rect 2301 4612 2581 4613
rect 2448 4614 2585 4615
rect 2451 4616 2534 4617
rect 2457 4618 2531 4619
rect 2460 4620 2680 4621
rect 2463 4622 2540 4623
rect 2466 4624 2543 4625
rect 2469 4626 2552 4627
rect 2475 4628 2546 4629
rect 2395 4630 2545 4631
rect 2478 4632 2513 4633
rect 2487 4634 2618 4635
rect 2490 4636 2621 4637
rect 2493 4638 2564 4639
rect 2499 4640 2570 4641
rect 2505 4642 2594 4643
rect 2509 4644 2539 4645
rect 2511 4646 2716 4647
rect 2518 4648 2806 4649
rect 2523 4650 2600 4651
rect 2529 4652 2760 4653
rect 2535 4654 2790 4655
rect 2541 4656 2548 4657
rect 2550 4656 2624 4657
rect 2568 4658 2651 4659
rect 2583 4660 2666 4661
rect 2425 4662 2666 4663
rect 2589 4664 2730 4665
rect 2575 4666 2730 4667
rect 2601 4668 2648 4669
rect 2605 4670 2736 4671
rect 2565 4672 2605 4673
rect 2614 4672 2691 4673
rect 2617 4674 2694 4675
rect 2620 4676 2697 4677
rect 2626 4678 2645 4679
rect 2626 4680 2721 4681
rect 2638 4682 2800 4683
rect 2641 4684 2709 4685
rect 2650 4686 2733 4687
rect 2659 4688 2786 4689
rect 2662 4690 2727 4691
rect 2672 4692 2706 4693
rect 2699 4694 2770 4695
rect 2702 4696 2767 4697
rect 2587 4698 2703 4699
rect 2586 4700 2669 4701
rect 2623 4702 2669 4703
rect 2705 4702 2773 4703
rect 2060 4711 2226 4712
rect 2074 4713 2192 4714
rect 2077 4715 2189 4716
rect 2081 4717 2167 4718
rect 2093 4719 2101 4720
rect 2106 4719 2236 4720
rect 2084 4721 2106 4722
rect 2084 4723 2134 4724
rect 2109 4725 2235 4726
rect 2108 4727 2126 4728
rect 2113 4729 2142 4730
rect 2116 4731 2158 4732
rect 2130 4733 2290 4734
rect 2138 4735 2208 4736
rect 2151 4737 2296 4738
rect 2152 4739 2185 4740
rect 2154 4741 2467 4742
rect 2158 4743 2170 4744
rect 2164 4745 2242 4746
rect 2067 4747 2241 4748
rect 2067 4749 2183 4750
rect 2193 4749 2244 4750
rect 2167 4751 2195 4752
rect 2196 4751 2247 4752
rect 2211 4753 2621 4754
rect 2214 4755 2651 4756
rect 2217 4757 2262 4758
rect 2229 4759 2289 4760
rect 2202 4761 2229 4762
rect 2238 4761 2286 4762
rect 2199 4763 2238 4764
rect 2253 4763 2304 4764
rect 2112 4765 2253 4766
rect 2256 4765 2298 4766
rect 2205 4767 2256 4768
rect 2259 4767 2581 4768
rect 2265 4769 2319 4770
rect 2220 4771 2265 4772
rect 2063 4773 2220 4774
rect 2274 4773 2322 4774
rect 2279 4775 2644 4776
rect 2283 4777 2551 4778
rect 2309 4779 2491 4780
rect 2325 4781 2648 4782
rect 2277 4783 2325 4784
rect 2331 4783 2373 4784
rect 2330 4785 2350 4786
rect 2313 4787 2349 4788
rect 2271 4789 2313 4790
rect 2343 4789 2716 4790
rect 2307 4791 2343 4792
rect 2361 4791 2391 4792
rect 2367 4793 2403 4794
rect 2397 4795 2713 4796
rect 2415 4797 2430 4798
rect 2379 4799 2415 4800
rect 2355 4801 2379 4802
rect 2301 4803 2355 4804
rect 2250 4805 2301 4806
rect 2120 4807 2250 4808
rect 2417 4807 2446 4808
rect 2420 4809 2449 4810
rect 2436 4811 2439 4812
rect 2433 4813 2436 4814
rect 2441 4813 2458 4814
rect 2444 4815 2461 4816
rect 2451 4817 2466 4818
rect 2453 4819 2479 4820
rect 2459 4821 2464 4822
rect 2462 4823 2578 4824
rect 2469 4825 2478 4826
rect 2471 4827 2569 4828
rect 2475 4829 2484 4830
rect 2487 4829 2508 4830
rect 2493 4831 2577 4832
rect 2495 4833 2669 4834
rect 2499 4835 2520 4836
rect 2505 4837 2514 4838
rect 2511 4839 2532 4840
rect 2306 4841 2511 4842
rect 2523 4841 2709 4842
rect 2529 4843 2694 4844
rect 2535 4845 2556 4846
rect 2538 4847 2559 4848
rect 2544 4849 2613 4850
rect 2543 4851 2548 4852
rect 2541 4853 2547 4854
rect 2567 4853 2630 4854
rect 2573 4855 2618 4856
rect 2579 4857 2605 4858
rect 2589 4859 2595 4860
rect 2586 4861 2589 4862
rect 2583 4863 2586 4864
rect 2565 4865 2583 4866
rect 2591 4865 2709 4866
rect 2606 4867 2624 4868
rect 2360 4869 2625 4870
rect 2614 4871 2730 4872
rect 2618 4873 2697 4874
rect 2626 4875 2653 4876
rect 2636 4877 2673 4878
rect 2498 4879 2674 4880
rect 2638 4881 2737 4882
rect 2641 4883 2734 4884
rect 2409 4885 2735 4886
rect 2385 4887 2409 4888
rect 2649 4887 2695 4888
rect 2659 4889 2668 4890
rect 2609 4891 2659 4892
rect 2662 4891 2688 4892
rect 2670 4893 2691 4894
rect 2699 4893 2715 4894
rect 2702 4895 2718 4896
rect 2726 4895 2738 4896
rect 2053 4904 2226 4905
rect 2060 4906 2241 4907
rect 2063 4908 2165 4909
rect 2066 4910 2189 4911
rect 2070 4912 2238 4913
rect 2069 4914 2082 4915
rect 2074 4916 2183 4917
rect 2077 4918 2192 4919
rect 2076 4920 2081 4921
rect 2083 4920 2201 4921
rect 2095 4922 2247 4923
rect 2105 4924 2235 4925
rect 2108 4926 2265 4927
rect 2115 4928 2256 4929
rect 2119 4930 2235 4931
rect 2122 4932 2244 4933
rect 2125 4934 2139 4935
rect 2134 4936 2208 4937
rect 2135 4938 2159 4939
rect 2141 4940 2152 4941
rect 2141 4942 2397 4943
rect 2155 4944 2325 4945
rect 2155 4946 2286 4947
rect 2158 4948 2280 4949
rect 2161 4950 2220 4951
rect 2170 4952 2217 4953
rect 2179 4954 2229 4955
rect 2185 4956 2250 4957
rect 2188 4958 2253 4959
rect 2197 4960 2388 4961
rect 2197 4962 2262 4963
rect 2204 4964 2580 4965
rect 2222 4966 2289 4967
rect 2231 4968 2298 4969
rect 2243 4970 2301 4971
rect 2246 4972 2304 4973
rect 2255 4974 2319 4975
rect 2261 4976 2331 4977
rect 2273 4978 2361 4979
rect 2279 4980 2616 4981
rect 2285 4982 2349 4983
rect 2303 4984 2373 4985
rect 2309 4986 2379 4987
rect 2315 4988 2600 4989
rect 2321 4990 2400 4991
rect 2321 4992 2391 4993
rect 2327 4994 2445 4995
rect 2342 4996 2550 4997
rect 2345 4998 2409 4999
rect 2351 5000 2415 5001
rect 2354 5002 2581 5003
rect 2366 5004 2430 5005
rect 2372 5006 2436 5007
rect 2375 5008 2439 5009
rect 2378 5010 2617 5011
rect 2384 5012 2559 5013
rect 2390 5014 2460 5015
rect 2393 5016 2681 5017
rect 2402 5018 2738 5019
rect 2408 5020 2478 5021
rect 2432 5022 2496 5023
rect 2435 5024 2499 5025
rect 2438 5026 2577 5027
rect 2441 5028 2445 5029
rect 2441 5030 2466 5031
rect 2420 5032 2466 5033
rect 2420 5034 2484 5035
rect 2447 5036 2553 5037
rect 2453 5038 2702 5039
rect 2456 5040 2520 5041
rect 2462 5042 2647 5043
rect 2417 5044 2463 5045
rect 2468 5044 2728 5045
rect 2471 5046 2520 5047
rect 2474 5048 2532 5049
rect 2486 5050 2508 5051
rect 2297 5052 2508 5053
rect 2489 5054 2511 5055
rect 2492 5056 2547 5057
rect 2495 5058 2572 5059
rect 2510 5060 2568 5061
rect 2513 5062 2625 5063
rect 2516 5064 2583 5065
rect 2522 5066 2586 5067
rect 2525 5068 2589 5069
rect 2528 5070 2592 5071
rect 2531 5072 2621 5073
rect 2546 5074 2610 5075
rect 2555 5076 2643 5077
rect 2543 5078 2557 5079
rect 2312 5080 2544 5081
rect 2562 5080 2619 5081
rect 2565 5082 2595 5083
rect 2586 5084 2650 5085
rect 2589 5086 2653 5087
rect 2592 5088 2671 5089
rect 2606 5090 2656 5091
rect 2573 5092 2607 5093
rect 2627 5092 2640 5093
rect 2626 5094 2721 5095
rect 2629 5096 2718 5097
rect 2667 5098 2691 5099
rect 2714 5098 2724 5099
rect 2054 5107 2162 5108
rect 2057 5109 2120 5110
rect 2062 5111 2165 5112
rect 2071 5113 2136 5114
rect 2078 5115 2093 5116
rect 2081 5117 2096 5118
rect 2098 5117 2201 5118
rect 2101 5119 2198 5120
rect 2102 5121 2115 5122
rect 2105 5123 2132 5124
rect 2111 5125 2186 5126
rect 2122 5127 2139 5128
rect 2126 5129 2145 5130
rect 2128 5131 2276 5132
rect 2137 5133 2152 5134
rect 2141 5135 2235 5136
rect 2144 5137 2517 5138
rect 2155 5139 2587 5140
rect 2167 5141 2400 5142
rect 2167 5143 2180 5144
rect 2170 5145 2397 5146
rect 2170 5147 2189 5148
rect 2191 5147 2223 5148
rect 2200 5149 2232 5150
rect 2203 5151 2244 5152
rect 2206 5153 2247 5154
rect 2210 5155 2282 5156
rect 2148 5157 2210 5158
rect 2216 5157 2219 5158
rect 2215 5159 2256 5160
rect 2221 5161 2262 5162
rect 2233 5163 2280 5164
rect 2236 5165 2466 5166
rect 2254 5167 2304 5168
rect 2260 5169 2328 5170
rect 2266 5171 2603 5172
rect 2273 5173 2553 5174
rect 2272 5175 2463 5176
rect 2278 5177 2487 5178
rect 2290 5179 2322 5180
rect 2297 5181 2541 5182
rect 2296 5183 2596 5184
rect 2302 5185 2346 5186
rect 2309 5187 2572 5188
rect 2308 5189 2569 5190
rect 2329 5191 2385 5192
rect 2338 5193 2607 5194
rect 2344 5195 2388 5196
rect 2347 5197 2445 5198
rect 2359 5199 2433 5200
rect 2362 5201 2367 5202
rect 2372 5201 2498 5202
rect 2371 5203 2593 5204
rect 2375 5205 2486 5206
rect 2285 5207 2375 5208
rect 2284 5209 2316 5210
rect 2314 5211 2352 5212
rect 2350 5213 2448 5214
rect 2378 5215 2610 5216
rect 2377 5217 2457 5218
rect 2383 5219 2439 5220
rect 2386 5221 2458 5222
rect 2390 5223 2557 5224
rect 2393 5225 2425 5226
rect 2392 5227 2643 5228
rect 2408 5229 2434 5230
rect 2410 5231 2550 5232
rect 2420 5233 2516 5234
rect 2257 5235 2421 5236
rect 2430 5235 2523 5236
rect 2441 5237 2544 5238
rect 2442 5239 2547 5240
rect 2445 5241 2461 5242
rect 2454 5243 2529 5244
rect 2464 5245 2526 5246
rect 2468 5247 2530 5248
rect 2470 5249 2563 5250
rect 2476 5251 2633 5252
rect 2479 5253 2630 5254
rect 2489 5255 2505 5256
rect 2488 5257 2590 5258
rect 2495 5259 2508 5260
rect 2492 5261 2495 5262
rect 2491 5263 2511 5264
rect 2482 5265 2512 5266
rect 2519 5265 2537 5266
rect 2435 5267 2519 5268
rect 2531 5267 2614 5268
rect 2474 5269 2533 5270
rect 2473 5271 2566 5272
rect 2620 5271 2627 5272
rect 2047 5280 2120 5281
rect 2074 5282 2093 5283
rect 2075 5284 2123 5285
rect 2079 5286 2086 5287
rect 2082 5288 2090 5289
rect 2092 5288 2100 5289
rect 2102 5288 2171 5289
rect 2106 5290 2219 5291
rect 2113 5292 2135 5293
rect 2116 5294 2197 5295
rect 2119 5296 2152 5297
rect 2122 5298 2129 5299
rect 2128 5300 2132 5301
rect 2131 5302 2142 5303
rect 2138 5304 2227 5305
rect 2148 5306 2164 5307
rect 2155 5308 2222 5309
rect 2157 5310 2273 5311
rect 2167 5312 2176 5313
rect 2169 5314 2210 5315
rect 2203 5316 2209 5317
rect 2206 5318 2212 5319
rect 2215 5318 2224 5319
rect 2200 5320 2215 5321
rect 2191 5322 2200 5323
rect 2217 5322 2248 5323
rect 2229 5324 2279 5325
rect 2233 5326 2245 5327
rect 2238 5328 2276 5329
rect 2241 5330 2282 5331
rect 2254 5332 2287 5333
rect 2257 5334 2509 5335
rect 2260 5336 2411 5337
rect 2259 5338 2375 5339
rect 2266 5340 2278 5341
rect 2265 5342 2351 5343
rect 2271 5344 2403 5345
rect 2296 5346 2332 5347
rect 2302 5348 2547 5349
rect 2308 5350 2335 5351
rect 2290 5352 2308 5353
rect 2289 5354 2512 5355
rect 2314 5356 2523 5357
rect 2319 5358 2399 5359
rect 2322 5360 2348 5361
rect 2325 5362 2363 5363
rect 2338 5364 2341 5365
rect 2344 5364 2353 5365
rect 2359 5364 2516 5365
rect 2368 5366 2418 5367
rect 2367 5368 2461 5369
rect 2371 5370 2380 5371
rect 2370 5372 2446 5373
rect 2386 5374 2526 5375
rect 2383 5376 2386 5377
rect 2382 5378 2396 5379
rect 2388 5380 2443 5381
rect 2392 5382 2530 5383
rect 2414 5384 2431 5385
rect 2417 5386 2434 5387
rect 2420 5388 2477 5389
rect 2313 5390 2421 5391
rect 2427 5390 2443 5391
rect 2430 5392 2483 5393
rect 2329 5394 2483 5395
rect 2328 5396 2486 5397
rect 2433 5398 2471 5399
rect 2436 5400 2502 5401
rect 2445 5402 2489 5403
rect 2448 5404 2492 5405
rect 2454 5406 2466 5407
rect 2473 5406 2537 5407
rect 2284 5408 2473 5409
rect 2283 5410 2425 5411
rect 2377 5412 2424 5413
rect 2479 5412 2533 5413
rect 2491 5414 2501 5415
rect 2494 5416 2498 5417
rect 2065 5425 2073 5426
rect 2079 5425 2129 5426
rect 2099 5427 2114 5428
rect 2106 5429 2173 5430
rect 2111 5431 2179 5432
rect 2115 5433 2215 5434
rect 2119 5435 2182 5436
rect 2125 5437 2252 5438
rect 2127 5439 2209 5440
rect 2131 5441 2221 5442
rect 2130 5443 2212 5444
rect 2141 5445 2233 5446
rect 2145 5447 2158 5448
rect 2138 5449 2145 5450
rect 2148 5449 2242 5450
rect 2151 5451 2258 5452
rect 2163 5453 2167 5454
rect 2175 5453 2206 5454
rect 2196 5455 2222 5456
rect 2118 5457 2197 5458
rect 2223 5457 2255 5458
rect 2199 5459 2225 5460
rect 2184 5461 2200 5462
rect 2169 5463 2185 5464
rect 2229 5463 2306 5464
rect 2238 5465 2276 5466
rect 2247 5467 2266 5468
rect 2248 5469 2323 5470
rect 2134 5471 2324 5472
rect 2259 5473 2469 5474
rect 2260 5475 2383 5476
rect 2218 5477 2384 5478
rect 2277 5479 2339 5480
rect 2215 5481 2279 5482
rect 2283 5481 2392 5482
rect 2284 5483 2360 5484
rect 2286 5485 2297 5486
rect 2287 5487 2314 5488
rect 2289 5489 2420 5490
rect 2307 5491 2455 5492
rect 2244 5493 2309 5494
rect 2245 5495 2320 5496
rect 2317 5497 2390 5498
rect 2328 5499 2411 5500
rect 2271 5501 2330 5502
rect 2235 5503 2273 5504
rect 2347 5503 2424 5504
rect 2352 5505 2405 5506
rect 2370 5507 2403 5508
rect 2374 5509 2418 5510
rect 2379 5511 2396 5512
rect 2380 5513 2439 5514
rect 2385 5515 2484 5516
rect 2365 5517 2387 5518
rect 2407 5517 2431 5518
rect 2340 5519 2432 5520
rect 2341 5521 2423 5522
rect 2414 5523 2456 5524
rect 2413 5525 2434 5526
rect 2353 5527 2435 5528
rect 2416 5529 2437 5530
rect 2425 5531 2453 5532
rect 2428 5533 2446 5534
rect 2367 5535 2446 5536
rect 2441 5537 2449 5538
rect 2325 5539 2449 5540
rect 2326 5541 2399 5542
rect 2331 5543 2399 5544
rect 2476 5543 2495 5544
rect 2487 5545 2495 5546
rect 2491 5547 2515 5548
rect 2500 5549 2505 5550
rect 2089 5558 2193 5559
rect 2092 5560 2190 5561
rect 2101 5562 2206 5563
rect 2111 5564 2173 5565
rect 2104 5566 2112 5567
rect 2118 5566 2197 5567
rect 2132 5568 2154 5569
rect 2134 5570 2249 5571
rect 2137 5572 2222 5573
rect 2141 5574 2279 5575
rect 2148 5576 2273 5577
rect 2159 5578 2200 5579
rect 2162 5580 2185 5581
rect 2166 5582 2223 5583
rect 2171 5584 2179 5585
rect 2174 5586 2182 5587
rect 2183 5586 2258 5587
rect 2195 5588 2212 5589
rect 2198 5590 2439 5591
rect 2204 5592 2225 5593
rect 2208 5594 2327 5595
rect 2144 5596 2208 5597
rect 2216 5596 2228 5597
rect 2225 5598 2276 5599
rect 2228 5600 2255 5601
rect 2231 5602 2242 5603
rect 2233 5604 2290 5605
rect 2234 5606 2252 5607
rect 2236 5608 2293 5609
rect 2237 5610 2263 5611
rect 2247 5612 2306 5613
rect 2245 5614 2305 5615
rect 2284 5616 2324 5617
rect 2283 5618 2339 5619
rect 2287 5620 2318 5621
rect 2286 5622 2330 5623
rect 2296 5624 2299 5625
rect 2260 5626 2296 5627
rect 2259 5628 2309 5629
rect 2307 5630 2366 5631
rect 2310 5632 2420 5633
rect 2322 5634 2449 5635
rect 2325 5636 2342 5637
rect 2335 5638 2366 5639
rect 2340 5640 2345 5641
rect 2347 5640 2394 5641
rect 2350 5642 2417 5643
rect 2353 5644 2401 5645
rect 2356 5646 2384 5647
rect 2359 5648 2379 5649
rect 2359 5650 2375 5651
rect 2369 5652 2381 5653
rect 2372 5654 2388 5655
rect 2375 5656 2408 5657
rect 2390 5658 2414 5659
rect 2404 5660 2488 5661
rect 2406 5662 2426 5663
rect 2410 5664 2446 5665
rect 2428 5666 2442 5667
rect 2473 5666 2484 5667
rect 2089 5675 2193 5676
rect 2092 5677 2100 5678
rect 2104 5677 2172 5678
rect 2096 5679 2104 5680
rect 2106 5679 2217 5680
rect 2108 5681 2175 5682
rect 2109 5683 2190 5684
rect 2115 5685 2123 5686
rect 2118 5687 2196 5688
rect 2125 5689 2154 5690
rect 2126 5691 2205 5692
rect 2129 5693 2208 5694
rect 2138 5695 2199 5696
rect 2141 5697 2184 5698
rect 2132 5699 2142 5700
rect 2144 5699 2232 5700
rect 2144 5701 2229 5702
rect 2151 5703 2191 5704
rect 2154 5705 2226 5706
rect 2157 5707 2260 5708
rect 2163 5709 2263 5710
rect 2172 5711 2290 5712
rect 2181 5713 2296 5714
rect 2184 5715 2299 5716
rect 2193 5717 2363 5718
rect 2196 5719 2284 5720
rect 2205 5721 2293 5722
rect 2208 5723 2248 5724
rect 2211 5725 2360 5726
rect 2222 5727 2401 5728
rect 2221 5729 2323 5730
rect 2228 5731 2326 5732
rect 2234 5733 2376 5734
rect 2237 5735 2379 5736
rect 2244 5737 2305 5738
rect 2246 5739 2397 5740
rect 2249 5741 2388 5742
rect 2255 5743 2311 5744
rect 2262 5745 2391 5746
rect 2286 5747 2341 5748
rect 2307 5749 2414 5750
rect 2350 5751 2394 5752
rect 2356 5753 2370 5754
rect 2065 5762 2073 5763
rect 2089 5762 2110 5763
rect 2119 5762 2142 5763
rect 2122 5764 2158 5765
rect 2126 5766 2139 5767
rect 2147 5766 2152 5767
rect 2153 5766 2157 5767
rect 2159 5766 2235 5767
rect 2166 5768 2182 5769
rect 2169 5770 2215 5771
rect 2172 5772 2191 5773
rect 2184 5774 2222 5775
rect 2193 5776 2209 5777
rect 2196 5778 2225 5779
rect 2211 5780 2232 5781
rect 2237 5780 2256 5781
rect 2246 5782 2263 5783
rect 2249 5784 2260 5785
rect 2146 5793 2151 5794
rect 2156 5793 2160 5794
rect 2143 5802 2154 5803
<< metal2 >>
rect 2134 1007 2135 1011
rect 2137 1007 2138 1011
rect 2077 1017 2078 1054
rect 2147 1017 2148 1054
rect 2087 1019 2088 1054
rect 2120 1019 2121 1054
rect 2101 1021 2102 1054
rect 2129 1021 2130 1054
rect 2108 1023 2109 1054
rect 2111 1023 2112 1054
rect 2131 1015 2132 1024
rect 2174 1023 2175 1054
rect 2091 1025 2092 1054
rect 2132 1025 2133 1054
rect 2134 1015 2135 1026
rect 2198 1025 2199 1054
rect 2135 1027 2136 1054
rect 2207 1027 2208 1054
rect 2137 1015 2138 1030
rect 2183 1029 2184 1054
rect 2138 1031 2139 1054
rect 2159 1031 2160 1054
rect 2140 1015 2141 1034
rect 2211 1033 2212 1054
rect 2143 1015 2144 1036
rect 2180 1035 2181 1054
rect 2150 1037 2151 1054
rect 2171 1037 2172 1054
rect 2155 1015 2156 1040
rect 2201 1039 2202 1054
rect 2156 1041 2157 1054
rect 2227 1041 2228 1054
rect 2162 1043 2163 1054
rect 2214 1043 2215 1054
rect 2195 1045 2196 1054
rect 2221 1045 2222 1054
rect 2224 1045 2225 1054
rect 2243 1045 2244 1054
rect 2233 1047 2234 1054
rect 2236 1047 2237 1054
rect 2246 1047 2247 1054
rect 2274 1047 2275 1054
rect 2255 1049 2256 1054
rect 2264 1049 2265 1054
rect 2258 1051 2259 1054
rect 2261 1051 2262 1054
rect 2084 1058 2085 1061
rect 2230 1060 2231 1139
rect 2084 1062 2085 1139
rect 2143 1062 2144 1139
rect 2087 1058 2088 1065
rect 2159 1058 2160 1065
rect 2077 1058 2078 1067
rect 2158 1066 2159 1139
rect 2078 1068 2079 1139
rect 2389 1068 2390 1139
rect 2098 1058 2099 1071
rect 2311 1070 2312 1139
rect 2114 1058 2115 1073
rect 2251 1072 2252 1139
rect 2124 1074 2125 1139
rect 2156 1058 2157 1075
rect 2129 1058 2130 1077
rect 2176 1076 2177 1139
rect 2138 1058 2139 1079
rect 2155 1078 2156 1139
rect 2152 1080 2153 1139
rect 2162 1058 2163 1081
rect 2120 1058 2121 1083
rect 2161 1082 2162 1139
rect 2111 1058 2112 1085
rect 2121 1084 2122 1139
rect 2165 1058 2166 1085
rect 2218 1058 2219 1085
rect 2168 1058 2169 1087
rect 2266 1086 2267 1139
rect 2174 1058 2175 1089
rect 2218 1088 2219 1139
rect 2180 1058 2181 1091
rect 2278 1090 2279 1139
rect 2095 1092 2096 1139
rect 2179 1092 2180 1139
rect 2201 1058 2202 1093
rect 2227 1058 2228 1093
rect 2207 1058 2208 1095
rect 2281 1094 2282 1139
rect 2185 1096 2186 1139
rect 2206 1096 2207 1139
rect 2221 1058 2222 1097
rect 2290 1096 2291 1139
rect 2224 1058 2225 1099
rect 2323 1098 2324 1139
rect 2233 1058 2234 1101
rect 2317 1100 2318 1139
rect 2091 1102 2092 1139
rect 2233 1102 2234 1139
rect 2236 1058 2237 1103
rect 2353 1102 2354 1139
rect 2147 1058 2148 1105
rect 2236 1104 2237 1139
rect 2239 1058 2240 1105
rect 2350 1104 2351 1139
rect 2167 1106 2168 1139
rect 2239 1106 2240 1139
rect 2243 1058 2244 1107
rect 2341 1106 2342 1139
rect 2171 1058 2172 1109
rect 2242 1108 2243 1139
rect 2132 1058 2133 1111
rect 2170 1110 2171 1139
rect 2246 1058 2247 1111
rect 2338 1110 2339 1139
rect 2183 1058 2184 1113
rect 2245 1112 2246 1139
rect 2182 1114 2183 1139
rect 2195 1058 2196 1115
rect 2080 1058 2081 1117
rect 2194 1116 2195 1139
rect 2081 1118 2082 1139
rect 2127 1118 2128 1139
rect 2255 1058 2256 1119
rect 2380 1118 2381 1139
rect 2211 1058 2212 1121
rect 2254 1120 2255 1139
rect 2198 1058 2199 1123
rect 2212 1122 2213 1139
rect 2258 1058 2259 1123
rect 2383 1122 2384 1139
rect 2268 1058 2269 1125
rect 2362 1124 2363 1139
rect 2088 1126 2089 1139
rect 2269 1126 2270 1139
rect 2271 1058 2272 1127
rect 2386 1126 2387 1139
rect 2274 1058 2275 1129
rect 2406 1128 2407 1139
rect 2299 1130 2300 1139
rect 2430 1130 2431 1139
rect 2335 1132 2336 1139
rect 2393 1132 2394 1139
rect 2371 1134 2372 1139
rect 2440 1134 2441 1139
rect 2409 1136 2410 1139
rect 2416 1136 2417 1139
rect 2068 1143 2069 1146
rect 2248 1145 2249 1254
rect 2072 1143 2073 1148
rect 2275 1147 2276 1254
rect 2078 1143 2079 1150
rect 2093 1149 2094 1254
rect 2084 1143 2085 1152
rect 2272 1151 2273 1254
rect 2087 1153 2088 1254
rect 2302 1153 2303 1254
rect 2098 1143 2099 1156
rect 2293 1155 2294 1254
rect 2099 1157 2100 1254
rect 2230 1143 2231 1158
rect 2108 1159 2109 1254
rect 2179 1143 2180 1160
rect 2117 1143 2118 1162
rect 2145 1161 2146 1254
rect 2121 1163 2122 1254
rect 2404 1163 2405 1254
rect 2124 1165 2125 1254
rect 2278 1143 2279 1166
rect 2135 1167 2136 1254
rect 2266 1143 2267 1168
rect 2137 1143 2138 1170
rect 2284 1169 2285 1254
rect 2143 1143 2144 1172
rect 2172 1171 2173 1254
rect 2152 1143 2153 1174
rect 2199 1173 2200 1254
rect 2155 1143 2156 1176
rect 2287 1175 2288 1254
rect 2081 1143 2082 1178
rect 2154 1177 2155 1254
rect 2161 1143 2162 1178
rect 2278 1177 2279 1254
rect 2127 1143 2128 1180
rect 2160 1179 2161 1254
rect 2128 1181 2129 1254
rect 2314 1181 2315 1254
rect 2167 1143 2168 1184
rect 2245 1143 2246 1184
rect 2065 1143 2066 1186
rect 2245 1185 2246 1254
rect 2062 1187 2063 1254
rect 2066 1187 2067 1254
rect 2176 1143 2177 1188
rect 2220 1187 2221 1254
rect 2178 1189 2179 1254
rect 2389 1143 2390 1190
rect 2182 1143 2183 1192
rect 2194 1143 2195 1192
rect 2206 1143 2207 1192
rect 2263 1191 2264 1254
rect 2212 1143 2213 1194
rect 2296 1193 2297 1254
rect 2170 1143 2171 1196
rect 2211 1195 2212 1254
rect 2233 1143 2234 1196
rect 2308 1195 2309 1254
rect 2236 1143 2237 1198
rect 2257 1197 2258 1254
rect 2239 1143 2240 1200
rect 2329 1199 2330 1254
rect 2242 1143 2243 1202
rect 2332 1201 2333 1254
rect 2251 1143 2252 1204
rect 2326 1203 2327 1254
rect 2269 1143 2270 1206
rect 2356 1205 2357 1254
rect 2080 1207 2081 1254
rect 2269 1207 2270 1254
rect 2281 1143 2282 1208
rect 2359 1207 2360 1254
rect 2281 1209 2282 1254
rect 2443 1143 2444 1210
rect 2290 1143 2291 1212
rect 2374 1211 2375 1254
rect 2114 1143 2115 1214
rect 2290 1213 2291 1254
rect 2114 1215 2115 1254
rect 2181 1215 2182 1254
rect 2299 1143 2300 1216
rect 2386 1215 2387 1254
rect 2311 1143 2312 1218
rect 2398 1217 2399 1254
rect 2117 1219 2118 1254
rect 2311 1219 2312 1254
rect 2317 1143 2318 1220
rect 2446 1219 2447 1254
rect 2131 1221 2132 1254
rect 2317 1221 2318 1254
rect 2335 1143 2336 1222
rect 2443 1221 2444 1254
rect 2218 1143 2219 1224
rect 2335 1223 2336 1254
rect 2158 1143 2159 1226
rect 2217 1225 2218 1254
rect 2338 1143 2339 1226
rect 2518 1225 2519 1254
rect 2341 1143 2342 1228
rect 2428 1227 2429 1254
rect 2254 1143 2255 1230
rect 2341 1229 2342 1254
rect 2350 1143 2351 1230
rect 2458 1229 2459 1254
rect 2353 1143 2354 1232
rect 2461 1231 2462 1254
rect 2142 1233 2143 1254
rect 2353 1233 2354 1254
rect 2362 1143 2363 1234
rect 2464 1233 2465 1254
rect 2371 1143 2372 1236
rect 2486 1235 2487 1254
rect 2380 1143 2381 1238
rect 2502 1237 2503 1254
rect 2383 1143 2384 1240
rect 2489 1239 2490 1254
rect 2377 1241 2378 1254
rect 2383 1241 2384 1254
rect 2396 1143 2397 1242
rect 2440 1241 2441 1254
rect 2406 1143 2407 1244
rect 2409 1143 2410 1244
rect 2410 1245 2411 1254
rect 2470 1245 2471 1254
rect 2430 1143 2431 1248
rect 2492 1247 2493 1254
rect 2323 1143 2324 1250
rect 2431 1249 2432 1254
rect 2433 1143 2434 1250
rect 2467 1249 2468 1254
rect 2483 1249 2484 1254
rect 2563 1249 2564 1254
rect 2515 1251 2516 1254
rect 2521 1251 2522 1254
rect 2059 1258 2060 1261
rect 2281 1258 2282 1261
rect 2068 1262 2069 1387
rect 2108 1258 2109 1263
rect 2073 1258 2074 1265
rect 2345 1264 2346 1387
rect 2072 1266 2073 1387
rect 2245 1258 2246 1267
rect 2080 1258 2081 1269
rect 2204 1268 2205 1387
rect 2086 1270 2087 1387
rect 2201 1270 2202 1387
rect 2093 1258 2094 1273
rect 2112 1272 2113 1387
rect 2096 1258 2097 1275
rect 2369 1274 2370 1387
rect 2118 1276 2119 1387
rect 2302 1258 2303 1277
rect 2124 1258 2125 1279
rect 2408 1278 2409 1387
rect 2125 1280 2126 1387
rect 2311 1258 2312 1281
rect 2128 1258 2129 1283
rect 2351 1282 2352 1387
rect 2142 1258 2143 1285
rect 2326 1258 2327 1285
rect 2131 1258 2132 1287
rect 2141 1286 2142 1387
rect 2160 1258 2161 1287
rect 2231 1286 2232 1387
rect 2165 1288 2166 1387
rect 2172 1258 2173 1289
rect 2181 1258 2182 1289
rect 2207 1288 2208 1387
rect 2189 1290 2190 1387
rect 2199 1258 2200 1291
rect 2211 1258 2212 1291
rect 2240 1290 2241 1387
rect 2220 1258 2221 1293
rect 2252 1292 2253 1387
rect 2226 1258 2227 1295
rect 2329 1258 2330 1295
rect 2178 1258 2179 1297
rect 2225 1296 2226 1387
rect 2154 1258 2155 1299
rect 2177 1298 2178 1387
rect 2233 1258 2234 1299
rect 2353 1258 2354 1299
rect 2217 1258 2218 1301
rect 2234 1300 2235 1387
rect 2272 1258 2273 1301
rect 2312 1300 2313 1387
rect 2138 1258 2139 1303
rect 2273 1302 2274 1387
rect 2275 1258 2276 1303
rect 2321 1302 2322 1387
rect 2248 1258 2249 1305
rect 2276 1304 2277 1387
rect 2278 1258 2279 1305
rect 2348 1304 2349 1387
rect 2284 1258 2285 1307
rect 2392 1258 2393 1307
rect 2287 1258 2288 1309
rect 2390 1308 2391 1387
rect 2290 1258 2291 1311
rect 2327 1310 2328 1387
rect 2079 1312 2080 1387
rect 2291 1312 2292 1387
rect 2293 1258 2294 1313
rect 2372 1312 2373 1387
rect 2296 1258 2297 1315
rect 2363 1314 2364 1387
rect 2257 1258 2258 1317
rect 2297 1316 2298 1387
rect 2096 1318 2097 1387
rect 2258 1318 2259 1387
rect 2314 1258 2315 1319
rect 2339 1318 2340 1387
rect 2263 1258 2264 1321
rect 2315 1320 2316 1387
rect 2093 1322 2094 1387
rect 2264 1322 2265 1387
rect 2317 1258 2318 1323
rect 2354 1322 2355 1387
rect 2335 1258 2336 1325
rect 2381 1324 2382 1387
rect 2236 1258 2237 1327
rect 2336 1326 2337 1387
rect 2341 1258 2342 1327
rect 2393 1326 2394 1387
rect 2356 1258 2357 1329
rect 2396 1328 2397 1387
rect 2308 1258 2309 1331
rect 2357 1330 2358 1387
rect 2269 1258 2270 1333
rect 2309 1332 2310 1387
rect 2100 1334 2101 1387
rect 2270 1334 2271 1387
rect 2359 1258 2360 1335
rect 2417 1334 2418 1387
rect 2114 1258 2115 1337
rect 2360 1336 2361 1387
rect 2374 1258 2375 1337
rect 2438 1336 2439 1387
rect 2332 1258 2333 1339
rect 2375 1338 2376 1387
rect 2121 1258 2122 1341
rect 2333 1340 2334 1387
rect 2377 1258 2378 1341
rect 2426 1340 2427 1387
rect 2410 1258 2411 1343
rect 2471 1342 2472 1387
rect 2435 1344 2436 1387
rect 2589 1344 2590 1387
rect 2440 1258 2441 1347
rect 2534 1346 2535 1387
rect 2386 1258 2387 1349
rect 2441 1348 2442 1387
rect 2090 1258 2091 1351
rect 2387 1350 2388 1387
rect 2443 1258 2444 1351
rect 2495 1350 2496 1387
rect 2446 1258 2447 1353
rect 2507 1352 2508 1387
rect 2447 1354 2448 1387
rect 2555 1354 2556 1387
rect 2458 1258 2459 1357
rect 2519 1356 2520 1387
rect 2398 1258 2399 1359
rect 2459 1358 2460 1387
rect 2145 1258 2146 1361
rect 2399 1360 2400 1387
rect 2461 1258 2462 1361
rect 2522 1360 2523 1387
rect 2464 1258 2465 1363
rect 2525 1362 2526 1387
rect 2404 1258 2405 1365
rect 2465 1364 2466 1387
rect 2229 1258 2230 1367
rect 2405 1366 2406 1387
rect 2467 1258 2468 1367
rect 2528 1366 2529 1387
rect 2483 1258 2484 1369
rect 2543 1368 2544 1387
rect 2486 1258 2487 1371
rect 2546 1370 2547 1387
rect 2489 1258 2490 1373
rect 2576 1372 2577 1387
rect 2428 1258 2429 1375
rect 2489 1374 2490 1387
rect 2492 1258 2493 1375
rect 2564 1374 2565 1387
rect 2431 1258 2432 1377
rect 2492 1376 2493 1387
rect 2365 1258 2366 1379
rect 2432 1378 2433 1387
rect 2502 1258 2503 1379
rect 2549 1378 2550 1387
rect 2515 1258 2516 1381
rect 2607 1380 2608 1387
rect 2531 1382 2532 1387
rect 2586 1382 2587 1387
rect 2567 1384 2568 1387
rect 2621 1384 2622 1387
rect 2645 1384 2646 1387
rect 2648 1384 2649 1387
rect 2065 1391 2066 1394
rect 2324 1393 2325 1574
rect 2072 1395 2073 1574
rect 2342 1395 2343 1574
rect 2082 1391 2083 1398
rect 2318 1397 2319 1574
rect 2086 1399 2087 1574
rect 2201 1391 2202 1400
rect 2093 1401 2094 1574
rect 2327 1391 2328 1402
rect 2096 1391 2097 1404
rect 2252 1391 2253 1404
rect 2096 1405 2097 1574
rect 2240 1391 2241 1406
rect 2105 1407 2106 1574
rect 2112 1391 2113 1408
rect 2108 1409 2109 1574
rect 2147 1409 2148 1574
rect 2111 1411 2112 1574
rect 2201 1411 2202 1574
rect 2115 1391 2116 1414
rect 2252 1413 2253 1574
rect 2115 1415 2116 1574
rect 2402 1415 2403 1574
rect 2118 1391 2119 1418
rect 2504 1417 2505 1574
rect 2118 1419 2119 1574
rect 2384 1419 2385 1574
rect 2122 1421 2123 1574
rect 2366 1421 2367 1574
rect 2132 1391 2133 1424
rect 2336 1391 2337 1424
rect 2134 1425 2135 1574
rect 2141 1391 2142 1426
rect 2140 1427 2141 1574
rect 2189 1391 2190 1428
rect 2143 1429 2144 1574
rect 2390 1391 2391 1430
rect 2159 1431 2160 1574
rect 2165 1391 2166 1432
rect 2177 1391 2178 1432
rect 2189 1431 2190 1574
rect 2177 1433 2178 1574
rect 2474 1433 2475 1574
rect 2195 1435 2196 1574
rect 2207 1391 2208 1436
rect 2204 1391 2205 1438
rect 2222 1437 2223 1574
rect 2219 1391 2220 1440
rect 2399 1391 2400 1440
rect 2089 1441 2090 1574
rect 2219 1441 2220 1574
rect 2225 1391 2226 1442
rect 2243 1441 2244 1574
rect 2225 1443 2226 1574
rect 2408 1391 2409 1444
rect 2228 1391 2229 1446
rect 2393 1391 2394 1446
rect 2231 1391 2232 1448
rect 2246 1447 2247 1574
rect 2234 1391 2235 1450
rect 2237 1449 2238 1574
rect 2258 1391 2259 1450
rect 2282 1449 2283 1574
rect 2068 1391 2069 1452
rect 2258 1451 2259 1574
rect 2068 1453 2069 1574
rect 2291 1391 2292 1454
rect 2264 1391 2265 1456
rect 2288 1455 2289 1574
rect 2264 1457 2265 1574
rect 2270 1391 2271 1458
rect 2276 1391 2277 1458
rect 2327 1457 2328 1574
rect 2279 1459 2280 1574
rect 2393 1459 2394 1574
rect 2297 1391 2298 1462
rect 2330 1461 2331 1574
rect 2321 1391 2322 1464
rect 2336 1463 2337 1574
rect 2333 1391 2334 1466
rect 2390 1465 2391 1574
rect 2339 1391 2340 1468
rect 2408 1467 2409 1574
rect 2354 1391 2355 1470
rect 2411 1469 2412 1574
rect 2345 1391 2346 1472
rect 2354 1471 2355 1574
rect 2369 1391 2370 1472
rect 2378 1471 2379 1574
rect 2375 1391 2376 1474
rect 2444 1473 2445 1574
rect 2405 1391 2406 1476
rect 2456 1475 2457 1574
rect 2273 1391 2274 1478
rect 2405 1477 2406 1574
rect 2414 1391 2415 1478
rect 2498 1477 2499 1574
rect 2363 1391 2364 1480
rect 2414 1479 2415 1574
rect 2417 1391 2418 1480
rect 2486 1479 2487 1574
rect 2426 1391 2427 1482
rect 2450 1481 2451 1574
rect 2156 1391 2157 1484
rect 2426 1483 2427 1574
rect 2435 1391 2436 1484
rect 2585 1483 2586 1574
rect 2396 1391 2397 1486
rect 2435 1485 2436 1574
rect 2351 1391 2352 1488
rect 2396 1487 2397 1574
rect 2312 1391 2313 1490
rect 2351 1489 2352 1574
rect 2312 1491 2313 1574
rect 2432 1391 2433 1492
rect 2381 1391 2382 1494
rect 2432 1493 2433 1574
rect 2372 1391 2373 1496
rect 2381 1495 2382 1574
rect 2357 1391 2358 1498
rect 2372 1497 2373 1574
rect 2348 1391 2349 1500
rect 2357 1499 2358 1574
rect 2309 1391 2310 1502
rect 2348 1501 2349 1574
rect 2438 1391 2439 1502
rect 2667 1501 2668 1574
rect 2125 1391 2126 1504
rect 2438 1503 2439 1574
rect 2441 1391 2442 1504
rect 2468 1503 2469 1574
rect 2387 1391 2388 1506
rect 2441 1505 2442 1574
rect 2360 1391 2361 1508
rect 2387 1507 2388 1574
rect 2315 1391 2316 1510
rect 2360 1509 2361 1574
rect 2447 1391 2448 1510
rect 2462 1509 2463 1574
rect 2453 1391 2454 1512
rect 2582 1511 2583 1574
rect 2459 1391 2460 1514
rect 2516 1513 2517 1574
rect 2459 1515 2460 1574
rect 2552 1391 2553 1516
rect 2471 1391 2472 1518
rect 2594 1517 2595 1574
rect 2501 1519 2502 1574
rect 2573 1391 2574 1520
rect 2507 1391 2508 1522
rect 2600 1521 2601 1574
rect 2510 1523 2511 1574
rect 2728 1523 2729 1574
rect 2519 1391 2520 1526
rect 2636 1525 2637 1574
rect 2522 1391 2523 1528
rect 2639 1527 2640 1574
rect 2522 1529 2523 1574
rect 2725 1529 2726 1574
rect 2525 1391 2526 1532
rect 2606 1531 2607 1574
rect 2528 1391 2529 1534
rect 2609 1533 2610 1574
rect 2465 1391 2466 1536
rect 2528 1535 2529 1574
rect 2531 1391 2532 1536
rect 2654 1535 2655 1574
rect 2534 1391 2535 1538
rect 2657 1537 2658 1574
rect 2537 1391 2538 1540
rect 2660 1539 2661 1574
rect 2540 1541 2541 1574
rect 2591 1541 2592 1574
rect 2543 1391 2544 1544
rect 2612 1543 2613 1574
rect 2276 1545 2277 1574
rect 2543 1545 2544 1574
rect 2546 1391 2547 1546
rect 2627 1545 2628 1574
rect 2546 1547 2547 1574
rect 2663 1547 2664 1574
rect 2549 1391 2550 1550
rect 2633 1549 2634 1574
rect 2564 1391 2565 1552
rect 2624 1391 2625 1552
rect 2495 1391 2496 1554
rect 2564 1553 2565 1574
rect 2306 1391 2307 1556
rect 2495 1555 2496 1574
rect 2306 1557 2307 1574
rect 2690 1557 2691 1574
rect 2567 1391 2568 1560
rect 2651 1559 2652 1574
rect 2576 1391 2577 1562
rect 2674 1561 2675 1574
rect 2489 1391 2490 1564
rect 2576 1563 2577 1574
rect 2579 1391 2580 1564
rect 2680 1563 2681 1574
rect 2492 1391 2493 1566
rect 2579 1565 2580 1574
rect 2261 1567 2262 1574
rect 2492 1567 2493 1574
rect 2630 1567 2631 1574
rect 2735 1567 2736 1574
rect 2648 1391 2649 1570
rect 2745 1569 2746 1574
rect 2621 1391 2622 1572
rect 2648 1571 2649 1574
rect 2057 1580 2058 1761
rect 2122 1580 2123 1761
rect 2072 1578 2073 1583
rect 2094 1582 2095 1761
rect 2075 1578 2076 1585
rect 2096 1578 2097 1585
rect 2075 1586 2076 1761
rect 2306 1578 2307 1587
rect 2089 1578 2090 1589
rect 2222 1578 2223 1589
rect 2101 1590 2102 1761
rect 2219 1578 2220 1591
rect 2105 1578 2106 1593
rect 2131 1592 2132 1761
rect 2111 1578 2112 1595
rect 2195 1578 2196 1595
rect 2116 1596 2117 1761
rect 2327 1578 2328 1597
rect 2119 1598 2120 1761
rect 2360 1578 2361 1599
rect 2128 1600 2129 1761
rect 2159 1578 2160 1601
rect 2134 1578 2135 1603
rect 2153 1602 2154 1761
rect 2134 1604 2135 1761
rect 2303 1604 2304 1761
rect 2140 1578 2141 1607
rect 2183 1606 2184 1761
rect 2143 1578 2144 1609
rect 2465 1608 2466 1761
rect 2171 1610 2172 1761
rect 2564 1578 2565 1611
rect 2189 1578 2190 1613
rect 2219 1612 2220 1761
rect 2201 1578 2202 1615
rect 2234 1614 2235 1761
rect 2225 1578 2226 1617
rect 2240 1616 2241 1761
rect 2231 1618 2232 1761
rect 2683 1578 2684 1619
rect 2237 1578 2238 1621
rect 2267 1620 2268 1761
rect 2258 1578 2259 1623
rect 2414 1578 2415 1623
rect 2243 1578 2244 1625
rect 2258 1624 2259 1761
rect 2261 1578 2262 1625
rect 2480 1624 2481 1761
rect 2252 1578 2253 1627
rect 2261 1626 2262 1761
rect 2246 1578 2247 1629
rect 2252 1628 2253 1761
rect 2264 1578 2265 1629
rect 2273 1628 2274 1761
rect 2276 1578 2277 1629
rect 2639 1578 2640 1629
rect 2282 1578 2283 1631
rect 2291 1630 2292 1761
rect 2285 1632 2286 1761
rect 2357 1578 2358 1633
rect 2288 1578 2289 1635
rect 2297 1634 2298 1761
rect 2315 1634 2316 1761
rect 2704 1578 2705 1635
rect 2318 1578 2319 1637
rect 2321 1636 2322 1761
rect 2324 1578 2325 1637
rect 2327 1636 2328 1761
rect 2330 1636 2331 1761
rect 2330 1578 2331 1637
rect 2336 1636 2337 1761
rect 2336 1578 2337 1637
rect 2342 1636 2343 1761
rect 2342 1578 2343 1637
rect 2351 1578 2352 1637
rect 2369 1636 2370 1761
rect 2098 1638 2099 1761
rect 2351 1638 2352 1761
rect 2363 1638 2364 1761
rect 2504 1578 2505 1639
rect 2378 1638 2379 1761
rect 2378 1578 2379 1639
rect 2381 1638 2382 1761
rect 2381 1578 2382 1639
rect 2396 1578 2397 1641
rect 2414 1640 2415 1761
rect 2396 1642 2397 1761
rect 2402 1578 2403 1643
rect 2390 1578 2391 1645
rect 2402 1644 2403 1761
rect 2384 1578 2385 1647
rect 2390 1646 2391 1761
rect 2372 1578 2373 1649
rect 2384 1648 2385 1761
rect 2366 1578 2367 1651
rect 2372 1650 2373 1761
rect 2082 1578 2083 1653
rect 2366 1652 2367 1761
rect 2068 1578 2069 1655
rect 2081 1654 2082 1761
rect 2068 1656 2069 1761
rect 2165 1656 2166 1761
rect 2399 1656 2400 1761
rect 2405 1578 2406 1657
rect 2393 1578 2394 1659
rect 2405 1658 2406 1761
rect 2387 1578 2388 1661
rect 2393 1660 2394 1761
rect 2408 1578 2409 1661
rect 2420 1660 2421 1761
rect 2408 1662 2409 1761
rect 2426 1578 2427 1663
rect 2411 1578 2412 1665
rect 2423 1664 2424 1761
rect 2432 1578 2433 1665
rect 2552 1664 2553 1761
rect 2432 1666 2433 1761
rect 2441 1578 2442 1667
rect 2435 1578 2436 1669
rect 2555 1668 2556 1761
rect 2450 1668 2451 1761
rect 2450 1578 2451 1669
rect 2459 1578 2460 1671
rect 2489 1670 2490 1761
rect 2462 1578 2463 1673
rect 2726 1672 2727 1761
rect 2438 1578 2439 1675
rect 2462 1674 2463 1761
rect 2438 1676 2439 1761
rect 2670 1578 2671 1677
rect 2468 1578 2469 1679
rect 2667 1578 2668 1679
rect 2456 1578 2457 1681
rect 2468 1680 2469 1761
rect 2456 1682 2457 1761
rect 2669 1682 2670 1761
rect 2474 1578 2475 1685
rect 2588 1684 2589 1761
rect 2150 1578 2151 1687
rect 2474 1686 2475 1761
rect 2486 1578 2487 1687
rect 2531 1686 2532 1761
rect 2444 1578 2445 1689
rect 2486 1688 2487 1761
rect 2162 1690 2163 1761
rect 2444 1690 2445 1761
rect 2492 1578 2493 1691
rect 2558 1690 2559 1761
rect 2495 1578 2496 1693
rect 2561 1692 2562 1761
rect 2504 1694 2505 1761
rect 2510 1578 2511 1695
rect 2501 1578 2502 1697
rect 2510 1696 2511 1761
rect 2516 1578 2517 1697
rect 2525 1696 2526 1761
rect 2498 1578 2499 1699
rect 2516 1698 2517 1761
rect 2519 1698 2520 1761
rect 2784 1698 2785 1761
rect 2522 1578 2523 1701
rect 2537 1700 2538 1761
rect 2543 1578 2544 1701
rect 2570 1700 2571 1761
rect 2543 1702 2544 1761
rect 2609 1578 2610 1703
rect 2546 1578 2547 1705
rect 2591 1578 2592 1705
rect 2528 1578 2529 1707
rect 2546 1706 2547 1761
rect 2564 1706 2565 1761
rect 2791 1706 2792 1761
rect 2582 1578 2583 1709
rect 2666 1708 2667 1761
rect 2582 1710 2583 1761
rect 2674 1578 2675 1711
rect 2585 1578 2586 1713
rect 2663 1712 2664 1761
rect 2594 1578 2595 1715
rect 2684 1714 2685 1761
rect 2540 1578 2541 1717
rect 2594 1716 2595 1761
rect 2600 1578 2601 1717
rect 2711 1716 2712 1761
rect 2579 1578 2580 1719
rect 2600 1718 2601 1761
rect 2606 1578 2607 1719
rect 2697 1578 2698 1719
rect 2624 1720 2625 1761
rect 2794 1720 2795 1761
rect 2627 1578 2628 1723
rect 2675 1722 2676 1761
rect 2576 1578 2577 1725
rect 2627 1724 2628 1761
rect 2360 1726 2361 1761
rect 2576 1726 2577 1761
rect 2630 1578 2631 1727
rect 2787 1726 2788 1761
rect 2633 1578 2634 1729
rect 2678 1728 2679 1761
rect 2636 1578 2637 1731
rect 2708 1730 2709 1761
rect 2636 1732 2637 1761
rect 2766 1732 2767 1761
rect 2639 1734 2640 1761
rect 2763 1734 2764 1761
rect 2642 1736 2643 1761
rect 2756 1736 2757 1761
rect 2648 1578 2649 1739
rect 2696 1738 2697 1761
rect 2651 1578 2652 1741
rect 2699 1740 2700 1761
rect 2654 1578 2655 1743
rect 2720 1742 2721 1761
rect 2612 1578 2613 1745
rect 2654 1744 2655 1761
rect 2657 1578 2658 1745
rect 2723 1744 2724 1761
rect 2312 1578 2313 1747
rect 2657 1746 2658 1761
rect 2159 1748 2160 1761
rect 2312 1748 2313 1761
rect 2660 1578 2661 1749
rect 2714 1748 2715 1761
rect 2279 1578 2280 1751
rect 2660 1750 2661 1761
rect 2137 1752 2138 1761
rect 2279 1752 2280 1761
rect 2680 1578 2681 1753
rect 2739 1752 2740 1761
rect 2681 1754 2682 1761
rect 2718 1578 2719 1755
rect 2513 1756 2514 1761
rect 2717 1756 2718 1761
rect 2745 1578 2746 1757
rect 2818 1756 2819 1761
rect 2808 1758 2809 1761
rect 2812 1758 2813 1761
rect 2047 1765 2048 1768
rect 2122 1765 2123 1768
rect 2054 1765 2055 1770
rect 2075 1765 2076 1770
rect 2059 1771 2060 2014
rect 2075 1771 2076 2014
rect 2061 1765 2062 1774
rect 2081 1765 2082 1774
rect 2071 1765 2072 1776
rect 2454 1775 2455 2014
rect 2064 1765 2065 1778
rect 2072 1777 2073 2014
rect 2078 1777 2079 2014
rect 2165 1765 2166 1778
rect 2087 1765 2088 1780
rect 2348 1765 2349 1780
rect 2089 1781 2090 2014
rect 2234 1765 2235 1782
rect 2082 1783 2083 2014
rect 2235 1783 2236 2014
rect 2092 1785 2093 2014
rect 2376 1785 2377 2014
rect 2113 1787 2114 2014
rect 2354 1765 2355 1788
rect 2116 1765 2117 1790
rect 2384 1765 2385 1790
rect 2119 1765 2120 1792
rect 2390 1765 2391 1792
rect 2119 1793 2120 2014
rect 2131 1765 2132 1794
rect 2125 1765 2126 1796
rect 2423 1765 2424 1796
rect 2128 1765 2129 1798
rect 2460 1797 2461 2014
rect 2129 1799 2130 2014
rect 2153 1765 2154 1800
rect 2134 1765 2135 1802
rect 2256 1801 2257 2014
rect 2137 1765 2138 1804
rect 2273 1765 2274 1804
rect 2144 1765 2145 1806
rect 2444 1765 2445 1806
rect 2125 1807 2126 2014
rect 2144 1807 2145 2014
rect 2148 1807 2149 2014
rect 2499 1807 2500 2014
rect 2171 1765 2172 1810
rect 2378 1765 2379 1810
rect 2174 1765 2175 1812
rect 2279 1765 2280 1812
rect 2181 1813 2182 2014
rect 2489 1765 2490 1814
rect 2202 1815 2203 2014
rect 2231 1765 2232 1816
rect 2205 1817 2206 2014
rect 2219 1765 2220 1818
rect 2207 1765 2208 1820
rect 2486 1765 2487 1820
rect 2210 1765 2211 1822
rect 2673 1821 2674 2014
rect 2223 1823 2224 2014
rect 2252 1765 2253 1824
rect 2229 1825 2230 2014
rect 2393 1765 2394 1826
rect 2240 1765 2241 1828
rect 2472 1827 2473 2014
rect 2241 1829 2242 2014
rect 2258 1765 2259 1830
rect 2244 1831 2245 2014
rect 2309 1765 2310 1832
rect 2250 1833 2251 2014
rect 2267 1765 2268 1834
rect 2268 1835 2269 2014
rect 2291 1765 2292 1836
rect 2274 1837 2275 2014
rect 2297 1765 2298 1838
rect 2280 1839 2281 2014
rect 2303 1765 2304 1840
rect 2289 1841 2290 2014
rect 2627 1765 2628 1842
rect 2292 1843 2293 2014
rect 2315 1765 2316 1844
rect 2310 1845 2311 2014
rect 2321 1765 2322 1846
rect 2312 1765 2313 1848
rect 2715 1847 2716 2014
rect 2316 1849 2317 2014
rect 2330 1765 2331 1850
rect 2322 1851 2323 2014
rect 2372 1765 2373 1852
rect 2327 1765 2328 1854
rect 2391 1853 2392 2014
rect 2328 1855 2329 2014
rect 2402 1765 2403 1856
rect 2151 1857 2152 2014
rect 2403 1857 2404 2014
rect 2331 1859 2332 2014
rect 2405 1765 2406 1860
rect 2334 1861 2335 2014
rect 2570 1765 2571 1862
rect 2346 1863 2347 2014
rect 2438 1765 2439 1864
rect 2351 1765 2352 1866
rect 2436 1865 2437 2014
rect 2352 1867 2353 2014
rect 2552 1765 2553 1868
rect 2355 1869 2356 2014
rect 2555 1765 2556 1870
rect 2360 1765 2361 1872
rect 2588 1765 2589 1872
rect 2363 1765 2364 1874
rect 2594 1765 2595 1874
rect 2364 1875 2365 2014
rect 2561 1765 2562 1876
rect 2379 1877 2380 2014
rect 2657 1765 2658 1878
rect 2385 1879 2386 2014
rect 2462 1765 2463 1880
rect 2366 1765 2367 1882
rect 2463 1881 2464 2014
rect 2396 1765 2397 1884
rect 2487 1883 2488 2014
rect 2101 1885 2102 2014
rect 2397 1885 2398 2014
rect 2399 1765 2400 1886
rect 2490 1885 2491 2014
rect 2381 1765 2382 1888
rect 2400 1887 2401 2014
rect 2420 1765 2421 1888
rect 2445 1887 2446 2014
rect 2068 1765 2069 1890
rect 2421 1889 2422 2014
rect 2069 1891 2070 2014
rect 2319 1891 2320 2014
rect 2427 1891 2428 2014
rect 2808 1765 2809 1892
rect 2432 1765 2433 1894
rect 2493 1893 2494 2014
rect 2342 1765 2343 1896
rect 2433 1895 2434 2014
rect 2439 1895 2440 2014
rect 2468 1765 2469 1896
rect 2098 1765 2099 1898
rect 2469 1897 2470 2014
rect 2465 1765 2466 1900
rect 2508 1899 2509 2014
rect 2369 1765 2370 1902
rect 2466 1901 2467 2014
rect 2370 1903 2371 2014
rect 2531 1765 2532 1904
rect 2474 1765 2475 1906
rect 2733 1765 2734 1906
rect 2475 1907 2476 2014
rect 2564 1765 2565 1908
rect 2480 1765 2481 1910
rect 2481 1909 2482 2014
rect 2484 1909 2485 2014
rect 2558 1765 2559 1910
rect 2504 1765 2505 1912
rect 2589 1911 2590 2014
rect 2408 1765 2409 1914
rect 2505 1913 2506 2014
rect 2159 1765 2160 1916
rect 2409 1915 2410 2014
rect 2160 1917 2161 2014
rect 2183 1765 2184 1918
rect 2510 1765 2511 1918
rect 2586 1917 2587 2014
rect 2511 1919 2512 2014
rect 2729 1765 2730 1920
rect 2516 1765 2517 1922
rect 2541 1921 2542 2014
rect 2141 1765 2142 1924
rect 2517 1923 2518 2014
rect 2141 1925 2142 2014
rect 2298 1925 2299 2014
rect 2523 1925 2524 2014
rect 2546 1765 2547 1926
rect 2525 1765 2526 1928
rect 2553 1927 2554 2014
rect 2529 1929 2530 2014
rect 2537 1765 2538 1930
rect 2547 1929 2548 2014
rect 2642 1765 2643 1930
rect 2550 1931 2551 2014
rect 2660 1765 2661 1932
rect 2559 1933 2560 2014
rect 2582 1765 2583 1934
rect 2571 1935 2572 2014
rect 2749 1765 2750 1936
rect 2580 1937 2581 2014
rect 2775 1937 2776 2014
rect 2613 1939 2614 2014
rect 2663 1765 2664 1940
rect 2616 1941 2617 2014
rect 2666 1765 2667 1942
rect 2619 1943 2620 2014
rect 2850 1943 2851 2014
rect 2624 1765 2625 1946
rect 2634 1945 2635 2014
rect 2628 1947 2629 2014
rect 2723 1765 2724 1948
rect 2636 1765 2637 1950
rect 2661 1949 2662 2014
rect 2600 1765 2601 1952
rect 2637 1951 2638 2014
rect 2519 1765 2520 1954
rect 2601 1953 2602 2014
rect 2639 1765 2640 1954
rect 2649 1953 2650 2014
rect 2640 1955 2641 2014
rect 2839 1955 2840 2014
rect 2667 1957 2668 2014
rect 2763 1765 2764 1958
rect 2576 1765 2577 1960
rect 2763 1959 2764 2014
rect 2543 1765 2544 1962
rect 2577 1961 2578 2014
rect 2513 1765 2514 1964
rect 2544 1963 2545 2014
rect 2675 1765 2676 1964
rect 2703 1963 2704 2014
rect 2678 1765 2679 1966
rect 2724 1965 2725 2014
rect 2654 1765 2655 1968
rect 2679 1967 2680 2014
rect 2681 1765 2682 1968
rect 2752 1765 2753 1968
rect 2682 1969 2683 2014
rect 2843 1969 2844 2014
rect 2684 1765 2685 1972
rect 2685 1971 2686 2014
rect 2696 1765 2697 1972
rect 2760 1971 2761 2014
rect 2697 1973 2698 2014
rect 2708 1765 2709 1974
rect 2699 1765 2700 1976
rect 2727 1975 2728 2014
rect 2700 1977 2701 2014
rect 2711 1765 2712 1978
rect 2706 1979 2707 2014
rect 2791 1765 2792 1980
rect 2720 1765 2721 1982
rect 2784 1981 2785 2014
rect 2736 1765 2737 1984
rect 2742 1765 2743 1984
rect 2739 1765 2740 1986
rect 2769 1985 2770 2014
rect 2739 1987 2740 2014
rect 2801 1987 2802 2014
rect 2742 1989 2743 2014
rect 2766 1765 2767 1990
rect 2450 1765 2451 1992
rect 2766 1991 2767 2014
rect 2084 1765 2085 1994
rect 2451 1993 2452 2014
rect 2085 1995 2086 2014
rect 2261 1765 2262 1996
rect 2262 1997 2263 2014
rect 2285 1765 2286 1998
rect 2286 1999 2287 2014
rect 2456 1765 2457 2000
rect 2414 1765 2415 2002
rect 2457 2001 2458 2014
rect 2336 1765 2337 2004
rect 2415 2003 2416 2014
rect 2757 2003 2758 2014
rect 2829 2003 2830 2014
rect 2772 2005 2773 2014
rect 2778 2005 2779 2014
rect 2781 2005 2782 2014
rect 2790 2005 2791 2014
rect 2797 2005 2798 2014
rect 2808 2005 2809 2014
rect 2812 1765 2813 2006
rect 2821 1765 2822 2006
rect 2811 2007 2812 2014
rect 2825 2007 2826 2014
rect 2818 1765 2819 2010
rect 2856 2009 2857 2014
rect 2721 2011 2722 2014
rect 2818 2011 2819 2014
rect 2822 2011 2823 2014
rect 2846 2011 2847 2014
rect 2011 2020 2012 2251
rect 2447 2020 2448 2251
rect 2066 2018 2067 2023
rect 2463 2018 2464 2023
rect 2069 2018 2070 2025
rect 2451 2018 2452 2025
rect 2072 2018 2073 2027
rect 2381 2026 2382 2251
rect 2078 2018 2079 2029
rect 2171 2028 2172 2251
rect 2092 2018 2093 2031
rect 2122 2018 2123 2031
rect 2104 2018 2105 2033
rect 2160 2018 2161 2033
rect 2110 2034 2111 2251
rect 2436 2018 2437 2035
rect 2113 2018 2114 2037
rect 2409 2018 2410 2037
rect 2119 2018 2120 2039
rect 2135 2038 2136 2251
rect 2129 2018 2130 2041
rect 2490 2018 2491 2041
rect 2141 2018 2142 2043
rect 2501 2042 2502 2251
rect 2141 2044 2142 2251
rect 2415 2018 2416 2045
rect 2144 2018 2145 2047
rect 2439 2018 2440 2047
rect 2148 2018 2149 2049
rect 2385 2018 2386 2049
rect 2148 2050 2149 2251
rect 2229 2018 2230 2051
rect 2152 2052 2153 2251
rect 2310 2018 2311 2053
rect 2155 2054 2156 2251
rect 2493 2018 2494 2055
rect 2159 2056 2160 2251
rect 2489 2056 2490 2251
rect 2178 2018 2179 2059
rect 2207 2058 2208 2251
rect 2075 2018 2076 2061
rect 2177 2060 2178 2251
rect 2181 2018 2182 2061
rect 2492 2060 2493 2251
rect 2190 2018 2191 2063
rect 2715 2018 2716 2063
rect 2202 2018 2203 2065
rect 2450 2064 2451 2251
rect 2205 2018 2206 2067
rect 2231 2066 2232 2251
rect 2222 2068 2223 2251
rect 2223 2018 2224 2069
rect 2243 2068 2244 2251
rect 2472 2018 2473 2069
rect 2256 2018 2257 2071
rect 2324 2070 2325 2251
rect 2219 2072 2220 2251
rect 2255 2072 2256 2251
rect 2262 2018 2263 2073
rect 2306 2072 2307 2251
rect 2264 2074 2265 2251
rect 2603 2074 2604 2251
rect 2268 2018 2269 2077
rect 2312 2076 2313 2251
rect 2082 2018 2083 2079
rect 2267 2078 2268 2251
rect 2276 2078 2277 2251
rect 2466 2018 2467 2079
rect 2280 2018 2281 2081
rect 2849 2080 2850 2251
rect 2250 2018 2251 2083
rect 2279 2082 2280 2251
rect 2289 2018 2290 2083
rect 2697 2018 2698 2083
rect 2292 2018 2293 2085
rect 2342 2084 2343 2251
rect 2241 2018 2242 2087
rect 2291 2086 2292 2251
rect 2298 2018 2299 2087
rect 2348 2086 2349 2251
rect 2316 2018 2317 2089
rect 2360 2088 2361 2251
rect 2322 2018 2323 2091
rect 2366 2090 2367 2251
rect 2328 2018 2329 2093
rect 2372 2092 2373 2251
rect 2346 2018 2347 2095
rect 2384 2094 2385 2251
rect 2352 2018 2353 2097
rect 2408 2096 2409 2251
rect 2364 2018 2365 2099
rect 2414 2098 2415 2251
rect 2319 2018 2320 2101
rect 2363 2100 2364 2251
rect 2274 2018 2275 2103
rect 2318 2102 2319 2251
rect 2235 2018 2236 2105
rect 2273 2104 2274 2251
rect 2370 2018 2371 2105
rect 2429 2104 2430 2251
rect 2397 2018 2398 2107
rect 2465 2106 2466 2251
rect 2379 2018 2380 2109
rect 2396 2108 2397 2251
rect 2059 2110 2060 2251
rect 2378 2110 2379 2251
rect 2427 2018 2428 2111
rect 2471 2110 2472 2251
rect 2376 2018 2377 2113
rect 2426 2112 2427 2251
rect 2331 2018 2332 2115
rect 2375 2114 2376 2251
rect 2125 2018 2126 2117
rect 2330 2116 2331 2251
rect 2125 2118 2126 2251
rect 2195 2118 2196 2251
rect 2433 2018 2434 2119
rect 2495 2118 2496 2251
rect 2445 2018 2446 2121
rect 2519 2120 2520 2251
rect 2444 2122 2445 2251
rect 2484 2018 2485 2123
rect 2421 2018 2422 2125
rect 2483 2124 2484 2251
rect 2193 2018 2194 2127
rect 2420 2126 2421 2251
rect 2457 2018 2458 2127
rect 2525 2126 2526 2251
rect 2469 2018 2470 2129
rect 2477 2128 2478 2251
rect 2475 2018 2476 2131
rect 2513 2130 2514 2251
rect 2481 2018 2482 2133
rect 2531 2132 2532 2251
rect 2499 2018 2500 2135
rect 2537 2134 2538 2251
rect 2076 2136 2077 2251
rect 2498 2136 2499 2251
rect 2505 2018 2506 2137
rect 2561 2136 2562 2251
rect 2400 2018 2401 2139
rect 2504 2138 2505 2251
rect 2508 2018 2509 2139
rect 2564 2138 2565 2251
rect 2116 2018 2117 2141
rect 2507 2140 2508 2251
rect 2511 2018 2512 2141
rect 2789 2140 2790 2251
rect 2355 2018 2356 2143
rect 2510 2142 2511 2251
rect 2334 2018 2335 2145
rect 2354 2144 2355 2251
rect 2517 2018 2518 2145
rect 2852 2144 2853 2251
rect 2523 2018 2524 2147
rect 2573 2146 2574 2251
rect 2541 2018 2542 2149
rect 2597 2148 2598 2251
rect 2544 2018 2545 2151
rect 2801 2150 2802 2251
rect 2487 2018 2488 2153
rect 2543 2152 2544 2251
rect 2069 2154 2070 2251
rect 2486 2154 2487 2251
rect 2547 2018 2548 2155
rect 2567 2154 2568 2251
rect 2286 2018 2287 2157
rect 2546 2156 2547 2251
rect 2555 2156 2556 2251
rect 2559 2018 2560 2157
rect 2586 2018 2587 2157
rect 2642 2156 2643 2251
rect 2261 2158 2262 2251
rect 2585 2158 2586 2251
rect 2609 2158 2610 2251
rect 2775 2018 2776 2159
rect 2619 2018 2620 2161
rect 2832 2018 2833 2161
rect 2621 2162 2622 2251
rect 2772 2018 2773 2163
rect 2640 2018 2641 2165
rect 2708 2164 2709 2251
rect 2577 2018 2578 2167
rect 2639 2166 2640 2251
rect 2649 2018 2650 2167
rect 2750 2166 2751 2251
rect 2589 2018 2590 2169
rect 2648 2168 2649 2251
rect 2247 2018 2248 2171
rect 2588 2170 2589 2251
rect 2667 2018 2668 2171
rect 2762 2170 2763 2251
rect 2637 2018 2638 2173
rect 2666 2172 2667 2251
rect 2673 2018 2674 2173
rect 2865 2172 2866 2251
rect 2672 2174 2673 2251
rect 2942 2174 2943 2251
rect 2676 2018 2677 2177
rect 2706 2018 2707 2177
rect 2682 2018 2683 2179
rect 2771 2178 2772 2251
rect 2685 2018 2686 2181
rect 2859 2180 2860 2251
rect 2628 2018 2629 2183
rect 2684 2182 2685 2251
rect 2571 2018 2572 2185
rect 2627 2184 2628 2251
rect 2550 2018 2551 2187
rect 2570 2186 2571 2251
rect 2690 2186 2691 2251
rect 2907 2186 2908 2251
rect 2693 2188 2694 2251
rect 2889 2188 2890 2251
rect 2696 2190 2697 2251
rect 2900 2190 2901 2251
rect 2703 2018 2704 2193
rect 2804 2192 2805 2251
rect 2711 2194 2712 2251
rect 2754 2018 2755 2195
rect 2718 2018 2719 2197
rect 2798 2196 2799 2251
rect 2721 2018 2722 2199
rect 2819 2198 2820 2251
rect 2724 2018 2725 2201
rect 2822 2200 2823 2251
rect 2729 2202 2730 2251
rect 2935 2202 2936 2251
rect 2739 2018 2740 2205
rect 2837 2204 2838 2251
rect 2616 2018 2617 2207
rect 2738 2206 2739 2251
rect 2553 2018 2554 2209
rect 2615 2208 2616 2251
rect 2742 2018 2743 2209
rect 2840 2208 2841 2251
rect 2747 2210 2748 2251
rect 2954 2210 2955 2251
rect 2757 2018 2758 2213
rect 2825 2018 2826 2213
rect 2661 2018 2662 2215
rect 2756 2214 2757 2251
rect 2601 2018 2602 2217
rect 2660 2216 2661 2251
rect 2727 2018 2728 2217
rect 2825 2216 2826 2251
rect 2760 2018 2761 2219
rect 2877 2218 2878 2251
rect 2766 2018 2767 2221
rect 2896 2220 2897 2251
rect 2769 2018 2770 2223
rect 2862 2222 2863 2251
rect 2679 2018 2680 2225
rect 2768 2224 2769 2251
rect 2781 2018 2782 2225
rect 2880 2224 2881 2251
rect 2613 2018 2614 2227
rect 2780 2226 2781 2251
rect 2784 2018 2785 2227
rect 2883 2226 2884 2251
rect 2735 2228 2736 2251
rect 2783 2228 2784 2251
rect 2787 2018 2788 2229
rect 2794 2018 2795 2229
rect 2634 2018 2635 2231
rect 2795 2230 2796 2251
rect 2580 2018 2581 2233
rect 2633 2232 2634 2251
rect 2529 2018 2530 2235
rect 2579 2234 2580 2251
rect 2460 2018 2461 2237
rect 2528 2236 2529 2251
rect 2391 2018 2392 2239
rect 2459 2238 2460 2251
rect 2390 2240 2391 2251
rect 2454 2018 2455 2241
rect 2403 2018 2404 2243
rect 2453 2242 2454 2251
rect 2145 2244 2146 2251
rect 2402 2244 2403 2251
rect 2700 2018 2701 2245
rect 2786 2244 2787 2251
rect 2792 2244 2793 2251
rect 2868 2244 2869 2251
rect 2856 2018 2857 2247
rect 2948 2246 2949 2251
rect 2702 2248 2703 2251
rect 2856 2248 2857 2251
rect 2874 2248 2875 2251
rect 2921 2248 2922 2251
rect 2045 2257 2046 2512
rect 2049 2257 2050 2512
rect 2062 2255 2063 2258
rect 2483 2255 2484 2258
rect 2066 2255 2067 2260
rect 2390 2255 2391 2260
rect 2070 2261 2071 2512
rect 2486 2255 2487 2262
rect 2080 2263 2081 2512
rect 2110 2255 2111 2264
rect 2088 2255 2089 2266
rect 2229 2265 2230 2512
rect 2089 2267 2090 2512
rect 2498 2255 2499 2268
rect 2097 2255 2098 2270
rect 2400 2269 2401 2512
rect 2098 2271 2099 2512
rect 2322 2271 2323 2512
rect 2107 2255 2108 2274
rect 2171 2255 2172 2274
rect 2107 2275 2108 2512
rect 2231 2255 2232 2276
rect 2117 2277 2118 2512
rect 2418 2277 2419 2512
rect 2125 2255 2126 2280
rect 2363 2255 2364 2280
rect 2126 2281 2127 2512
rect 2366 2255 2367 2282
rect 2129 2255 2130 2284
rect 2525 2255 2526 2284
rect 2138 2255 2139 2286
rect 2154 2285 2155 2512
rect 2141 2255 2142 2288
rect 2465 2255 2466 2288
rect 2143 2289 2144 2512
rect 2495 2255 2496 2290
rect 2157 2291 2158 2512
rect 2469 2291 2470 2512
rect 2159 2255 2160 2294
rect 2288 2255 2289 2294
rect 2135 2255 2136 2296
rect 2160 2295 2161 2512
rect 2162 2255 2163 2296
rect 2477 2255 2478 2296
rect 2152 2255 2153 2298
rect 2163 2297 2164 2512
rect 2177 2255 2178 2298
rect 2193 2297 2194 2512
rect 2187 2299 2188 2512
rect 2564 2255 2565 2300
rect 2195 2255 2196 2302
rect 2211 2301 2212 2512
rect 2199 2303 2200 2512
rect 2207 2255 2208 2304
rect 2217 2303 2218 2512
rect 2528 2255 2529 2304
rect 2219 2255 2220 2306
rect 2510 2255 2511 2306
rect 2222 2255 2223 2308
rect 2607 2307 2608 2512
rect 2243 2255 2244 2310
rect 2289 2309 2290 2512
rect 2250 2311 2251 2512
rect 2496 2311 2497 2512
rect 2255 2255 2256 2314
rect 2346 2313 2347 2512
rect 2259 2315 2260 2512
rect 2279 2255 2280 2316
rect 2267 2255 2268 2318
rect 2271 2317 2272 2512
rect 2276 2255 2277 2318
rect 2280 2317 2281 2512
rect 2273 2255 2274 2320
rect 2277 2319 2278 2512
rect 2291 2255 2292 2320
rect 2295 2319 2296 2512
rect 2304 2319 2305 2512
rect 2312 2255 2313 2320
rect 2076 2255 2077 2322
rect 2313 2321 2314 2512
rect 2306 2255 2307 2324
rect 2310 2323 2311 2512
rect 2316 2323 2317 2512
rect 2318 2255 2319 2324
rect 2324 2255 2325 2324
rect 2328 2323 2329 2512
rect 2330 2255 2331 2324
rect 2334 2323 2335 2512
rect 2340 2323 2341 2512
rect 2342 2255 2343 2324
rect 2348 2255 2349 2324
rect 2364 2323 2365 2512
rect 2352 2325 2353 2512
rect 2447 2255 2448 2326
rect 2166 2327 2167 2512
rect 2448 2327 2449 2512
rect 2358 2329 2359 2512
rect 2378 2255 2379 2330
rect 2360 2255 2361 2332
rect 2370 2331 2371 2512
rect 2361 2333 2362 2512
rect 2381 2255 2382 2334
rect 2372 2255 2373 2336
rect 2394 2335 2395 2512
rect 2122 2255 2123 2338
rect 2373 2337 2374 2512
rect 2382 2337 2383 2512
rect 2459 2255 2460 2338
rect 2148 2255 2149 2340
rect 2460 2339 2461 2512
rect 2147 2341 2148 2512
rect 2265 2341 2266 2512
rect 2384 2255 2385 2342
rect 2385 2341 2386 2512
rect 2391 2341 2392 2512
rect 2426 2255 2427 2342
rect 2247 2343 2248 2512
rect 2427 2343 2428 2512
rect 2402 2255 2403 2346
rect 2478 2345 2479 2512
rect 2406 2347 2407 2512
rect 2501 2255 2502 2348
rect 2412 2349 2413 2512
rect 2745 2349 2746 2512
rect 2424 2351 2425 2512
rect 2519 2255 2520 2352
rect 2429 2255 2430 2354
rect 2592 2353 2593 2512
rect 2436 2355 2437 2512
rect 2453 2255 2454 2356
rect 2442 2357 2443 2512
rect 2543 2255 2544 2358
rect 2136 2359 2137 2512
rect 2544 2359 2545 2512
rect 2454 2361 2455 2512
rect 2561 2255 2562 2362
rect 2466 2363 2467 2512
rect 2871 2255 2872 2364
rect 2475 2365 2476 2512
rect 2492 2255 2493 2366
rect 2484 2367 2485 2512
rect 2585 2255 2586 2368
rect 2502 2369 2503 2512
rect 2507 2255 2508 2370
rect 2420 2255 2421 2372
rect 2508 2371 2509 2512
rect 2421 2373 2422 2512
rect 2504 2255 2505 2374
rect 2520 2373 2521 2512
rect 2573 2255 2574 2374
rect 2526 2375 2527 2512
rect 2889 2255 2890 2376
rect 2550 2377 2551 2512
rect 2648 2255 2649 2378
rect 2574 2379 2575 2512
rect 2945 2255 2946 2380
rect 2609 2255 2610 2382
rect 2655 2381 2656 2512
rect 2619 2383 2620 2512
rect 2693 2255 2694 2384
rect 2621 2255 2622 2386
rect 2649 2385 2650 2512
rect 2627 2255 2628 2388
rect 2903 2387 2904 2512
rect 2628 2389 2629 2512
rect 2708 2255 2709 2390
rect 2537 2255 2538 2392
rect 2709 2391 2710 2512
rect 2414 2255 2415 2394
rect 2538 2393 2539 2512
rect 2415 2395 2416 2512
rect 2622 2395 2623 2512
rect 2631 2395 2632 2512
rect 2633 2255 2634 2396
rect 2637 2395 2638 2512
rect 2702 2255 2703 2396
rect 2555 2255 2556 2398
rect 2703 2397 2704 2512
rect 2556 2399 2557 2512
rect 2642 2255 2643 2400
rect 2639 2255 2640 2402
rect 2844 2401 2845 2512
rect 2679 2403 2680 2512
rect 2747 2255 2748 2404
rect 2588 2255 2589 2406
rect 2748 2405 2749 2512
rect 2684 2255 2685 2408
rect 2900 2407 2901 2512
rect 2471 2255 2472 2410
rect 2685 2409 2686 2512
rect 2472 2411 2473 2512
rect 2489 2255 2490 2412
rect 2490 2413 2491 2512
rect 2531 2255 2532 2414
rect 2532 2415 2533 2512
rect 2579 2255 2580 2416
rect 2580 2417 2581 2512
rect 2660 2255 2661 2418
rect 2444 2255 2445 2420
rect 2661 2419 2662 2512
rect 2445 2421 2446 2512
rect 2546 2255 2547 2422
rect 2696 2255 2697 2422
rect 2935 2421 2936 2512
rect 2697 2423 2698 2512
rect 2958 2255 2959 2424
rect 2241 2425 2242 2512
rect 2959 2425 2960 2512
rect 2700 2427 2701 2512
rect 2966 2427 2967 2512
rect 2715 2429 2716 2512
rect 2914 2255 2915 2430
rect 2729 2255 2730 2432
rect 2733 2431 2734 2512
rect 2735 2255 2736 2432
rect 2829 2431 2830 2512
rect 2738 2255 2739 2434
rect 2832 2433 2833 2512
rect 2750 2255 2751 2436
rect 2931 2435 2932 2512
rect 2396 2255 2397 2438
rect 2751 2437 2752 2512
rect 2375 2255 2376 2440
rect 2397 2439 2398 2512
rect 2100 2255 2101 2442
rect 2376 2441 2377 2512
rect 2756 2255 2757 2442
rect 2938 2255 2939 2442
rect 2757 2443 2758 2512
rect 2762 2255 2763 2444
rect 2666 2255 2667 2446
rect 2763 2445 2764 2512
rect 2667 2447 2668 2512
rect 2945 2447 2946 2512
rect 2760 2449 2761 2512
rect 2795 2255 2796 2450
rect 2771 2255 2772 2452
rect 2775 2451 2776 2512
rect 2768 2255 2769 2454
rect 2772 2453 2773 2512
rect 2784 2453 2785 2512
rect 2813 2255 2814 2454
rect 2786 2255 2787 2456
rect 2847 2455 2848 2512
rect 2597 2255 2598 2458
rect 2787 2457 2788 2512
rect 2513 2255 2514 2460
rect 2598 2459 2599 2512
rect 2789 2255 2790 2460
rect 2850 2459 2851 2512
rect 2570 2255 2571 2462
rect 2790 2461 2791 2512
rect 2796 2461 2797 2512
rect 2804 2255 2805 2462
rect 2567 2255 2568 2464
rect 2805 2463 2806 2512
rect 2568 2465 2569 2512
rect 2672 2255 2673 2466
rect 2673 2467 2674 2512
rect 2711 2255 2712 2468
rect 2798 2255 2799 2468
rect 2870 2467 2871 2512
rect 2801 2255 2802 2470
rect 2816 2255 2817 2470
rect 2811 2471 2812 2512
rect 2819 2255 2820 2472
rect 2814 2473 2815 2512
rect 2822 2255 2823 2474
rect 2817 2475 2818 2512
rect 2825 2255 2826 2476
rect 2823 2477 2824 2512
rect 2877 2255 2878 2478
rect 2837 2255 2838 2480
rect 2891 2479 2892 2512
rect 2840 2255 2841 2482
rect 2868 2255 2869 2482
rect 2792 2255 2793 2484
rect 2867 2483 2868 2512
rect 2354 2255 2355 2486
rect 2793 2485 2794 2512
rect 2355 2487 2356 2512
rect 2450 2255 2451 2488
rect 2841 2487 2842 2512
rect 2893 2255 2894 2488
rect 2852 2255 2853 2490
rect 2856 2255 2857 2490
rect 2603 2255 2604 2492
rect 2856 2491 2857 2512
rect 2408 2255 2409 2494
rect 2604 2493 2605 2512
rect 2865 2255 2866 2494
rect 2888 2493 2889 2512
rect 2874 2255 2875 2496
rect 2918 2495 2919 2512
rect 2873 2497 2874 2512
rect 2952 2497 2953 2512
rect 2880 2255 2881 2500
rect 2897 2499 2898 2512
rect 2879 2501 2880 2512
rect 2938 2501 2939 2512
rect 2883 2255 2884 2504
rect 2886 2255 2887 2504
rect 2862 2255 2863 2506
rect 2885 2505 2886 2512
rect 2615 2255 2616 2508
rect 2863 2507 2864 2512
rect 2616 2509 2617 2512
rect 2690 2255 2691 2510
rect 2915 2509 2916 2512
rect 2921 2255 2922 2510
rect 2948 2255 2949 2510
rect 2969 2509 2970 2512
rect 2035 2516 2036 2519
rect 2361 2516 2362 2519
rect 2038 2516 2039 2521
rect 2042 2516 2043 2521
rect 2049 2516 2050 2521
rect 2056 2516 2057 2521
rect 2063 2516 2064 2521
rect 2358 2516 2359 2521
rect 2080 2516 2081 2523
rect 2104 2522 2105 2801
rect 2084 2524 2085 2801
rect 2089 2516 2090 2525
rect 2093 2524 2094 2801
rect 2336 2524 2337 2801
rect 2095 2516 2096 2527
rect 2538 2516 2539 2527
rect 2098 2516 2099 2529
rect 2793 2516 2794 2529
rect 2100 2530 2101 2801
rect 2418 2516 2419 2531
rect 2110 2516 2111 2533
rect 2480 2532 2481 2801
rect 2077 2516 2078 2535
rect 2110 2534 2111 2801
rect 2114 2516 2115 2535
rect 2187 2516 2188 2535
rect 2129 2516 2130 2537
rect 2508 2516 2509 2537
rect 2133 2516 2134 2539
rect 2424 2516 2425 2539
rect 2139 2540 2140 2801
rect 2237 2540 2238 2801
rect 2142 2542 2143 2801
rect 2160 2516 2161 2543
rect 2145 2544 2146 2801
rect 2394 2516 2395 2545
rect 2147 2516 2148 2547
rect 2259 2516 2260 2547
rect 2148 2548 2149 2801
rect 2402 2548 2403 2801
rect 2176 2550 2177 2801
rect 2199 2516 2200 2551
rect 2188 2552 2189 2801
rect 2211 2516 2212 2553
rect 2206 2554 2207 2801
rect 2229 2516 2230 2555
rect 2224 2556 2225 2801
rect 2478 2516 2479 2557
rect 2227 2558 2228 2801
rect 2265 2516 2266 2559
rect 2231 2560 2232 2801
rect 2552 2560 2553 2801
rect 2243 2562 2244 2801
rect 2289 2516 2290 2563
rect 2247 2516 2248 2565
rect 2502 2516 2503 2565
rect 2255 2566 2256 2801
rect 2561 2566 2562 2801
rect 2261 2568 2262 2801
rect 2271 2516 2272 2569
rect 2267 2570 2268 2801
rect 2277 2516 2278 2571
rect 2291 2570 2292 2801
rect 2328 2516 2329 2571
rect 2297 2572 2298 2801
rect 2322 2516 2323 2573
rect 2304 2516 2305 2575
rect 2318 2574 2319 2801
rect 2303 2576 2304 2801
rect 2385 2516 2386 2577
rect 2310 2516 2311 2579
rect 2330 2578 2331 2801
rect 2316 2516 2317 2581
rect 2324 2580 2325 2801
rect 2295 2516 2296 2583
rect 2315 2582 2316 2801
rect 2340 2516 2341 2583
rect 2360 2582 2361 2801
rect 2342 2584 2343 2801
rect 2751 2516 2752 2585
rect 2352 2516 2353 2587
rect 2498 2586 2499 2801
rect 2355 2516 2356 2589
rect 2501 2588 2502 2801
rect 2334 2516 2335 2591
rect 2354 2590 2355 2801
rect 2313 2516 2314 2593
rect 2333 2592 2334 2801
rect 2366 2592 2367 2801
rect 2604 2516 2605 2593
rect 2373 2516 2374 2595
rect 2486 2594 2487 2801
rect 2364 2516 2365 2597
rect 2372 2596 2373 2801
rect 2376 2516 2377 2597
rect 2384 2596 2385 2801
rect 2375 2598 2376 2801
rect 2427 2516 2428 2599
rect 2066 2516 2067 2601
rect 2426 2600 2427 2801
rect 2391 2516 2392 2603
rect 2477 2602 2478 2801
rect 2390 2604 2391 2801
rect 2745 2516 2746 2605
rect 2406 2516 2407 2607
rect 2528 2606 2529 2801
rect 2408 2608 2409 2801
rect 2860 2516 2861 2609
rect 2412 2516 2413 2611
rect 2429 2610 2430 2801
rect 2397 2516 2398 2613
rect 2411 2612 2412 2801
rect 2370 2516 2371 2615
rect 2396 2614 2397 2801
rect 2415 2516 2416 2615
rect 2661 2516 2662 2615
rect 2400 2516 2401 2617
rect 2414 2616 2415 2801
rect 2436 2516 2437 2617
rect 2585 2616 2586 2801
rect 2435 2618 2436 2801
rect 2622 2516 2623 2619
rect 2442 2516 2443 2621
rect 2594 2620 2595 2801
rect 2166 2516 2167 2623
rect 2441 2622 2442 2801
rect 2167 2624 2168 2801
rect 2454 2516 2455 2625
rect 2448 2516 2449 2627
rect 2453 2626 2454 2801
rect 2163 2516 2164 2629
rect 2447 2628 2448 2801
rect 2164 2630 2165 2801
rect 2624 2630 2625 2801
rect 2460 2516 2461 2633
rect 2576 2632 2577 2801
rect 2466 2516 2467 2635
rect 2582 2634 2583 2801
rect 2097 2636 2098 2801
rect 2465 2636 2466 2801
rect 2472 2516 2473 2637
rect 2534 2636 2535 2801
rect 2475 2516 2476 2639
rect 2537 2638 2538 2801
rect 2474 2640 2475 2801
rect 2832 2516 2833 2641
rect 2490 2516 2491 2643
rect 2546 2642 2547 2801
rect 2489 2644 2490 2801
rect 2685 2516 2686 2645
rect 2496 2516 2497 2647
rect 2935 2516 2936 2647
rect 2382 2516 2383 2649
rect 2495 2648 2496 2801
rect 2510 2648 2511 2801
rect 2709 2516 2710 2649
rect 2516 2650 2517 2801
rect 2835 2650 2836 2801
rect 2520 2516 2521 2653
rect 2735 2652 2736 2801
rect 2522 2654 2523 2801
rect 2598 2516 2599 2655
rect 2445 2516 2446 2657
rect 2597 2656 2598 2801
rect 2544 2516 2545 2659
rect 2558 2658 2559 2801
rect 2568 2516 2569 2659
rect 2720 2658 2721 2801
rect 2567 2660 2568 2801
rect 2784 2516 2785 2661
rect 2570 2662 2571 2801
rect 2703 2516 2704 2663
rect 2550 2516 2551 2665
rect 2702 2664 2703 2801
rect 2574 2516 2575 2667
rect 2726 2666 2727 2801
rect 2592 2516 2593 2669
rect 2877 2668 2878 2801
rect 2607 2516 2608 2671
rect 2805 2516 2806 2671
rect 2532 2516 2533 2673
rect 2606 2672 2607 2801
rect 2421 2516 2422 2675
rect 2531 2674 2532 2801
rect 2420 2676 2421 2801
rect 2715 2516 2716 2677
rect 2580 2516 2581 2679
rect 2714 2678 2715 2801
rect 2612 2680 2613 2801
rect 2655 2516 2656 2681
rect 2616 2516 2617 2683
rect 2711 2682 2712 2801
rect 2619 2516 2620 2685
rect 2690 2684 2691 2801
rect 2618 2686 2619 2801
rect 2856 2516 2857 2687
rect 2628 2516 2629 2689
rect 2750 2688 2751 2801
rect 2346 2516 2347 2691
rect 2627 2690 2628 2801
rect 2639 2690 2640 2801
rect 2748 2516 2749 2691
rect 2654 2692 2655 2801
rect 2891 2516 2892 2693
rect 2657 2694 2658 2801
rect 2760 2516 2761 2695
rect 2621 2696 2622 2801
rect 2759 2696 2760 2801
rect 2667 2516 2668 2699
rect 2906 2516 2907 2699
rect 2673 2516 2674 2701
rect 2945 2516 2946 2701
rect 2526 2516 2527 2703
rect 2672 2702 2673 2801
rect 2525 2704 2526 2801
rect 2829 2516 2830 2705
rect 2679 2516 2680 2707
rect 2938 2706 2939 2801
rect 2469 2516 2470 2709
rect 2678 2708 2679 2801
rect 2280 2516 2281 2711
rect 2468 2710 2469 2801
rect 2129 2712 2130 2801
rect 2279 2712 2280 2801
rect 2684 2712 2685 2801
rect 2733 2516 2734 2713
rect 2697 2516 2698 2715
rect 2982 2516 2983 2715
rect 2556 2516 2557 2717
rect 2696 2716 2697 2801
rect 2700 2516 2701 2717
rect 2979 2516 2980 2717
rect 2708 2718 2709 2801
rect 2891 2718 2892 2801
rect 2732 2720 2733 2801
rect 2847 2516 2848 2721
rect 2738 2722 2739 2801
rect 2972 2516 2973 2723
rect 2744 2724 2745 2801
rect 2912 2724 2913 2801
rect 2757 2516 2758 2727
rect 2863 2516 2864 2727
rect 2763 2516 2764 2729
rect 2894 2516 2895 2729
rect 2631 2516 2632 2731
rect 2894 2730 2895 2801
rect 2630 2732 2631 2801
rect 2649 2516 2650 2733
rect 2648 2734 2649 2801
rect 2900 2516 2901 2735
rect 2637 2516 2638 2737
rect 2901 2736 2902 2801
rect 2484 2516 2485 2739
rect 2636 2738 2637 2801
rect 2126 2516 2127 2741
rect 2483 2740 2484 2801
rect 2125 2742 2126 2801
rect 2193 2516 2194 2743
rect 2194 2744 2195 2801
rect 2217 2516 2218 2745
rect 2218 2746 2219 2801
rect 2241 2516 2242 2747
rect 2772 2516 2773 2747
rect 2777 2746 2778 2801
rect 2783 2746 2784 2801
rect 2796 2516 2797 2747
rect 2787 2516 2788 2749
rect 2853 2516 2854 2749
rect 2786 2750 2787 2801
rect 2966 2516 2967 2751
rect 2792 2752 2793 2801
rect 2844 2516 2845 2753
rect 2122 2754 2123 2801
rect 2844 2754 2845 2801
rect 2795 2756 2796 2801
rect 2811 2516 2812 2757
rect 2154 2516 2155 2759
rect 2810 2758 2811 2801
rect 2798 2760 2799 2801
rect 2814 2516 2815 2761
rect 2790 2516 2791 2763
rect 2814 2762 2815 2801
rect 2789 2764 2790 2801
rect 2841 2516 2842 2765
rect 2801 2766 2802 2801
rect 2823 2516 2824 2767
rect 2808 2516 2809 2769
rect 2838 2516 2839 2769
rect 2807 2770 2808 2801
rect 2850 2516 2851 2771
rect 2817 2516 2818 2773
rect 2963 2516 2964 2773
rect 2820 2774 2821 2801
rect 2885 2516 2886 2775
rect 2823 2776 2824 2801
rect 2888 2516 2889 2777
rect 2826 2778 2827 2801
rect 2908 2778 2909 2801
rect 2829 2780 2830 2801
rect 2873 2516 2874 2781
rect 2841 2782 2842 2801
rect 2897 2516 2898 2783
rect 2859 2784 2860 2801
rect 2942 2516 2943 2785
rect 2862 2786 2863 2801
rect 2928 2786 2929 2801
rect 2871 2788 2872 2801
rect 2915 2516 2916 2789
rect 2775 2516 2776 2791
rect 2915 2790 2916 2801
rect 2874 2792 2875 2801
rect 2918 2516 2919 2793
rect 2879 2516 2880 2795
rect 2949 2516 2950 2795
rect 2918 2796 2919 2801
rect 2969 2516 2970 2797
rect 2935 2798 2936 2801
rect 2942 2798 2943 2801
rect 2059 2807 2060 3086
rect 2154 2807 2155 3086
rect 2065 2805 2066 2810
rect 2480 2805 2481 2810
rect 2068 2805 2069 2812
rect 2084 2805 2085 2812
rect 2069 2813 2070 3086
rect 2110 2805 2111 2814
rect 2075 2805 2076 2816
rect 2261 2805 2262 2816
rect 2076 2817 2077 3086
rect 2495 2805 2496 2818
rect 2083 2819 2084 3086
rect 2465 2805 2466 2820
rect 2087 2821 2088 3086
rect 2426 2805 2427 2822
rect 2093 2805 2094 2824
rect 2627 2805 2628 2824
rect 2094 2825 2095 3086
rect 2188 2805 2189 2826
rect 2097 2827 2098 3086
rect 2477 2805 2478 2828
rect 2104 2805 2105 2830
rect 2525 2805 2526 2830
rect 2119 2831 2120 3086
rect 2372 2805 2373 2832
rect 2122 2805 2123 2834
rect 2333 2805 2334 2834
rect 2125 2805 2126 2836
rect 2396 2805 2397 2836
rect 2080 2837 2081 3086
rect 2125 2837 2126 3086
rect 2129 2805 2130 2838
rect 2468 2805 2469 2838
rect 2112 2839 2113 3086
rect 2469 2839 2470 3086
rect 2131 2841 2132 3086
rect 2447 2805 2448 2842
rect 2136 2805 2137 2844
rect 2384 2805 2385 2844
rect 2135 2845 2136 3086
rect 2214 2845 2215 3086
rect 2142 2805 2143 2848
rect 2157 2847 2158 3086
rect 2142 2849 2143 3086
rect 2534 2805 2535 2850
rect 2145 2805 2146 2852
rect 2334 2851 2335 3086
rect 2145 2853 2146 3086
rect 2582 2805 2583 2854
rect 2160 2855 2161 3086
rect 2486 2805 2487 2856
rect 2163 2857 2164 3086
rect 2194 2805 2195 2858
rect 2167 2805 2168 2860
rect 2594 2805 2595 2860
rect 2176 2805 2177 2862
rect 2190 2861 2191 3086
rect 2178 2863 2179 3086
rect 2218 2805 2219 2864
rect 2196 2865 2197 3086
rect 2366 2805 2367 2866
rect 2199 2867 2200 3086
rect 2624 2805 2625 2868
rect 2202 2869 2203 3086
rect 2243 2805 2244 2870
rect 2206 2805 2207 2872
rect 2289 2871 2290 3086
rect 2208 2873 2209 3086
rect 2237 2805 2238 2874
rect 2220 2875 2221 3086
rect 2406 2875 2407 3086
rect 2224 2805 2225 2878
rect 2706 2877 2707 3086
rect 2223 2879 2224 3086
rect 2639 2805 2640 2880
rect 2227 2805 2228 2882
rect 2328 2881 2329 3086
rect 2231 2805 2232 2884
rect 2435 2805 2436 2884
rect 2152 2805 2153 2886
rect 2436 2885 2437 3086
rect 2232 2887 2233 3086
rect 2267 2805 2268 2888
rect 2244 2889 2245 3086
rect 2279 2805 2280 2890
rect 2262 2891 2263 3086
rect 2291 2805 2292 2892
rect 2268 2893 2269 3086
rect 2315 2805 2316 2894
rect 2271 2895 2272 3086
rect 2318 2805 2319 2896
rect 2277 2897 2278 3086
rect 2324 2805 2325 2898
rect 2283 2899 2284 3086
rect 2330 2805 2331 2900
rect 2286 2901 2287 3086
rect 2336 2805 2337 2902
rect 2297 2805 2298 2904
rect 2394 2903 2395 3086
rect 2303 2805 2304 2906
rect 2331 2905 2332 3086
rect 2304 2907 2305 3086
rect 2354 2805 2355 2908
rect 2310 2909 2311 3086
rect 2360 2805 2361 2910
rect 2313 2911 2314 3086
rect 2375 2805 2376 2912
rect 2072 2805 2073 2914
rect 2376 2913 2377 3086
rect 2322 2915 2323 3086
rect 2342 2805 2343 2916
rect 2340 2917 2341 3086
rect 2498 2805 2499 2918
rect 2343 2919 2344 3086
rect 2501 2805 2502 2920
rect 2346 2921 2347 3086
rect 2402 2805 2403 2922
rect 2352 2923 2353 3086
rect 2414 2805 2415 2924
rect 2355 2925 2356 3086
rect 2597 2805 2598 2926
rect 2358 2927 2359 3086
rect 2408 2805 2409 2928
rect 2364 2929 2365 3086
rect 2420 2805 2421 2930
rect 2370 2931 2371 3086
rect 2429 2805 2430 2932
rect 2379 2933 2380 3086
rect 2453 2805 2454 2934
rect 2382 2935 2383 3086
rect 2537 2805 2538 2936
rect 2385 2937 2386 3086
rect 2390 2805 2391 2938
rect 2391 2939 2392 3086
rect 2483 2805 2484 2940
rect 2397 2941 2398 3086
rect 2528 2805 2529 2942
rect 2400 2943 2401 3086
rect 2531 2805 2532 2944
rect 2403 2945 2404 3086
rect 2762 2805 2763 2946
rect 2411 2805 2412 2948
rect 2439 2947 2440 3086
rect 2424 2949 2425 3086
rect 2489 2805 2490 2950
rect 2430 2951 2431 3086
rect 2516 2805 2517 2952
rect 2441 2805 2442 2954
rect 2484 2953 2485 3086
rect 2442 2955 2443 3086
rect 2576 2805 2577 2956
rect 2445 2957 2446 3086
rect 2585 2805 2586 2958
rect 2448 2959 2449 3086
rect 2522 2805 2523 2960
rect 2454 2961 2455 3086
rect 2552 2805 2553 2962
rect 2460 2963 2461 3086
rect 2546 2805 2547 2964
rect 2466 2965 2467 3086
rect 2636 2805 2637 2966
rect 2472 2967 2473 3086
rect 2558 2805 2559 2968
rect 2474 2805 2475 2970
rect 2481 2969 2482 3086
rect 2475 2971 2476 3086
rect 2561 2805 2562 2972
rect 2478 2973 2479 3086
rect 2510 2805 2511 2974
rect 2490 2975 2491 3086
rect 2735 2805 2736 2976
rect 2496 2977 2497 3086
rect 2810 2805 2811 2978
rect 2508 2979 2509 3086
rect 2630 2805 2631 2980
rect 2514 2981 2515 3086
rect 2730 2981 2731 3086
rect 2526 2983 2527 3086
rect 2877 2805 2878 2984
rect 2532 2985 2533 3086
rect 2696 2805 2697 2986
rect 2544 2987 2545 3086
rect 2702 2805 2703 2988
rect 2550 2989 2551 3086
rect 2894 2805 2895 2990
rect 2553 2991 2554 3086
rect 2708 2805 2709 2992
rect 2556 2993 2557 3086
rect 2612 2805 2613 2994
rect 2562 2995 2563 3086
rect 2720 2805 2721 2996
rect 2567 2805 2568 2998
rect 2688 2997 2689 3086
rect 2241 2999 2242 3086
rect 2568 2999 2569 3086
rect 2570 2805 2571 3000
rect 2759 2805 2760 3000
rect 2574 3001 2575 3086
rect 2838 2805 2839 3002
rect 2580 3003 2581 3086
rect 2648 2805 2649 3004
rect 2592 3005 2593 3086
rect 2853 3005 2854 3086
rect 2595 3007 2596 3086
rect 2846 3007 2847 3086
rect 2598 3009 2599 3086
rect 2901 2805 2902 3010
rect 2604 3011 2605 3086
rect 2744 2805 2745 3012
rect 2606 2805 2607 3014
rect 2718 3013 2719 3086
rect 2610 3015 2611 3086
rect 2750 2805 2751 3016
rect 2613 3017 2614 3086
rect 2823 2805 2824 3018
rect 2618 2805 2619 3020
rect 2817 2805 2818 3020
rect 2631 3021 2632 3086
rect 2654 2805 2655 3022
rect 2634 3023 2635 3086
rect 2657 2805 2658 3024
rect 2637 3025 2638 3086
rect 2850 2805 2851 3026
rect 2643 3027 2644 3086
rect 2697 3027 2698 3086
rect 2672 2805 2673 3030
rect 2835 2805 2836 3030
rect 2673 3031 2674 3086
rect 2798 2805 2799 3032
rect 2676 3033 2677 3086
rect 2684 2805 2685 3034
rect 2621 2805 2622 3036
rect 2685 3035 2686 3086
rect 2678 2805 2679 3038
rect 2757 3037 2758 3086
rect 2679 3039 2680 3086
rect 2783 2805 2784 3040
rect 2682 3041 2683 3086
rect 2786 2805 2787 3042
rect 2502 3043 2503 3086
rect 2785 3043 2786 3086
rect 2690 2805 2691 3046
rect 2891 2805 2892 3046
rect 2691 3047 2692 3086
rect 2844 2805 2845 3048
rect 2703 3049 2704 3086
rect 2732 2805 2733 3050
rect 2709 3051 2710 3086
rect 2789 2805 2790 3052
rect 2711 2805 2712 3054
rect 2788 3053 2789 3086
rect 2712 3055 2713 3086
rect 2792 2805 2793 3056
rect 2733 3057 2734 3086
rect 2820 2805 2821 3058
rect 2736 3059 2737 3086
rect 2748 3059 2749 3086
rect 2738 2805 2739 3062
rect 2912 2805 2913 3062
rect 2739 3063 2740 3086
rect 2826 2805 2827 3064
rect 2754 3065 2755 3086
rect 2841 2805 2842 3066
rect 2760 3067 2761 3086
rect 2862 2805 2863 3068
rect 2763 3069 2764 3086
rect 2777 2805 2778 3070
rect 2772 3071 2773 3086
rect 2871 2805 2872 3072
rect 2775 3073 2776 3086
rect 2874 2805 2875 3074
rect 2781 3075 2782 3086
rect 2795 2805 2796 3076
rect 2801 2805 2802 3076
rect 2884 2805 2885 3076
rect 2826 3077 2827 3086
rect 2918 2805 2919 3078
rect 2829 2805 2830 3080
rect 2938 2805 2939 3080
rect 2726 2805 2727 3082
rect 2829 3081 2830 3086
rect 2714 2805 2715 3084
rect 2727 3083 2728 3086
rect 2859 2805 2860 3084
rect 2931 2805 2932 3084
rect 2062 3090 2063 3093
rect 2190 3090 2191 3093
rect 2065 3094 2066 3323
rect 2374 3094 2375 3323
rect 2087 3090 2088 3097
rect 2277 3090 2278 3097
rect 2097 3090 2098 3099
rect 2289 3090 2290 3099
rect 2079 3100 2080 3323
rect 2098 3100 2099 3323
rect 2101 3100 2102 3323
rect 2304 3090 2305 3101
rect 2104 3102 2105 3323
rect 2125 3090 2126 3103
rect 2110 3104 2111 3323
rect 2400 3090 2401 3105
rect 2115 3090 2116 3107
rect 2394 3090 2395 3107
rect 2073 3090 2074 3109
rect 2395 3108 2396 3323
rect 2114 3110 2115 3323
rect 2313 3090 2314 3111
rect 2120 3112 2121 3323
rect 2154 3090 2155 3113
rect 2123 3114 2124 3323
rect 2157 3090 2158 3115
rect 2126 3116 2127 3323
rect 2346 3090 2347 3117
rect 2135 3090 2136 3119
rect 2176 3118 2177 3323
rect 2138 3090 2139 3121
rect 2208 3090 2209 3121
rect 2142 3090 2143 3123
rect 2262 3090 2263 3123
rect 2141 3124 2142 3323
rect 2305 3124 2306 3323
rect 2145 3090 2146 3127
rect 2442 3090 2443 3127
rect 2157 3128 2158 3323
rect 2178 3090 2179 3129
rect 2173 3130 2174 3323
rect 2281 3130 2282 3323
rect 2182 3132 2183 3323
rect 2214 3090 2215 3133
rect 2202 3090 2203 3135
rect 2368 3134 2369 3323
rect 2218 3136 2219 3323
rect 2244 3090 2245 3137
rect 2224 3138 2225 3323
rect 2355 3090 2356 3139
rect 2232 3090 2233 3141
rect 2362 3140 2363 3323
rect 2236 3142 2237 3323
rect 2385 3090 2386 3143
rect 2238 3090 2239 3145
rect 2382 3090 2383 3145
rect 2241 3090 2242 3147
rect 2472 3090 2473 3147
rect 2242 3148 2243 3323
rect 2268 3090 2269 3149
rect 2263 3150 2264 3323
rect 2286 3090 2287 3151
rect 2269 3152 2270 3323
rect 2310 3090 2311 3153
rect 2138 3154 2139 3323
rect 2311 3154 2312 3323
rect 2283 3090 2284 3157
rect 2410 3156 2411 3323
rect 2293 3158 2294 3323
rect 2328 3090 2329 3159
rect 2296 3160 2297 3323
rect 2331 3090 2332 3161
rect 2317 3162 2318 3323
rect 2358 3090 2359 3163
rect 2083 3090 2084 3165
rect 2359 3164 2360 3323
rect 2329 3166 2330 3323
rect 2334 3090 2335 3167
rect 2335 3168 2336 3323
rect 2340 3090 2341 3169
rect 2338 3170 2339 3323
rect 2343 3090 2344 3171
rect 2341 3172 2342 3323
rect 2370 3090 2371 3173
rect 2347 3174 2348 3323
rect 2364 3090 2365 3175
rect 2365 3176 2366 3323
rect 2379 3090 2380 3177
rect 2371 3178 2372 3323
rect 2376 3090 2377 3179
rect 2383 3178 2384 3323
rect 2406 3090 2407 3179
rect 2072 3180 2073 3323
rect 2407 3180 2408 3323
rect 2389 3182 2390 3323
rect 2391 3090 2392 3183
rect 2112 3090 2113 3185
rect 2392 3184 2393 3323
rect 2397 3090 2398 3185
rect 2401 3184 2402 3323
rect 2076 3090 2077 3187
rect 2398 3186 2399 3323
rect 2075 3188 2076 3323
rect 2271 3090 2272 3189
rect 2403 3090 2404 3189
rect 2413 3188 2414 3323
rect 2094 3090 2095 3191
rect 2404 3190 2405 3323
rect 2094 3192 2095 3323
rect 2272 3192 2273 3323
rect 2422 3192 2423 3323
rect 2478 3090 2479 3193
rect 2428 3194 2429 3323
rect 2445 3090 2446 3195
rect 2436 3090 2437 3197
rect 2443 3196 2444 3323
rect 2424 3090 2425 3199
rect 2437 3198 2438 3323
rect 2439 3090 2440 3199
rect 2446 3198 2447 3323
rect 2448 3090 2449 3199
rect 2650 3198 2651 3323
rect 2160 3090 2161 3201
rect 2449 3200 2450 3323
rect 2466 3090 2467 3201
rect 2473 3200 2474 3323
rect 2460 3090 2461 3203
rect 2467 3202 2468 3323
rect 2454 3090 2455 3205
rect 2461 3204 2462 3323
rect 2430 3090 2431 3207
rect 2455 3206 2456 3323
rect 2131 3090 2132 3209
rect 2431 3208 2432 3323
rect 2479 3208 2480 3323
rect 2653 3208 2654 3323
rect 2481 3090 2482 3211
rect 2482 3210 2483 3323
rect 2490 3090 2491 3211
rect 2718 3090 2719 3211
rect 2287 3212 2288 3323
rect 2491 3212 2492 3323
rect 2496 3090 2497 3213
rect 2730 3090 2731 3213
rect 2484 3090 2485 3215
rect 2497 3214 2498 3323
rect 2502 3090 2503 3215
rect 2696 3214 2697 3323
rect 2503 3216 2504 3323
rect 2508 3090 2509 3217
rect 2521 3216 2522 3323
rect 2712 3090 2713 3217
rect 2524 3218 2525 3323
rect 2568 3090 2569 3219
rect 2532 3090 2533 3221
rect 2539 3220 2540 3323
rect 2536 3222 2537 3323
rect 2550 3090 2551 3223
rect 2542 3224 2543 3323
rect 2544 3090 2545 3225
rect 2553 3090 2554 3225
rect 2820 3090 2821 3225
rect 2554 3226 2555 3323
rect 2580 3090 2581 3227
rect 2556 3090 2557 3229
rect 2711 3228 2712 3323
rect 2560 3230 2561 3323
rect 2562 3090 2563 3231
rect 2572 3230 2573 3323
rect 2631 3090 2632 3231
rect 2574 3090 2575 3233
rect 2660 3232 2661 3323
rect 2575 3234 2576 3323
rect 2634 3090 2635 3235
rect 2578 3236 2579 3323
rect 2669 3236 2670 3323
rect 2590 3238 2591 3323
rect 2800 3238 2801 3323
rect 2592 3090 2593 3241
rect 2846 3090 2847 3241
rect 2593 3242 2594 3323
rect 2610 3090 2611 3243
rect 2595 3090 2596 3245
rect 2839 3090 2840 3245
rect 2475 3090 2476 3247
rect 2596 3246 2597 3323
rect 2469 3090 2470 3249
rect 2476 3248 2477 3323
rect 2598 3090 2599 3249
rect 2836 3090 2837 3249
rect 2322 3090 2323 3251
rect 2599 3250 2600 3323
rect 2323 3252 2324 3323
rect 2352 3090 2353 3253
rect 2128 3090 2129 3255
rect 2353 3254 2354 3323
rect 2129 3256 2130 3323
rect 2434 3256 2435 3323
rect 2602 3256 2603 3323
rect 2832 3090 2833 3257
rect 2604 3090 2605 3259
rect 2803 3258 2804 3323
rect 2613 3090 2614 3261
rect 2720 3260 2721 3323
rect 2620 3262 2621 3323
rect 2685 3090 2686 3263
rect 2623 3264 2624 3323
rect 2643 3090 2644 3265
rect 2632 3266 2633 3323
rect 2806 3090 2807 3267
rect 2635 3268 2636 3323
rect 2823 3090 2824 3269
rect 2641 3270 2642 3323
rect 2682 3090 2683 3271
rect 2644 3272 2645 3323
rect 2741 3272 2742 3323
rect 2663 3274 2664 3323
rect 2703 3090 2704 3275
rect 2666 3276 2667 3323
rect 2706 3090 2707 3277
rect 2673 3090 2674 3279
rect 2777 3278 2778 3323
rect 2676 3090 2677 3281
rect 2809 3090 2810 3281
rect 2675 3282 2676 3323
rect 2787 3282 2788 3323
rect 2681 3284 2682 3323
rect 2817 3284 2818 3323
rect 2684 3286 2685 3323
rect 2813 3090 2814 3287
rect 2688 3090 2689 3289
rect 2700 3090 2701 3289
rect 2702 3288 2703 3323
rect 2791 3288 2792 3323
rect 2709 3090 2710 3291
rect 2784 3290 2785 3323
rect 2708 3292 2709 3323
rect 2733 3090 2734 3293
rect 2723 3294 2724 3323
rect 2748 3090 2749 3295
rect 2726 3296 2727 3323
rect 2754 3090 2755 3297
rect 2729 3298 2730 3323
rect 2757 3090 2758 3299
rect 2732 3300 2733 3323
rect 2760 3090 2761 3301
rect 2514 3090 2515 3303
rect 2759 3302 2760 3323
rect 2515 3304 2516 3323
rect 2637 3090 2638 3305
rect 2638 3306 2639 3323
rect 2679 3090 2680 3307
rect 2736 3090 2737 3307
rect 2751 3090 2752 3307
rect 2735 3308 2736 3323
rect 2763 3090 2764 3309
rect 2739 3090 2740 3311
rect 2766 3310 2767 3323
rect 2691 3090 2692 3313
rect 2738 3312 2739 3323
rect 2690 3314 2691 3323
rect 2780 3314 2781 3323
rect 2750 3316 2751 3323
rect 2772 3090 2773 3317
rect 2526 3090 2527 3319
rect 2773 3318 2774 3323
rect 2753 3320 2754 3323
rect 2775 3090 2776 3321
rect 2797 3320 2798 3323
rect 2826 3090 2827 3321
rect 2011 3327 2012 3330
rect 2338 3327 2339 3330
rect 2065 3327 2066 3332
rect 2395 3327 2396 3332
rect 2068 3327 2069 3334
rect 2267 3333 2268 3548
rect 2068 3335 2069 3548
rect 2398 3327 2399 3336
rect 2072 3327 2073 3338
rect 2138 3327 2139 3338
rect 2079 3327 2080 3340
rect 2389 3327 2390 3340
rect 2082 3327 2083 3342
rect 2387 3341 2388 3548
rect 2094 3327 2095 3344
rect 2263 3327 2264 3344
rect 2098 3327 2099 3346
rect 2252 3345 2253 3548
rect 2108 3347 2109 3548
rect 2120 3327 2121 3348
rect 2114 3327 2115 3350
rect 2261 3349 2262 3548
rect 2041 3351 2042 3548
rect 2114 3351 2115 3548
rect 2117 3327 2118 3352
rect 2272 3327 2273 3352
rect 2117 3353 2118 3548
rect 2123 3327 2124 3354
rect 2120 3355 2121 3548
rect 2309 3355 2310 3548
rect 2126 3327 2127 3358
rect 2323 3327 2324 3358
rect 2127 3359 2128 3548
rect 2218 3327 2219 3360
rect 2129 3327 2130 3362
rect 2148 3327 2149 3362
rect 2141 3327 2142 3364
rect 2285 3363 2286 3548
rect 2166 3327 2167 3366
rect 2392 3327 2393 3366
rect 2153 3367 2154 3548
rect 2393 3367 2394 3548
rect 2157 3327 2158 3370
rect 2165 3369 2166 3548
rect 2156 3371 2157 3548
rect 2585 3371 2586 3548
rect 2171 3373 2172 3548
rect 2368 3327 2369 3374
rect 2173 3327 2174 3376
rect 2296 3327 2297 3376
rect 2174 3377 2175 3548
rect 2663 3327 2664 3378
rect 2176 3327 2177 3380
rect 2287 3327 2288 3380
rect 2177 3381 2178 3548
rect 2182 3327 2183 3382
rect 2207 3381 2208 3548
rect 2449 3327 2450 3382
rect 2224 3327 2225 3384
rect 2234 3383 2235 3548
rect 2225 3385 2226 3548
rect 2242 3327 2243 3386
rect 2228 3387 2229 3548
rect 2410 3327 2411 3388
rect 2210 3389 2211 3548
rect 2411 3389 2412 3548
rect 2239 3327 2240 3392
rect 2357 3391 2358 3548
rect 2243 3393 2244 3548
rect 2365 3327 2366 3394
rect 2258 3395 2259 3548
rect 2269 3327 2270 3396
rect 2104 3327 2105 3398
rect 2270 3397 2271 3548
rect 2279 3397 2280 3548
rect 2293 3327 2294 3398
rect 2281 3327 2282 3400
rect 2282 3399 2283 3548
rect 2291 3399 2292 3548
rect 2305 3327 2306 3400
rect 2297 3401 2298 3548
rect 2311 3327 2312 3402
rect 2303 3403 2304 3548
rect 2317 3327 2318 3404
rect 2312 3405 2313 3548
rect 2329 3327 2330 3406
rect 2324 3407 2325 3548
rect 2341 3327 2342 3408
rect 2330 3409 2331 3548
rect 2347 3327 2348 3410
rect 2335 3327 2336 3412
rect 2336 3411 2337 3548
rect 2339 3411 2340 3548
rect 2353 3327 2354 3412
rect 2345 3413 2346 3548
rect 2359 3327 2360 3414
rect 2351 3415 2352 3548
rect 2383 3327 2384 3416
rect 2362 3327 2363 3418
rect 2390 3417 2391 3548
rect 2363 3419 2364 3548
rect 2437 3327 2438 3420
rect 2369 3421 2370 3548
rect 2371 3327 2372 3422
rect 2372 3423 2373 3548
rect 2374 3327 2375 3424
rect 2375 3425 2376 3548
rect 2401 3327 2402 3426
rect 2087 3427 2088 3548
rect 2402 3427 2403 3548
rect 2378 3429 2379 3548
rect 2404 3327 2405 3430
rect 2396 3431 2397 3548
rect 2428 3327 2429 3432
rect 2399 3433 2400 3548
rect 2413 3327 2414 3434
rect 2405 3435 2406 3548
rect 2407 3327 2408 3436
rect 2075 3327 2076 3438
rect 2408 3437 2409 3548
rect 2429 3437 2430 3548
rect 2431 3327 2432 3438
rect 2432 3439 2433 3548
rect 2434 3327 2435 3440
rect 2435 3441 2436 3548
rect 2461 3327 2462 3442
rect 2441 3443 2442 3548
rect 2491 3327 2492 3444
rect 2446 3327 2447 3446
rect 2450 3445 2451 3548
rect 2443 3327 2444 3448
rect 2447 3447 2448 3548
rect 2453 3447 2454 3548
rect 2467 3327 2468 3448
rect 2455 3327 2456 3450
rect 2650 3327 2651 3450
rect 2465 3451 2466 3548
rect 2669 3327 2670 3452
rect 2471 3453 2472 3548
rect 2473 3327 2474 3454
rect 2474 3455 2475 3548
rect 2476 3327 2477 3456
rect 2240 3457 2241 3548
rect 2477 3457 2478 3548
rect 2482 3327 2483 3458
rect 2501 3457 2502 3548
rect 2483 3459 2484 3548
rect 2696 3327 2697 3460
rect 2489 3461 2490 3548
rect 2596 3327 2597 3462
rect 2492 3463 2493 3548
rect 2599 3327 2600 3464
rect 2495 3465 2496 3548
rect 2711 3327 2712 3466
rect 2497 3327 2498 3468
rect 2612 3467 2613 3548
rect 2507 3469 2508 3548
rect 2723 3327 2724 3470
rect 2515 3327 2516 3472
rect 2660 3327 2661 3472
rect 2521 3327 2522 3474
rect 2528 3473 2529 3548
rect 2542 3327 2543 3474
rect 2549 3473 2550 3548
rect 2543 3475 2544 3548
rect 2572 3327 2573 3476
rect 2546 3477 2547 3548
rect 2575 3327 2576 3478
rect 2554 3327 2555 3480
rect 2737 3479 2738 3548
rect 2539 3327 2540 3482
rect 2555 3481 2556 3548
rect 2560 3327 2561 3482
rect 2567 3481 2568 3548
rect 2578 3327 2579 3482
rect 2657 3327 2658 3482
rect 2593 3327 2594 3484
rect 2606 3483 2607 3548
rect 2609 3483 2610 3548
rect 2666 3327 2667 3484
rect 2503 3327 2504 3486
rect 2667 3485 2668 3548
rect 2422 3327 2423 3488
rect 2504 3487 2505 3548
rect 2423 3489 2424 3548
rect 2479 3327 2480 3490
rect 2620 3327 2621 3490
rect 2657 3489 2658 3548
rect 2623 3327 2624 3492
rect 2648 3491 2649 3548
rect 2627 3493 2628 3548
rect 2780 3327 2781 3494
rect 2519 3495 2520 3548
rect 2780 3495 2781 3548
rect 2630 3497 2631 3548
rect 2635 3327 2636 3498
rect 2632 3327 2633 3500
rect 2777 3327 2778 3500
rect 2633 3501 2634 3548
rect 2638 3327 2639 3502
rect 2636 3503 2637 3548
rect 2641 3327 2642 3504
rect 2639 3505 2640 3548
rect 2740 3505 2741 3548
rect 2644 3327 2645 3508
rect 2832 3507 2833 3548
rect 2645 3509 2646 3548
rect 2660 3509 2661 3548
rect 2675 3327 2676 3510
rect 2695 3509 2696 3548
rect 2702 3327 2703 3510
rect 2713 3509 2714 3548
rect 2701 3511 2702 3548
rect 2811 3511 2812 3548
rect 2720 3327 2721 3514
rect 2804 3513 2805 3548
rect 2726 3327 2727 3516
rect 2743 3515 2744 3548
rect 2725 3517 2726 3548
rect 2759 3327 2760 3518
rect 2729 3327 2730 3520
rect 2746 3519 2747 3548
rect 2708 3327 2709 3522
rect 2728 3521 2729 3548
rect 2690 3327 2691 3524
rect 2707 3523 2708 3548
rect 2750 3327 2751 3524
rect 2761 3523 2762 3548
rect 2732 3327 2733 3526
rect 2749 3525 2750 3548
rect 2753 3327 2754 3526
rect 2764 3525 2765 3548
rect 2735 3327 2736 3528
rect 2752 3527 2753 3548
rect 2734 3529 2735 3548
rect 2787 3529 2788 3548
rect 2767 3531 2768 3548
rect 2807 3327 2808 3532
rect 2684 3327 2685 3534
rect 2808 3533 2809 3548
rect 2773 3327 2774 3536
rect 2784 3327 2785 3536
rect 2264 3537 2265 3548
rect 2773 3537 2774 3548
rect 2674 3539 2675 3548
rect 2783 3539 2784 3548
rect 2797 3327 2798 3540
rect 2838 3539 2839 3548
rect 2677 3541 2678 3548
rect 2797 3541 2798 3548
rect 2817 3327 2818 3542
rect 2825 3541 2826 3548
rect 2814 3327 2815 3544
rect 2818 3543 2819 3548
rect 2731 3545 2732 3548
rect 2815 3545 2816 3548
rect 2038 3554 2039 3797
rect 2225 3552 2226 3555
rect 2044 3552 2045 3557
rect 2108 3552 2109 3557
rect 2052 3558 2053 3797
rect 2059 3558 2060 3797
rect 2056 3560 2057 3797
rect 2345 3552 2346 3561
rect 2066 3562 2067 3797
rect 2270 3552 2271 3563
rect 2072 3552 2073 3565
rect 2429 3552 2430 3565
rect 2068 3552 2069 3567
rect 2073 3566 2074 3797
rect 2084 3552 2085 3567
rect 2390 3552 2391 3567
rect 2084 3568 2085 3797
rect 2199 3568 2200 3797
rect 2094 3570 2095 3797
rect 2402 3552 2403 3571
rect 2102 3552 2103 3573
rect 2378 3552 2379 3573
rect 2105 3552 2106 3575
rect 2220 3574 2221 3797
rect 2106 3576 2107 3797
rect 2375 3552 2376 3577
rect 2110 3578 2111 3797
rect 2252 3552 2253 3579
rect 2114 3552 2115 3581
rect 2123 3580 2124 3797
rect 2117 3552 2118 3583
rect 2126 3582 2127 3797
rect 2117 3584 2118 3797
rect 2277 3584 2278 3797
rect 2130 3552 2131 3587
rect 2289 3586 2290 3797
rect 2129 3588 2130 3797
rect 2655 3588 2656 3797
rect 2132 3590 2133 3797
rect 2234 3552 2235 3591
rect 2134 3552 2135 3593
rect 2253 3592 2254 3797
rect 2137 3552 2138 3595
rect 2483 3552 2484 3595
rect 2139 3596 2140 3797
rect 2291 3552 2292 3597
rect 2146 3552 2147 3599
rect 2376 3598 2377 3797
rect 2184 3600 2185 3797
rect 2282 3552 2283 3601
rect 2087 3602 2088 3797
rect 2283 3602 2284 3797
rect 2190 3604 2191 3797
rect 2228 3552 2229 3605
rect 2192 3552 2193 3607
rect 2435 3552 2436 3607
rect 2196 3608 2197 3797
rect 2267 3552 2268 3609
rect 2205 3610 2206 3797
rect 2336 3552 2337 3611
rect 2207 3552 2208 3613
rect 2367 3612 2368 3797
rect 2165 3552 2166 3615
rect 2208 3614 2209 3797
rect 2217 3614 2218 3797
rect 2355 3614 2356 3797
rect 2223 3616 2224 3797
rect 2258 3552 2259 3617
rect 2229 3618 2230 3797
rect 2339 3552 2340 3619
rect 2235 3620 2236 3797
rect 2369 3552 2370 3621
rect 2238 3622 2239 3797
rect 2372 3552 2373 3623
rect 2177 3552 2178 3625
rect 2373 3624 2374 3797
rect 2178 3626 2179 3797
rect 2450 3552 2451 3627
rect 2241 3628 2242 3797
rect 2432 3552 2433 3629
rect 2243 3552 2244 3631
rect 2453 3552 2454 3631
rect 2250 3632 2251 3797
rect 2387 3552 2388 3633
rect 2256 3634 2257 3797
rect 2309 3552 2310 3635
rect 2261 3552 2262 3637
rect 2292 3636 2293 3797
rect 2262 3638 2263 3797
rect 2405 3552 2406 3639
rect 2268 3640 2269 3797
rect 2399 3552 2400 3641
rect 2279 3552 2280 3643
rect 2454 3642 2455 3797
rect 2285 3552 2286 3645
rect 2343 3644 2344 3797
rect 2120 3552 2121 3647
rect 2286 3646 2287 3797
rect 2120 3648 2121 3797
rect 2301 3648 2302 3797
rect 2295 3650 2296 3797
rect 2297 3552 2298 3651
rect 2307 3650 2308 3797
rect 2447 3552 2448 3651
rect 2312 3552 2313 3653
rect 2319 3652 2320 3797
rect 2303 3552 2304 3655
rect 2313 3654 2314 3797
rect 2324 3552 2325 3655
rect 2535 3654 2536 3797
rect 2330 3552 2331 3657
rect 2523 3656 2524 3797
rect 2331 3658 2332 3797
rect 2396 3552 2397 3659
rect 2334 3660 2335 3797
rect 2393 3552 2394 3661
rect 2337 3662 2338 3797
rect 2471 3552 2472 3663
rect 2349 3664 2350 3797
rect 2477 3552 2478 3665
rect 2351 3552 2352 3667
rect 2457 3666 2458 3797
rect 2357 3552 2358 3669
rect 2541 3668 2542 3797
rect 2361 3670 2362 3797
rect 2411 3552 2412 3671
rect 2379 3672 2380 3797
rect 2667 3552 2668 3673
rect 2385 3674 2386 3797
rect 2519 3552 2520 3675
rect 2397 3676 2398 3797
rect 2537 3552 2538 3677
rect 2403 3678 2404 3797
rect 2423 3552 2424 3679
rect 2424 3680 2425 3797
rect 2528 3552 2529 3681
rect 2439 3682 2440 3797
rect 2495 3552 2496 3683
rect 2174 3552 2175 3685
rect 2496 3684 2497 3797
rect 2175 3686 2176 3797
rect 2451 3686 2452 3797
rect 2463 3686 2464 3797
rect 2737 3552 2738 3687
rect 2465 3552 2466 3689
rect 2585 3552 2586 3689
rect 2474 3552 2475 3691
rect 2559 3690 2560 3797
rect 2487 3692 2488 3797
rect 2612 3552 2613 3693
rect 2499 3694 2500 3797
rect 2603 3552 2604 3695
rect 2501 3552 2502 3697
rect 2598 3696 2599 3797
rect 2502 3698 2503 3797
rect 2606 3552 2607 3699
rect 2504 3552 2505 3701
rect 2601 3700 2602 3797
rect 2363 3552 2364 3703
rect 2505 3702 2506 3797
rect 2507 3552 2508 3703
rect 2511 3702 2512 3797
rect 2529 3702 2530 3797
rect 2670 3702 2671 3797
rect 2543 3552 2544 3705
rect 2689 3704 2690 3797
rect 2546 3552 2547 3707
rect 2589 3706 2590 3797
rect 2549 3552 2550 3709
rect 2776 3552 2777 3709
rect 2553 3710 2554 3797
rect 2752 3552 2753 3711
rect 2555 3552 2556 3713
rect 2686 3712 2687 3797
rect 2571 3714 2572 3797
rect 2591 3552 2592 3715
rect 2583 3716 2584 3797
rect 2633 3552 2634 3717
rect 2586 3718 2587 3797
rect 2692 3718 2693 3797
rect 2604 3720 2605 3797
rect 2639 3552 2640 3721
rect 2627 3552 2628 3723
rect 2661 3722 2662 3797
rect 2628 3724 2629 3797
rect 2664 3552 2665 3725
rect 2630 3552 2631 3727
rect 2778 3726 2779 3797
rect 2631 3728 2632 3797
rect 2657 3552 2658 3729
rect 2636 3552 2637 3731
rect 2818 3552 2819 3731
rect 2427 3732 2428 3797
rect 2818 3732 2819 3797
rect 2640 3734 2641 3797
rect 2645 3552 2646 3735
rect 2489 3552 2490 3737
rect 2646 3736 2647 3797
rect 2441 3552 2442 3739
rect 2490 3738 2491 3797
rect 2643 3738 2644 3797
rect 2648 3552 2649 3739
rect 2492 3552 2493 3741
rect 2649 3740 2650 3797
rect 2264 3552 2265 3743
rect 2493 3742 2494 3797
rect 2265 3744 2266 3797
rect 2408 3552 2409 3745
rect 2409 3746 2410 3797
rect 2752 3746 2753 3797
rect 2658 3748 2659 3797
rect 2808 3748 2809 3797
rect 2673 3750 2674 3797
rect 2716 3750 2717 3797
rect 2677 3552 2678 3753
rect 2683 3752 2684 3797
rect 2609 3552 2610 3755
rect 2677 3754 2678 3797
rect 2610 3756 2611 3797
rect 2734 3552 2735 3757
rect 2680 3552 2681 3759
rect 2801 3552 2802 3759
rect 2695 3552 2696 3761
rect 2758 3760 2759 3797
rect 2701 3552 2702 3763
rect 2815 3552 2816 3763
rect 2707 3552 2708 3765
rect 2811 3552 2812 3765
rect 2707 3766 2708 3797
rect 2773 3552 2774 3767
rect 2710 3768 2711 3797
rect 2713 3552 2714 3769
rect 2713 3770 2714 3797
rect 2728 3552 2729 3771
rect 2722 3772 2723 3797
rect 2725 3552 2726 3773
rect 2731 3772 2732 3797
rect 2731 3552 2732 3773
rect 2734 3772 2735 3797
rect 2790 3552 2791 3773
rect 2737 3774 2738 3797
rect 2746 3552 2747 3775
rect 2743 3552 2744 3777
rect 2787 3552 2788 3777
rect 2421 3778 2422 3797
rect 2787 3778 2788 3797
rect 2743 3780 2744 3797
rect 2767 3552 2768 3781
rect 2481 3782 2482 3797
rect 2768 3782 2769 3797
rect 2746 3784 2747 3797
rect 2770 3552 2771 3785
rect 2755 3786 2756 3797
rect 2761 3552 2762 3787
rect 2567 3552 2568 3789
rect 2761 3788 2762 3797
rect 2764 3552 2765 3789
rect 2783 3552 2784 3789
rect 2680 3790 2681 3797
rect 2764 3790 2765 3797
rect 2749 3552 2750 3793
rect 2784 3792 2785 3797
rect 2525 3552 2526 3795
rect 2749 3794 2750 3797
rect 2781 3794 2782 3797
rect 2811 3794 2812 3797
rect 2815 3794 2816 3797
rect 2832 3552 2833 3795
rect 2038 3801 2039 3804
rect 2123 3801 2124 3804
rect 2042 3801 2043 3806
rect 2126 3801 2127 3806
rect 2059 3801 2060 3808
rect 2235 3801 2236 3808
rect 2068 3809 2069 4022
rect 2225 3809 2226 4022
rect 2077 3801 2078 3812
rect 2229 3801 2230 3812
rect 2087 3801 2088 3814
rect 2250 3801 2251 3814
rect 2089 3815 2090 4022
rect 2216 3815 2217 4022
rect 2091 3801 2092 3818
rect 2112 3817 2113 4022
rect 2100 3819 2101 4022
rect 2283 3801 2284 3820
rect 2124 3821 2125 4022
rect 2339 3821 2340 4022
rect 2129 3801 2130 3824
rect 2241 3801 2242 3824
rect 2072 3825 2073 4022
rect 2240 3825 2241 4022
rect 2132 3801 2133 3828
rect 2258 3827 2259 4022
rect 2139 3801 2140 3830
rect 2313 3801 2314 3830
rect 2120 3801 2121 3832
rect 2312 3831 2313 4022
rect 2141 3833 2142 4022
rect 2355 3801 2356 3834
rect 2172 3801 2173 3836
rect 2598 3801 2599 3836
rect 2175 3801 2176 3838
rect 2334 3801 2335 3838
rect 2174 3839 2175 4022
rect 2178 3801 2179 3840
rect 2180 3839 2181 4022
rect 2238 3801 2239 3840
rect 2184 3801 2185 3842
rect 2337 3801 2338 3842
rect 2187 3801 2188 3844
rect 2262 3801 2263 3844
rect 2192 3845 2193 4022
rect 2496 3801 2497 3846
rect 2196 3801 2197 3848
rect 2234 3847 2235 4022
rect 2075 3849 2076 4022
rect 2195 3849 2196 4022
rect 2199 3801 2200 3850
rect 2210 3849 2211 4022
rect 2198 3851 2199 4022
rect 2208 3801 2209 3852
rect 2205 3801 2206 3854
rect 2237 3853 2238 4022
rect 2190 3801 2191 3856
rect 2204 3855 2205 4022
rect 2214 3801 2215 3856
rect 2529 3801 2530 3856
rect 2228 3857 2229 4022
rect 2454 3801 2455 3858
rect 2246 3859 2247 4022
rect 2373 3801 2374 3860
rect 2268 3801 2269 3862
rect 2297 3861 2298 4022
rect 2080 3801 2081 3864
rect 2267 3863 2268 4022
rect 2079 3865 2080 4022
rect 2220 3801 2221 3866
rect 2271 3801 2272 3866
rect 2559 3801 2560 3866
rect 2265 3801 2266 3868
rect 2270 3867 2271 4022
rect 2274 3801 2275 3868
rect 2516 3867 2517 4022
rect 2273 3869 2274 4022
rect 2343 3801 2344 3870
rect 2277 3801 2278 3872
rect 2309 3871 2310 4022
rect 2279 3873 2280 4022
rect 2286 3801 2287 3874
rect 2256 3801 2257 3876
rect 2285 3875 2286 4022
rect 2289 3801 2290 3876
rect 2315 3875 2316 4022
rect 2295 3801 2296 3878
rect 2303 3877 2304 4022
rect 2253 3801 2254 3880
rect 2294 3879 2295 4022
rect 2223 3801 2224 3882
rect 2252 3881 2253 4022
rect 2301 3801 2302 3882
rect 2345 3881 2346 4022
rect 2094 3801 2095 3884
rect 2300 3883 2301 4022
rect 2093 3885 2094 4022
rect 2222 3885 2223 4022
rect 2307 3801 2308 3886
rect 2333 3885 2334 4022
rect 2319 3801 2320 3888
rect 2321 3887 2322 4022
rect 2292 3801 2293 3890
rect 2318 3889 2319 4022
rect 2117 3801 2118 3892
rect 2291 3891 2292 4022
rect 2327 3891 2328 4022
rect 2349 3801 2350 3892
rect 2348 3893 2349 4022
rect 2376 3801 2377 3894
rect 2351 3895 2352 4022
rect 2535 3801 2536 3896
rect 2354 3897 2355 4022
rect 2493 3801 2494 3898
rect 2357 3899 2358 4022
rect 2451 3801 2452 3900
rect 2360 3901 2361 4022
rect 2361 3801 2362 3902
rect 2366 3901 2367 4022
rect 2367 3801 2368 3902
rect 2372 3901 2373 4022
rect 2457 3801 2458 3902
rect 2385 3801 2386 3904
rect 2727 3903 2728 4022
rect 2390 3905 2391 4022
rect 2764 3801 2765 3906
rect 2397 3801 2398 3908
rect 2815 3801 2816 3908
rect 2396 3909 2397 4022
rect 2403 3801 2404 3910
rect 2379 3801 2380 3912
rect 2402 3911 2403 4022
rect 2409 3801 2410 3912
rect 2617 3911 2618 4022
rect 2414 3913 2415 4022
rect 2601 3801 2602 3914
rect 2417 3915 2418 4022
rect 2505 3801 2506 3916
rect 2424 3801 2425 3918
rect 2749 3801 2750 3918
rect 2429 3919 2430 4022
rect 2752 3801 2753 3920
rect 2432 3921 2433 4022
rect 2686 3801 2687 3922
rect 2427 3801 2428 3924
rect 2686 3923 2687 4022
rect 2421 3801 2422 3926
rect 2426 3925 2427 4022
rect 2439 3801 2440 3926
rect 2771 3801 2772 3926
rect 2438 3927 2439 4022
rect 2463 3801 2464 3928
rect 2456 3929 2457 4022
rect 2490 3801 2491 3930
rect 2462 3931 2463 4022
rect 2655 3801 2656 3932
rect 2474 3933 2475 4022
rect 2502 3801 2503 3934
rect 2492 3935 2493 4022
rect 2511 3801 2512 3936
rect 2499 3801 2500 3938
rect 2513 3937 2514 4022
rect 2481 3801 2482 3940
rect 2498 3939 2499 4022
rect 2480 3941 2481 4022
rect 2523 3801 2524 3942
rect 2510 3943 2511 4022
rect 2801 3801 2802 3944
rect 2528 3945 2529 4022
rect 2628 3801 2629 3946
rect 2531 3947 2532 4022
rect 2631 3801 2632 3948
rect 2534 3949 2535 4022
rect 2586 3801 2587 3950
rect 2537 3951 2538 4022
rect 2571 3801 2572 3952
rect 2487 3801 2488 3954
rect 2570 3953 2571 4022
rect 2486 3955 2487 4022
rect 2541 3801 2542 3956
rect 2543 3955 2544 4022
rect 2640 3801 2641 3956
rect 2546 3957 2547 4022
rect 2601 3957 2602 4022
rect 2549 3959 2550 4022
rect 2553 3801 2554 3960
rect 2567 3959 2568 4022
rect 2677 3801 2678 3960
rect 2573 3961 2574 4022
rect 2604 3801 2605 3962
rect 2583 3801 2584 3964
rect 2692 3963 2693 4022
rect 2585 3965 2586 4022
rect 2646 3801 2647 3966
rect 2589 3801 2590 3968
rect 2689 3801 2690 3968
rect 2588 3969 2589 4022
rect 2649 3801 2650 3970
rect 2604 3971 2605 4022
rect 2811 3801 2812 3972
rect 2610 3801 2611 3974
rect 2668 3973 2669 4022
rect 2610 3975 2611 4022
rect 2734 3801 2735 3976
rect 2331 3801 2332 3978
rect 2734 3977 2735 4022
rect 2623 3979 2624 4022
rect 2658 3801 2659 3980
rect 2626 3981 2627 4022
rect 2661 3801 2662 3982
rect 2643 3801 2644 3984
rect 2673 3801 2674 3984
rect 2647 3985 2648 4022
rect 2707 3801 2708 3986
rect 2650 3987 2651 4022
rect 2710 3801 2711 3988
rect 2653 3989 2654 4022
rect 2720 3989 2721 4022
rect 2665 3991 2666 4022
rect 2731 3801 2732 3992
rect 2450 3993 2451 4022
rect 2730 3993 2731 4022
rect 2683 3801 2684 3996
rect 2808 3801 2809 3996
rect 2683 3997 2684 4022
rect 2743 3801 2744 3998
rect 2689 3999 2690 4022
rect 2794 3801 2795 4000
rect 2695 4001 2696 4022
rect 2775 3801 2776 4002
rect 2701 4003 2702 4022
rect 2755 3801 2756 4004
rect 2704 4005 2705 4022
rect 2758 3801 2759 4006
rect 2707 4007 2708 4022
rect 2713 3801 2714 4008
rect 2710 4009 2711 4022
rect 2716 3801 2717 4010
rect 2635 4011 2636 4022
rect 2716 4011 2717 4022
rect 2737 4011 2738 4022
rect 2763 4011 2764 4022
rect 2740 4013 2741 4022
rect 2781 3801 2782 4014
rect 2743 4015 2744 4022
rect 2784 3801 2785 4016
rect 2746 3801 2747 4018
rect 2787 3801 2788 4018
rect 2698 4019 2699 4022
rect 2746 4019 2747 4022
rect 2056 4026 2057 4029
rect 2267 4026 2268 4029
rect 2082 4026 2083 4031
rect 2285 4026 2286 4031
rect 2083 4032 2084 4241
rect 2291 4026 2292 4033
rect 2087 4034 2088 4241
rect 2163 4034 2164 4241
rect 2089 4026 2090 4037
rect 2300 4026 2301 4037
rect 2097 4038 2098 4241
rect 2127 4026 2128 4039
rect 2100 4026 2101 4041
rect 2385 4040 2386 4241
rect 2103 4026 2104 4043
rect 2318 4026 2319 4043
rect 2104 4044 2105 4241
rect 2312 4026 2313 4045
rect 2079 4026 2080 4047
rect 2313 4046 2314 4241
rect 2080 4048 2081 4241
rect 2094 4048 2095 4241
rect 2112 4026 2113 4049
rect 2370 4048 2371 4241
rect 2119 4050 2120 4241
rect 2315 4026 2316 4051
rect 2122 4052 2123 4241
rect 2343 4052 2344 4241
rect 2129 4054 2130 4241
rect 2222 4026 2223 4055
rect 2131 4026 2132 4057
rect 2303 4026 2304 4057
rect 2133 4058 2134 4241
rect 2246 4026 2247 4059
rect 2138 4026 2139 4061
rect 2339 4026 2340 4061
rect 2141 4026 2142 4063
rect 2345 4026 2346 4063
rect 2148 4064 2149 4241
rect 2340 4064 2341 4241
rect 2157 4066 2158 4241
rect 2193 4066 2194 4241
rect 2174 4026 2175 4069
rect 2175 4068 2176 4241
rect 2180 4026 2181 4069
rect 2181 4068 2182 4241
rect 2189 4026 2190 4069
rect 2265 4068 2266 4241
rect 2068 4026 2069 4071
rect 2190 4070 2191 4241
rect 2198 4026 2199 4071
rect 2202 4070 2203 4241
rect 2195 4026 2196 4073
rect 2199 4072 2200 4241
rect 2204 4026 2205 4073
rect 2208 4072 2209 4241
rect 2210 4026 2211 4073
rect 2214 4072 2215 4241
rect 2216 4026 2217 4073
rect 2220 4072 2221 4241
rect 2225 4026 2226 4073
rect 2388 4072 2389 4241
rect 2226 4074 2227 4241
rect 2546 4026 2547 4075
rect 2228 4026 2229 4077
rect 2304 4076 2305 4241
rect 2231 4026 2232 4079
rect 2357 4026 2358 4079
rect 2234 4026 2235 4081
rect 2268 4080 2269 4241
rect 2237 4026 2238 4083
rect 2301 4082 2302 4241
rect 2240 4026 2241 4085
rect 2244 4084 2245 4241
rect 2252 4026 2253 4085
rect 2346 4084 2347 4241
rect 2256 4086 2257 4241
rect 2421 4086 2422 4241
rect 2258 4026 2259 4089
rect 2406 4088 2407 4241
rect 2261 4026 2262 4091
rect 2480 4026 2481 4091
rect 2262 4092 2263 4241
rect 2354 4026 2355 4093
rect 2076 4094 2077 4241
rect 2355 4094 2356 4241
rect 2270 4026 2271 4097
rect 2358 4096 2359 4241
rect 2271 4098 2272 4241
rect 2273 4026 2274 4099
rect 2277 4098 2278 4241
rect 2321 4026 2322 4099
rect 2279 4026 2280 4101
rect 2376 4100 2377 4241
rect 2294 4026 2295 4103
rect 2316 4102 2317 4241
rect 2295 4104 2296 4241
rect 2486 4026 2487 4105
rect 2319 4106 2320 4241
rect 2372 4026 2373 4107
rect 2309 4026 2310 4109
rect 2373 4108 2374 4241
rect 2325 4110 2326 4241
rect 2516 4026 2517 4111
rect 2330 4026 2331 4113
rect 2583 4112 2584 4241
rect 2331 4114 2332 4241
rect 2417 4026 2418 4115
rect 2337 4116 2338 4241
rect 2351 4026 2352 4117
rect 2348 4026 2349 4119
rect 2418 4118 2419 4241
rect 2360 4026 2361 4121
rect 2379 4120 2380 4241
rect 2366 4026 2367 4123
rect 2594 4026 2595 4123
rect 2297 4026 2298 4125
rect 2367 4124 2368 4241
rect 2390 4026 2391 4125
rect 2478 4124 2479 4241
rect 2391 4126 2392 4241
rect 2528 4026 2529 4127
rect 2394 4128 2395 4241
rect 2531 4026 2532 4129
rect 2396 4026 2397 4131
rect 2409 4130 2410 4241
rect 2402 4026 2403 4133
rect 2490 4132 2491 4241
rect 2126 4134 2127 4241
rect 2403 4134 2404 4241
rect 2429 4026 2430 4135
rect 2502 4134 2503 4241
rect 2438 4026 2439 4137
rect 2610 4026 2611 4137
rect 2450 4026 2451 4139
rect 2520 4138 2521 4241
rect 2451 4140 2452 4241
rect 2543 4026 2544 4141
rect 2454 4142 2455 4241
rect 2534 4026 2535 4143
rect 2460 4144 2461 4241
rect 2567 4026 2568 4145
rect 2466 4146 2467 4241
rect 2585 4026 2586 4147
rect 2414 4026 2415 4149
rect 2586 4148 2587 4241
rect 2333 4026 2334 4151
rect 2415 4150 2416 4241
rect 2469 4150 2470 4241
rect 2588 4026 2589 4151
rect 2492 4026 2493 4153
rect 2718 4152 2719 4241
rect 2508 4154 2509 4241
rect 2730 4026 2731 4155
rect 2505 4156 2506 4241
rect 2731 4156 2732 4241
rect 2510 4026 2511 4159
rect 2568 4158 2569 4241
rect 2513 4026 2514 4161
rect 2773 4160 2774 4241
rect 2432 4026 2433 4163
rect 2514 4162 2515 4241
rect 2433 4164 2434 4241
rect 2637 4164 2638 4241
rect 2537 4026 2538 4167
rect 2544 4166 2545 4241
rect 2462 4026 2463 4169
rect 2538 4168 2539 4241
rect 2463 4170 2464 4241
rect 2570 4026 2571 4171
rect 2474 4026 2475 4173
rect 2571 4172 2572 4241
rect 2549 4026 2550 4175
rect 2595 4174 2596 4241
rect 2550 4176 2551 4241
rect 2573 4026 2574 4177
rect 2498 4026 2499 4179
rect 2574 4178 2575 4241
rect 2426 4026 2427 4181
rect 2499 4180 2500 4241
rect 2427 4182 2428 4241
rect 2456 4026 2457 4183
rect 2457 4184 2458 4241
rect 2617 4026 2618 4185
rect 2562 4186 2563 4241
rect 2668 4026 2669 4187
rect 2580 4188 2581 4241
rect 2692 4026 2693 4189
rect 2598 4026 2599 4191
rect 2613 4026 2614 4191
rect 2238 4192 2239 4241
rect 2613 4192 2614 4241
rect 2601 4194 2602 4241
rect 2781 4026 2782 4195
rect 2623 4026 2624 4197
rect 2755 4196 2756 4241
rect 2445 4198 2446 4241
rect 2622 4198 2623 4241
rect 2643 4198 2644 4241
rect 2753 4026 2754 4199
rect 2647 4026 2648 4201
rect 2673 4200 2674 4241
rect 2646 4202 2647 4241
rect 2767 4026 2768 4203
rect 2650 4026 2651 4205
rect 2727 4204 2728 4241
rect 2653 4026 2654 4207
rect 2713 4026 2714 4207
rect 2652 4208 2653 4241
rect 2676 4208 2677 4241
rect 2655 4210 2656 4241
rect 2724 4210 2725 4241
rect 2679 4212 2680 4241
rect 2743 4026 2744 4213
rect 2689 4026 2690 4215
rect 2760 4026 2761 4215
rect 2691 4216 2692 4241
rect 2707 4026 2708 4217
rect 2695 4026 2696 4219
rect 2749 4026 2750 4219
rect 2526 4220 2527 4241
rect 2748 4220 2749 4241
rect 2635 4026 2636 4223
rect 2694 4222 2695 4241
rect 2701 4026 2702 4223
rect 2721 4222 2722 4241
rect 2686 4026 2687 4225
rect 2700 4224 2701 4241
rect 2704 4026 2705 4225
rect 2777 4026 2778 4225
rect 2665 4026 2666 4227
rect 2703 4226 2704 4241
rect 2710 4026 2711 4227
rect 2716 4026 2717 4227
rect 2484 4228 2485 4241
rect 2715 4228 2716 4241
rect 2698 4026 2699 4231
rect 2709 4230 2710 4241
rect 2683 4026 2684 4233
rect 2697 4232 2698 4241
rect 2604 4026 2605 4235
rect 2682 4234 2683 4241
rect 2712 4234 2713 4241
rect 2734 4026 2735 4235
rect 2626 4026 2627 4237
rect 2734 4236 2735 4241
rect 2740 4026 2741 4237
rect 2780 4236 2781 4241
rect 2706 4238 2707 4241
rect 2741 4238 2742 4241
rect 2044 4247 2045 4464
rect 2190 4245 2191 4248
rect 2059 4245 2060 4250
rect 2087 4245 2088 4250
rect 2063 4251 2064 4464
rect 2268 4245 2269 4252
rect 2067 4253 2068 4464
rect 2199 4245 2200 4254
rect 2069 4245 2070 4256
rect 2206 4255 2207 4464
rect 2074 4257 2075 4464
rect 2233 4257 2234 4464
rect 2076 4245 2077 4260
rect 2083 4245 2084 4260
rect 2084 4261 2085 4464
rect 2293 4261 2294 4464
rect 2095 4263 2096 4464
rect 2365 4263 2366 4464
rect 2097 4245 2098 4266
rect 2388 4245 2389 4266
rect 2098 4267 2099 4464
rect 2403 4245 2404 4268
rect 2104 4245 2105 4270
rect 2311 4269 2312 4464
rect 2107 4271 2108 4464
rect 2116 4271 2117 4464
rect 2113 4273 2114 4464
rect 2373 4245 2374 4274
rect 2129 4245 2130 4276
rect 2353 4275 2354 4464
rect 2133 4245 2134 4278
rect 2415 4245 2416 4278
rect 2135 4279 2136 4464
rect 2275 4279 2276 4464
rect 2142 4281 2143 4464
rect 2202 4245 2203 4282
rect 2070 4283 2071 4464
rect 2203 4283 2204 4464
rect 2148 4245 2149 4286
rect 2271 4245 2272 4286
rect 2157 4287 2158 4464
rect 2316 4245 2317 4288
rect 2160 4245 2161 4290
rect 2265 4245 2266 4290
rect 2163 4245 2164 4292
rect 2317 4291 2318 4464
rect 2166 4293 2167 4464
rect 2284 4293 2285 4464
rect 2175 4245 2176 4296
rect 2176 4295 2177 4464
rect 2181 4245 2182 4296
rect 2188 4295 2189 4464
rect 2193 4245 2194 4296
rect 2226 4245 2227 4296
rect 2214 4245 2215 4298
rect 2227 4297 2228 4464
rect 2215 4299 2216 4464
rect 2220 4245 2221 4300
rect 2208 4245 2209 4302
rect 2221 4301 2222 4464
rect 2238 4245 2239 4302
rect 2325 4245 2326 4302
rect 2244 4245 2245 4304
rect 2254 4303 2255 4464
rect 2245 4305 2246 4464
rect 2301 4245 2302 4306
rect 2248 4307 2249 4464
rect 2626 4307 2627 4464
rect 2256 4245 2257 4310
rect 2370 4245 2371 4310
rect 2241 4245 2242 4312
rect 2371 4311 2372 4464
rect 2119 4245 2120 4314
rect 2242 4313 2243 4464
rect 2272 4313 2273 4464
rect 2406 4245 2407 4314
rect 2290 4315 2291 4464
rect 2313 4245 2314 4316
rect 2299 4317 2300 4464
rect 2418 4245 2419 4318
rect 2302 4319 2303 4464
rect 2355 4245 2356 4320
rect 2308 4321 2309 4464
rect 2376 4245 2377 4322
rect 2314 4323 2315 4464
rect 2367 4245 2368 4324
rect 2326 4325 2327 4464
rect 2385 4245 2386 4326
rect 2323 4327 2324 4464
rect 2386 4327 2387 4464
rect 2335 4329 2336 4464
rect 2343 4245 2344 4330
rect 2340 4245 2341 4332
rect 2356 4331 2357 4464
rect 2304 4245 2305 4334
rect 2341 4333 2342 4464
rect 2305 4335 2306 4464
rect 2358 4245 2359 4336
rect 2319 4245 2320 4338
rect 2359 4337 2360 4464
rect 2262 4245 2263 4340
rect 2320 4339 2321 4464
rect 2368 4339 2369 4464
rect 2718 4245 2719 4340
rect 2377 4341 2378 4464
rect 2445 4245 2446 4342
rect 2389 4343 2390 4464
rect 2409 4245 2410 4344
rect 2401 4345 2402 4464
rect 2586 4245 2587 4346
rect 2413 4347 2414 4464
rect 2478 4245 2479 4348
rect 2419 4349 2420 4464
rect 2484 4245 2485 4350
rect 2425 4351 2426 4464
rect 2490 4245 2491 4352
rect 2427 4245 2428 4354
rect 2637 4245 2638 4354
rect 2433 4245 2434 4356
rect 2437 4355 2438 4464
rect 2449 4355 2450 4464
rect 2514 4245 2515 4356
rect 2451 4245 2452 4358
rect 2530 4357 2531 4464
rect 2457 4245 2458 4360
rect 2619 4245 2620 4360
rect 2229 4245 2230 4362
rect 2620 4361 2621 4464
rect 2463 4245 2464 4364
rect 2640 4245 2641 4364
rect 2466 4245 2467 4366
rect 2617 4365 2618 4464
rect 2469 4245 2470 4368
rect 2518 4367 2519 4464
rect 2491 4369 2492 4464
rect 2796 4369 2797 4464
rect 2497 4371 2498 4464
rect 2684 4371 2685 4464
rect 2508 4245 2509 4374
rect 2512 4373 2513 4464
rect 2509 4375 2510 4464
rect 2571 4245 2572 4376
rect 2520 4245 2521 4378
rect 2745 4245 2746 4378
rect 2421 4245 2422 4380
rect 2745 4379 2746 4464
rect 2533 4381 2534 4464
rect 2574 4245 2575 4382
rect 2542 4383 2543 4464
rect 2652 4245 2653 4384
rect 2550 4245 2551 4386
rect 2605 4385 2606 4464
rect 2544 4245 2545 4388
rect 2551 4387 2552 4464
rect 2545 4389 2546 4464
rect 2649 4245 2650 4390
rect 2460 4245 2461 4392
rect 2650 4391 2651 4464
rect 2295 4245 2296 4394
rect 2461 4393 2462 4464
rect 2277 4245 2278 4396
rect 2296 4395 2297 4464
rect 2562 4245 2563 4396
rect 2599 4395 2600 4464
rect 2563 4397 2564 4464
rect 2595 4245 2596 4398
rect 2568 4245 2569 4400
rect 2773 4245 2774 4400
rect 2569 4401 2570 4464
rect 2580 4245 2581 4402
rect 2394 4245 2395 4404
rect 2581 4403 2582 4464
rect 2331 4245 2332 4406
rect 2395 4405 2396 4464
rect 2575 4405 2576 4464
rect 2601 4245 2602 4406
rect 2587 4407 2588 4464
rect 2687 4407 2688 4464
rect 2593 4409 2594 4464
rect 2738 4409 2739 4464
rect 2610 4245 2611 4412
rect 2622 4245 2623 4412
rect 2583 4245 2584 4414
rect 2623 4413 2624 4464
rect 2391 4245 2392 4416
rect 2584 4415 2585 4464
rect 2613 4245 2614 4416
rect 2668 4415 2669 4464
rect 2646 4245 2647 4418
rect 2755 4245 2756 4418
rect 2647 4419 2648 4464
rect 2734 4245 2735 4420
rect 2655 4245 2656 4422
rect 2665 4421 2666 4464
rect 2673 4245 2674 4422
rect 2727 4245 2728 4422
rect 2676 4245 2677 4424
rect 2724 4245 2725 4424
rect 2526 4245 2527 4426
rect 2723 4425 2724 4464
rect 2694 4245 2695 4428
rect 2741 4245 2742 4428
rect 2499 4245 2500 4430
rect 2742 4429 2743 4464
rect 2500 4431 2501 4464
rect 2505 4245 2506 4432
rect 2682 4245 2683 4432
rect 2693 4431 2694 4464
rect 2703 4245 2704 4432
rect 2726 4431 2727 4464
rect 2702 4433 2703 4464
rect 2785 4433 2786 4464
rect 2706 4245 2707 4436
rect 2729 4435 2730 4464
rect 2643 4245 2644 4438
rect 2705 4437 2706 4464
rect 2712 4245 2713 4438
rect 2756 4437 2757 4464
rect 2700 4245 2701 4440
rect 2711 4439 2712 4464
rect 2699 4441 2700 4464
rect 2715 4245 2716 4442
rect 2278 4443 2279 4464
rect 2714 4443 2715 4464
rect 2759 4443 2760 4464
rect 2759 4245 2760 4444
rect 2762 4245 2763 4444
rect 2766 4245 2767 4444
rect 2731 4245 2732 4446
rect 2763 4445 2764 4464
rect 2721 4245 2722 4448
rect 2732 4447 2733 4464
rect 2709 4245 2710 4450
rect 2720 4449 2721 4464
rect 2697 4245 2698 4452
rect 2708 4451 2709 4464
rect 2691 4245 2692 4454
rect 2696 4453 2697 4464
rect 2679 4245 2680 4456
rect 2690 4455 2691 4464
rect 2379 4245 2380 4458
rect 2680 4457 2681 4464
rect 2769 4245 2770 4458
rect 2787 4245 2788 4458
rect 2769 4459 2770 4464
rect 2776 4245 2777 4460
rect 2772 4461 2773 4464
rect 2782 4461 2783 4464
rect 2053 4470 2054 4705
rect 2060 4470 2061 4705
rect 2056 4468 2057 4473
rect 2188 4468 2189 4473
rect 2063 4474 2064 4705
rect 2199 4474 2200 4705
rect 2070 4468 2071 4477
rect 2206 4468 2207 4477
rect 2074 4468 2075 4479
rect 2227 4468 2228 4479
rect 2074 4480 2075 4705
rect 2299 4468 2300 4481
rect 2077 4468 2078 4483
rect 2221 4468 2222 4483
rect 2081 4484 2082 4705
rect 2193 4484 2194 4705
rect 2084 4468 2085 4487
rect 2272 4468 2273 4487
rect 2088 4468 2089 4489
rect 2311 4468 2312 4489
rect 2088 4490 2089 4705
rect 2205 4490 2206 4705
rect 2091 4492 2092 4705
rect 2335 4468 2336 4493
rect 2095 4468 2096 4495
rect 2302 4468 2303 4495
rect 2098 4468 2099 4497
rect 2254 4468 2255 4497
rect 2100 4498 2101 4705
rect 2107 4468 2108 4499
rect 2113 4468 2114 4499
rect 2135 4468 2136 4499
rect 2113 4500 2114 4705
rect 2317 4468 2318 4501
rect 2116 4468 2117 4503
rect 2296 4468 2297 4503
rect 2120 4468 2121 4505
rect 2308 4468 2309 4505
rect 2123 4468 2124 4507
rect 2256 4506 2257 4705
rect 2123 4508 2124 4705
rect 2290 4468 2291 4509
rect 2133 4510 2134 4705
rect 2157 4468 2158 4511
rect 2142 4512 2143 4705
rect 2176 4468 2177 4513
rect 2151 4514 2152 4705
rect 2356 4468 2357 4515
rect 2157 4516 2158 4705
rect 2203 4468 2204 4517
rect 2160 4518 2161 4705
rect 2245 4468 2246 4519
rect 2163 4468 2164 4521
rect 2353 4468 2354 4521
rect 2166 4468 2167 4523
rect 2251 4468 2252 4523
rect 2166 4524 2167 4705
rect 2233 4468 2234 4525
rect 2169 4526 2170 4705
rect 2305 4468 2306 4527
rect 2173 4468 2174 4529
rect 2284 4468 2285 4529
rect 2184 4530 2185 4705
rect 2275 4468 2276 4531
rect 2187 4532 2188 4705
rect 2371 4468 2372 4533
rect 2190 4534 2191 4705
rect 2271 4534 2272 4705
rect 2196 4536 2197 4705
rect 2293 4468 2294 4537
rect 2202 4538 2203 4705
rect 2338 4468 2339 4539
rect 2211 4540 2212 4705
rect 2283 4540 2284 4705
rect 2215 4468 2216 4543
rect 2220 4542 2221 4705
rect 2217 4544 2218 4705
rect 2314 4468 2315 4545
rect 2229 4546 2230 4705
rect 2278 4468 2279 4547
rect 2235 4548 2236 4705
rect 2326 4468 2327 4549
rect 2238 4550 2239 4705
rect 2320 4468 2321 4551
rect 2242 4468 2243 4553
rect 2629 4552 2630 4705
rect 2241 4554 2242 4705
rect 2323 4468 2324 4555
rect 2250 4556 2251 4705
rect 2684 4468 2685 4557
rect 2253 4558 2254 4705
rect 2347 4468 2348 4559
rect 2259 4560 2260 4705
rect 2341 4468 2342 4561
rect 2265 4562 2266 4705
rect 2365 4468 2366 4563
rect 2274 4564 2275 4705
rect 2368 4468 2369 4565
rect 2277 4566 2278 4705
rect 2359 4468 2360 4567
rect 2289 4568 2290 4705
rect 2386 4468 2387 4569
rect 2295 4570 2296 4705
rect 2389 4468 2390 4571
rect 2307 4572 2308 4705
rect 2749 4468 2750 4573
rect 2313 4574 2314 4705
rect 2687 4468 2688 4575
rect 2325 4576 2326 4705
rect 2413 4468 2414 4577
rect 2331 4578 2332 4705
rect 2680 4468 2681 4579
rect 2343 4580 2344 4705
rect 2699 4468 2700 4581
rect 2349 4582 2350 4705
rect 2461 4468 2462 4583
rect 2355 4584 2356 4705
rect 2437 4468 2438 4585
rect 2361 4586 2362 4705
rect 2449 4468 2450 4587
rect 2367 4588 2368 4705
rect 2455 4468 2456 4589
rect 2377 4468 2378 4591
rect 2383 4468 2384 4591
rect 2379 4592 2380 4705
rect 2711 4468 2712 4593
rect 2385 4594 2386 4705
rect 2745 4468 2746 4595
rect 2397 4596 2398 4705
rect 2723 4468 2724 4597
rect 2401 4468 2402 4599
rect 2641 4468 2642 4599
rect 2409 4600 2410 4705
rect 2491 4468 2492 4601
rect 2415 4602 2416 4705
rect 2503 4468 2504 4603
rect 2419 4468 2420 4605
rect 2608 4604 2609 4705
rect 2433 4606 2434 4705
rect 2497 4468 2498 4607
rect 2436 4608 2437 4705
rect 2500 4468 2501 4609
rect 2445 4610 2446 4705
rect 2581 4468 2582 4611
rect 2301 4612 2302 4705
rect 2580 4612 2581 4705
rect 2448 4614 2449 4705
rect 2584 4468 2585 4615
rect 2451 4616 2452 4705
rect 2533 4468 2534 4617
rect 2457 4618 2458 4705
rect 2530 4468 2531 4619
rect 2460 4620 2461 4705
rect 2679 4620 2680 4705
rect 2463 4622 2464 4705
rect 2539 4468 2540 4623
rect 2466 4624 2467 4705
rect 2542 4468 2543 4625
rect 2469 4626 2470 4705
rect 2551 4468 2552 4627
rect 2475 4628 2476 4705
rect 2545 4468 2546 4629
rect 2395 4468 2396 4631
rect 2544 4630 2545 4705
rect 2478 4632 2479 4705
rect 2512 4468 2513 4633
rect 2487 4634 2488 4705
rect 2617 4468 2618 4635
rect 2490 4636 2491 4705
rect 2620 4468 2621 4637
rect 2493 4638 2494 4705
rect 2563 4468 2564 4639
rect 2499 4640 2500 4705
rect 2569 4468 2570 4641
rect 2505 4642 2506 4705
rect 2593 4468 2594 4643
rect 2509 4468 2510 4645
rect 2538 4644 2539 4705
rect 2511 4646 2512 4705
rect 2715 4646 2716 4705
rect 2518 4468 2519 4649
rect 2805 4468 2806 4649
rect 2523 4650 2524 4705
rect 2599 4468 2600 4651
rect 2529 4652 2530 4705
rect 2759 4468 2760 4653
rect 2535 4654 2536 4705
rect 2789 4468 2790 4655
rect 2541 4656 2542 4705
rect 2547 4656 2548 4705
rect 2550 4656 2551 4705
rect 2623 4468 2624 4657
rect 2568 4658 2569 4705
rect 2650 4468 2651 4659
rect 2583 4660 2584 4705
rect 2665 4468 2666 4661
rect 2425 4468 2426 4663
rect 2665 4662 2666 4705
rect 2589 4664 2590 4705
rect 2729 4468 2730 4665
rect 2575 4468 2576 4667
rect 2729 4666 2730 4705
rect 2601 4668 2602 4705
rect 2647 4468 2648 4669
rect 2605 4468 2606 4671
rect 2735 4468 2736 4671
rect 2565 4672 2566 4705
rect 2604 4672 2605 4705
rect 2614 4672 2615 4705
rect 2690 4468 2691 4673
rect 2617 4674 2618 4705
rect 2693 4468 2694 4675
rect 2620 4676 2621 4705
rect 2696 4468 2697 4677
rect 2626 4468 2627 4679
rect 2644 4468 2645 4679
rect 2626 4680 2627 4705
rect 2720 4468 2721 4681
rect 2638 4682 2639 4705
rect 2799 4468 2800 4683
rect 2641 4684 2642 4705
rect 2708 4468 2709 4685
rect 2650 4686 2651 4705
rect 2732 4468 2733 4687
rect 2659 4688 2660 4705
rect 2785 4468 2786 4689
rect 2662 4690 2663 4705
rect 2726 4468 2727 4691
rect 2672 4692 2673 4705
rect 2705 4468 2706 4693
rect 2699 4694 2700 4705
rect 2769 4468 2770 4695
rect 2702 4468 2703 4697
rect 2766 4468 2767 4697
rect 2587 4468 2588 4699
rect 2702 4698 2703 4705
rect 2586 4700 2587 4705
rect 2668 4468 2669 4701
rect 2623 4702 2624 4705
rect 2668 4702 2669 4705
rect 2705 4702 2706 4705
rect 2772 4468 2773 4703
rect 2060 4709 2061 4712
rect 2225 4711 2226 4898
rect 2074 4709 2075 4714
rect 2191 4713 2192 4898
rect 2077 4715 2078 4898
rect 2188 4715 2189 4898
rect 2081 4709 2082 4718
rect 2166 4709 2167 4718
rect 2093 4719 2094 4898
rect 2100 4709 2101 4720
rect 2106 4709 2107 4720
rect 2235 4709 2236 4720
rect 2084 4709 2085 4722
rect 2105 4721 2106 4898
rect 2084 4723 2085 4898
rect 2133 4709 2134 4724
rect 2109 4709 2110 4726
rect 2234 4725 2235 4898
rect 2108 4727 2109 4898
rect 2125 4727 2126 4898
rect 2113 4709 2114 4730
rect 2141 4729 2142 4898
rect 2116 4709 2117 4732
rect 2157 4709 2158 4732
rect 2130 4709 2131 4734
rect 2289 4709 2290 4734
rect 2138 4735 2139 4898
rect 2207 4735 2208 4898
rect 2151 4709 2152 4738
rect 2295 4709 2296 4738
rect 2152 4739 2153 4898
rect 2184 4709 2185 4740
rect 2154 4709 2155 4742
rect 2466 4709 2467 4742
rect 2158 4743 2159 4898
rect 2169 4709 2170 4744
rect 2164 4745 2165 4898
rect 2241 4709 2242 4746
rect 2067 4709 2068 4748
rect 2240 4747 2241 4898
rect 2067 4749 2068 4898
rect 2182 4749 2183 4898
rect 2193 4709 2194 4750
rect 2243 4749 2244 4898
rect 2167 4751 2168 4898
rect 2194 4751 2195 4898
rect 2196 4709 2197 4752
rect 2246 4751 2247 4898
rect 2211 4709 2212 4754
rect 2620 4709 2621 4754
rect 2214 4709 2215 4756
rect 2650 4709 2651 4756
rect 2217 4709 2218 4758
rect 2261 4757 2262 4898
rect 2229 4709 2230 4760
rect 2288 4759 2289 4898
rect 2202 4709 2203 4762
rect 2228 4761 2229 4898
rect 2238 4709 2239 4762
rect 2285 4761 2286 4898
rect 2199 4709 2200 4764
rect 2237 4763 2238 4898
rect 2253 4709 2254 4764
rect 2303 4763 2304 4898
rect 2112 4765 2113 4898
rect 2252 4765 2253 4898
rect 2256 4709 2257 4766
rect 2297 4765 2298 4898
rect 2205 4709 2206 4768
rect 2255 4767 2256 4898
rect 2259 4709 2260 4768
rect 2580 4709 2581 4768
rect 2265 4709 2266 4770
rect 2318 4769 2319 4898
rect 2220 4709 2221 4772
rect 2264 4771 2265 4898
rect 2063 4773 2064 4898
rect 2219 4773 2220 4898
rect 2274 4709 2275 4774
rect 2321 4773 2322 4898
rect 2279 4775 2280 4898
rect 2643 4775 2644 4898
rect 2283 4709 2284 4778
rect 2550 4709 2551 4778
rect 2309 4779 2310 4898
rect 2490 4709 2491 4780
rect 2325 4709 2326 4782
rect 2647 4709 2648 4782
rect 2277 4709 2278 4784
rect 2324 4783 2325 4898
rect 2331 4709 2332 4784
rect 2372 4783 2373 4898
rect 2330 4785 2331 4898
rect 2349 4709 2350 4786
rect 2313 4709 2314 4788
rect 2348 4787 2349 4898
rect 2271 4709 2272 4790
rect 2312 4789 2313 4898
rect 2343 4709 2344 4790
rect 2715 4709 2716 4790
rect 2307 4709 2308 4792
rect 2342 4791 2343 4898
rect 2361 4709 2362 4792
rect 2390 4791 2391 4898
rect 2367 4709 2368 4794
rect 2402 4793 2403 4898
rect 2397 4709 2398 4796
rect 2712 4709 2713 4796
rect 2415 4709 2416 4798
rect 2429 4797 2430 4898
rect 2379 4709 2380 4800
rect 2414 4799 2415 4898
rect 2355 4709 2356 4802
rect 2378 4801 2379 4898
rect 2301 4709 2302 4804
rect 2354 4803 2355 4898
rect 2250 4709 2251 4806
rect 2300 4805 2301 4898
rect 2120 4709 2121 4808
rect 2249 4807 2250 4898
rect 2417 4807 2418 4898
rect 2445 4709 2446 4808
rect 2420 4809 2421 4898
rect 2448 4709 2449 4810
rect 2436 4709 2437 4812
rect 2438 4811 2439 4898
rect 2433 4709 2434 4814
rect 2435 4813 2436 4898
rect 2441 4813 2442 4898
rect 2457 4709 2458 4814
rect 2444 4815 2445 4898
rect 2460 4709 2461 4816
rect 2451 4709 2452 4818
rect 2465 4817 2466 4898
rect 2453 4819 2454 4898
rect 2478 4709 2479 4820
rect 2459 4821 2460 4898
rect 2463 4709 2464 4822
rect 2462 4823 2463 4898
rect 2577 4709 2578 4824
rect 2469 4709 2470 4826
rect 2477 4825 2478 4898
rect 2471 4827 2472 4898
rect 2568 4709 2569 4828
rect 2475 4709 2476 4830
rect 2483 4829 2484 4898
rect 2487 4709 2488 4830
rect 2507 4829 2508 4898
rect 2493 4709 2494 4832
rect 2576 4831 2577 4898
rect 2495 4833 2496 4898
rect 2668 4709 2669 4834
rect 2499 4709 2500 4836
rect 2519 4835 2520 4898
rect 2505 4709 2506 4838
rect 2513 4837 2514 4898
rect 2511 4709 2512 4840
rect 2531 4839 2532 4898
rect 2306 4841 2307 4898
rect 2510 4841 2511 4898
rect 2523 4709 2524 4842
rect 2708 4709 2709 4842
rect 2529 4709 2530 4844
rect 2693 4709 2694 4844
rect 2535 4709 2536 4846
rect 2555 4845 2556 4898
rect 2538 4709 2539 4848
rect 2558 4847 2559 4898
rect 2544 4709 2545 4850
rect 2612 4849 2613 4898
rect 2543 4851 2544 4898
rect 2547 4709 2548 4852
rect 2541 4709 2542 4854
rect 2546 4853 2547 4898
rect 2567 4853 2568 4898
rect 2629 4709 2630 4854
rect 2573 4855 2574 4898
rect 2617 4709 2618 4856
rect 2579 4857 2580 4898
rect 2604 4709 2605 4858
rect 2589 4709 2590 4860
rect 2594 4859 2595 4898
rect 2586 4709 2587 4862
rect 2588 4861 2589 4898
rect 2583 4709 2584 4864
rect 2585 4863 2586 4898
rect 2565 4709 2566 4866
rect 2582 4865 2583 4898
rect 2591 4865 2592 4898
rect 2708 4865 2709 4898
rect 2606 4867 2607 4898
rect 2623 4709 2624 4868
rect 2360 4869 2361 4898
rect 2624 4869 2625 4898
rect 2614 4709 2615 4872
rect 2729 4709 2730 4872
rect 2618 4873 2619 4898
rect 2696 4709 2697 4874
rect 2626 4709 2627 4876
rect 2652 4875 2653 4898
rect 2636 4877 2637 4898
rect 2672 4709 2673 4878
rect 2498 4879 2499 4898
rect 2673 4879 2674 4898
rect 2638 4709 2639 4882
rect 2736 4709 2737 4882
rect 2641 4709 2642 4884
rect 2733 4709 2734 4884
rect 2409 4709 2410 4886
rect 2734 4885 2735 4898
rect 2385 4709 2386 4888
rect 2408 4887 2409 4898
rect 2649 4887 2650 4898
rect 2694 4887 2695 4898
rect 2659 4709 2660 4890
rect 2667 4889 2668 4898
rect 2609 4891 2610 4898
rect 2658 4891 2659 4898
rect 2662 4709 2663 4892
rect 2687 4891 2688 4898
rect 2670 4893 2671 4898
rect 2690 4893 2691 4898
rect 2699 4709 2700 4894
rect 2714 4893 2715 4898
rect 2702 4709 2703 4896
rect 2717 4895 2718 4898
rect 2722 4709 2723 4896
rect 2723 4895 2724 4898
rect 2726 4709 2727 4896
rect 2737 4895 2738 4898
rect 2053 4902 2054 4905
rect 2225 4902 2226 4905
rect 2060 4902 2061 4907
rect 2240 4902 2241 4907
rect 2063 4902 2064 4909
rect 2164 4908 2165 5101
rect 2066 4910 2067 5101
rect 2188 4902 2189 4911
rect 2070 4902 2071 4913
rect 2237 4902 2238 4913
rect 2069 4914 2070 5101
rect 2081 4902 2082 4915
rect 2074 4902 2075 4917
rect 2182 4902 2183 4917
rect 2077 4902 2078 4919
rect 2191 4902 2192 4919
rect 2076 4920 2077 5101
rect 2080 4920 2081 5101
rect 2083 4920 2084 5101
rect 2200 4920 2201 5101
rect 2092 4922 2093 5101
rect 2093 4902 2094 4923
rect 2095 4922 2096 5101
rect 2246 4902 2247 4923
rect 2105 4924 2106 5101
rect 2234 4902 2235 4925
rect 2108 4926 2109 5101
rect 2264 4902 2265 4927
rect 2115 4902 2116 4929
rect 2255 4902 2256 4929
rect 2119 4902 2120 4931
rect 2234 4930 2235 5101
rect 2122 4902 2123 4933
rect 2243 4902 2244 4933
rect 2125 4902 2126 4935
rect 2138 4934 2139 5101
rect 2134 4902 2135 4937
rect 2207 4902 2208 4937
rect 2135 4938 2136 5101
rect 2158 4902 2159 4939
rect 2141 4902 2142 4941
rect 2151 4940 2152 5101
rect 2141 4942 2142 5101
rect 2396 4942 2397 5101
rect 2155 4902 2156 4945
rect 2324 4902 2325 4945
rect 2155 4946 2156 5101
rect 2285 4902 2286 4947
rect 2158 4948 2159 5101
rect 2279 4902 2280 4949
rect 2161 4950 2162 5101
rect 2219 4902 2220 4951
rect 2170 4952 2171 5101
rect 2216 4952 2217 5101
rect 2179 4954 2180 5101
rect 2228 4902 2229 4955
rect 2185 4956 2186 5101
rect 2249 4902 2250 4957
rect 2188 4958 2189 5101
rect 2252 4902 2253 4959
rect 2197 4902 2198 4961
rect 2387 4960 2388 5101
rect 2197 4962 2198 5101
rect 2261 4902 2262 4963
rect 2204 4902 2205 4965
rect 2579 4902 2580 4965
rect 2222 4966 2223 5101
rect 2288 4902 2289 4967
rect 2231 4968 2232 5101
rect 2297 4902 2298 4969
rect 2243 4970 2244 5101
rect 2300 4902 2301 4971
rect 2246 4972 2247 5101
rect 2303 4902 2304 4973
rect 2255 4974 2256 5101
rect 2318 4902 2319 4975
rect 2261 4976 2262 5101
rect 2330 4902 2331 4977
rect 2273 4978 2274 5101
rect 2360 4902 2361 4979
rect 2279 4980 2280 5101
rect 2615 4902 2616 4981
rect 2285 4982 2286 5101
rect 2348 4902 2349 4983
rect 2303 4984 2304 5101
rect 2372 4902 2373 4985
rect 2309 4986 2310 5101
rect 2378 4902 2379 4987
rect 2315 4988 2316 5101
rect 2599 4988 2600 5101
rect 2321 4902 2322 4991
rect 2399 4990 2400 5101
rect 2321 4992 2322 5101
rect 2390 4902 2391 4993
rect 2327 4994 2328 5101
rect 2444 4902 2445 4995
rect 2342 4902 2343 4997
rect 2549 4996 2550 5101
rect 2345 4998 2346 5101
rect 2408 4902 2409 4999
rect 2351 5000 2352 5101
rect 2414 4902 2415 5001
rect 2354 4902 2355 5003
rect 2580 5002 2581 5101
rect 2366 5004 2367 5101
rect 2429 4902 2430 5005
rect 2372 5006 2373 5101
rect 2435 4902 2436 5007
rect 2375 5008 2376 5101
rect 2438 4902 2439 5009
rect 2378 5010 2379 5101
rect 2616 5010 2617 5101
rect 2384 5012 2385 5101
rect 2558 4902 2559 5013
rect 2390 5014 2391 5101
rect 2459 4902 2460 5015
rect 2393 5016 2394 5101
rect 2680 4902 2681 5017
rect 2402 4902 2403 5019
rect 2737 4902 2738 5019
rect 2408 5020 2409 5101
rect 2477 4902 2478 5021
rect 2432 5022 2433 5101
rect 2495 4902 2496 5023
rect 2435 5024 2436 5101
rect 2498 4902 2499 5025
rect 2438 5026 2439 5101
rect 2576 4902 2577 5027
rect 2441 4902 2442 5029
rect 2444 5028 2445 5101
rect 2441 5030 2442 5101
rect 2465 4902 2466 5031
rect 2420 4902 2421 5033
rect 2465 5032 2466 5101
rect 2420 5034 2421 5101
rect 2483 4902 2484 5035
rect 2447 5036 2448 5101
rect 2552 5036 2553 5101
rect 2453 4902 2454 5039
rect 2701 4902 2702 5039
rect 2456 5040 2457 5101
rect 2519 4902 2520 5041
rect 2462 4902 2463 5043
rect 2646 4902 2647 5043
rect 2417 4902 2418 5045
rect 2462 5044 2463 5101
rect 2468 5044 2469 5101
rect 2727 4902 2728 5045
rect 2471 4902 2472 5047
rect 2519 5046 2520 5101
rect 2474 5048 2475 5101
rect 2531 4902 2532 5049
rect 2486 5050 2487 5101
rect 2507 4902 2508 5051
rect 2297 5052 2298 5101
rect 2507 5052 2508 5101
rect 2489 5054 2490 5101
rect 2510 4902 2511 5055
rect 2492 5056 2493 5101
rect 2546 4902 2547 5057
rect 2495 5058 2496 5101
rect 2571 5058 2572 5101
rect 2510 5060 2511 5101
rect 2567 4902 2568 5061
rect 2513 4902 2514 5063
rect 2624 4902 2625 5063
rect 2516 5064 2517 5101
rect 2582 4902 2583 5065
rect 2522 5066 2523 5101
rect 2585 4902 2586 5067
rect 2525 5068 2526 5101
rect 2588 4902 2589 5069
rect 2528 5070 2529 5101
rect 2591 4902 2592 5071
rect 2531 5072 2532 5101
rect 2620 5072 2621 5101
rect 2546 5074 2547 5101
rect 2609 4902 2610 5075
rect 2555 4902 2556 5077
rect 2642 5076 2643 5101
rect 2543 4902 2544 5079
rect 2556 5078 2557 5101
rect 2312 4902 2313 5081
rect 2543 5080 2544 5101
rect 2562 5080 2563 5101
rect 2618 4902 2619 5081
rect 2565 5082 2566 5101
rect 2594 4902 2595 5083
rect 2586 5084 2587 5101
rect 2649 4902 2650 5085
rect 2589 5086 2590 5101
rect 2652 4902 2653 5087
rect 2592 5088 2593 5101
rect 2670 4902 2671 5089
rect 2606 4902 2607 5091
rect 2655 4902 2656 5091
rect 2573 4902 2574 5093
rect 2606 5092 2607 5101
rect 2627 4902 2628 5093
rect 2639 4902 2640 5093
rect 2626 5094 2627 5101
rect 2720 4902 2721 5095
rect 2629 5096 2630 5101
rect 2717 4902 2718 5097
rect 2667 4902 2668 5099
rect 2690 4902 2691 5099
rect 2714 4902 2715 5099
rect 2723 4902 2724 5099
rect 2054 5107 2055 5274
rect 2161 5105 2162 5108
rect 2057 5109 2058 5274
rect 2119 5109 2120 5274
rect 2062 5105 2063 5112
rect 2164 5105 2165 5112
rect 2071 5113 2072 5274
rect 2135 5105 2136 5114
rect 2078 5115 2079 5274
rect 2092 5105 2093 5116
rect 2081 5117 2082 5274
rect 2095 5105 2096 5118
rect 2098 5105 2099 5118
rect 2200 5105 2201 5118
rect 2101 5105 2102 5120
rect 2197 5105 2198 5120
rect 2102 5121 2103 5274
rect 2114 5105 2115 5122
rect 2105 5105 2106 5124
rect 2131 5123 2132 5274
rect 2111 5105 2112 5126
rect 2185 5105 2186 5126
rect 2122 5127 2123 5274
rect 2138 5105 2139 5128
rect 2126 5105 2127 5130
rect 2144 5105 2145 5130
rect 2128 5131 2129 5274
rect 2275 5131 2276 5274
rect 2137 5133 2138 5274
rect 2151 5133 2152 5274
rect 2141 5105 2142 5136
rect 2234 5105 2235 5136
rect 2144 5137 2145 5274
rect 2516 5105 2517 5138
rect 2155 5105 2156 5140
rect 2586 5105 2587 5140
rect 2167 5105 2168 5142
rect 2399 5105 2400 5142
rect 2167 5143 2168 5274
rect 2179 5105 2180 5144
rect 2170 5105 2171 5146
rect 2396 5105 2397 5146
rect 2170 5147 2171 5274
rect 2188 5105 2189 5148
rect 2191 5147 2192 5274
rect 2222 5105 2223 5148
rect 2200 5149 2201 5274
rect 2231 5105 2232 5150
rect 2203 5151 2204 5274
rect 2243 5105 2244 5152
rect 2206 5153 2207 5274
rect 2246 5105 2247 5154
rect 2210 5105 2211 5156
rect 2281 5155 2282 5274
rect 2148 5105 2149 5158
rect 2209 5157 2210 5274
rect 2216 5105 2217 5158
rect 2218 5157 2219 5274
rect 2215 5159 2216 5274
rect 2255 5105 2256 5160
rect 2221 5161 2222 5274
rect 2261 5105 2262 5162
rect 2233 5163 2234 5274
rect 2279 5105 2280 5164
rect 2236 5165 2237 5274
rect 2465 5105 2466 5166
rect 2254 5167 2255 5274
rect 2303 5105 2304 5168
rect 2260 5169 2261 5274
rect 2327 5105 2328 5170
rect 2266 5171 2267 5274
rect 2602 5105 2603 5172
rect 2273 5105 2274 5174
rect 2552 5105 2553 5174
rect 2272 5175 2273 5274
rect 2462 5105 2463 5176
rect 2278 5177 2279 5274
rect 2486 5105 2487 5178
rect 2290 5179 2291 5274
rect 2321 5105 2322 5180
rect 2297 5105 2298 5182
rect 2540 5105 2541 5182
rect 2296 5183 2297 5274
rect 2595 5105 2596 5184
rect 2302 5185 2303 5274
rect 2345 5105 2346 5186
rect 2309 5105 2310 5188
rect 2571 5105 2572 5188
rect 2308 5189 2309 5274
rect 2568 5105 2569 5190
rect 2329 5191 2330 5274
rect 2384 5105 2385 5192
rect 2338 5193 2339 5274
rect 2606 5105 2607 5194
rect 2344 5195 2345 5274
rect 2387 5105 2388 5196
rect 2347 5197 2348 5274
rect 2444 5105 2445 5198
rect 2359 5199 2360 5274
rect 2432 5105 2433 5200
rect 2362 5201 2363 5274
rect 2366 5105 2367 5202
rect 2372 5105 2373 5202
rect 2497 5201 2498 5274
rect 2371 5203 2372 5274
rect 2592 5105 2593 5204
rect 2375 5105 2376 5206
rect 2485 5205 2486 5274
rect 2285 5105 2286 5208
rect 2374 5207 2375 5274
rect 2284 5209 2285 5274
rect 2315 5105 2316 5210
rect 2314 5211 2315 5274
rect 2351 5105 2352 5212
rect 2350 5213 2351 5274
rect 2447 5105 2448 5214
rect 2378 5105 2379 5216
rect 2609 5105 2610 5216
rect 2377 5217 2378 5274
rect 2456 5105 2457 5218
rect 2383 5219 2384 5274
rect 2438 5105 2439 5220
rect 2386 5221 2387 5274
rect 2457 5221 2458 5274
rect 2390 5105 2391 5224
rect 2556 5105 2557 5224
rect 2393 5105 2394 5226
rect 2424 5225 2425 5274
rect 2392 5227 2393 5274
rect 2642 5105 2643 5228
rect 2408 5105 2409 5230
rect 2433 5229 2434 5274
rect 2410 5231 2411 5274
rect 2549 5105 2550 5232
rect 2420 5105 2421 5234
rect 2515 5233 2516 5274
rect 2257 5235 2258 5274
rect 2420 5235 2421 5274
rect 2430 5235 2431 5274
rect 2522 5105 2523 5236
rect 2441 5105 2442 5238
rect 2543 5237 2544 5274
rect 2442 5239 2443 5274
rect 2546 5105 2547 5240
rect 2445 5241 2446 5274
rect 2460 5241 2461 5274
rect 2454 5243 2455 5274
rect 2528 5105 2529 5244
rect 2464 5245 2465 5274
rect 2525 5105 2526 5246
rect 2468 5105 2469 5248
rect 2529 5247 2530 5274
rect 2470 5249 2471 5274
rect 2562 5105 2563 5250
rect 2476 5251 2477 5274
rect 2632 5105 2633 5252
rect 2479 5253 2480 5274
rect 2629 5105 2630 5254
rect 2489 5105 2490 5256
rect 2504 5105 2505 5256
rect 2488 5257 2489 5274
rect 2589 5105 2590 5258
rect 2495 5105 2496 5260
rect 2507 5105 2508 5260
rect 2492 5105 2493 5262
rect 2494 5261 2495 5274
rect 2491 5263 2492 5274
rect 2510 5105 2511 5264
rect 2482 5265 2483 5274
rect 2511 5265 2512 5274
rect 2519 5105 2520 5266
rect 2536 5265 2537 5274
rect 2435 5105 2436 5268
rect 2518 5267 2519 5274
rect 2531 5105 2532 5268
rect 2613 5105 2614 5268
rect 2474 5105 2475 5270
rect 2532 5269 2533 5274
rect 2473 5271 2474 5274
rect 2565 5105 2566 5272
rect 2620 5105 2621 5272
rect 2626 5105 2627 5272
rect 2047 5278 2048 5281
rect 2119 5278 2120 5281
rect 2050 5280 2051 5419
rect 2050 5278 2051 5281
rect 2074 5278 2075 5283
rect 2092 5278 2093 5283
rect 2075 5284 2076 5419
rect 2122 5278 2123 5285
rect 2079 5286 2080 5419
rect 2085 5278 2086 5287
rect 2082 5288 2083 5419
rect 2089 5288 2090 5419
rect 2092 5288 2093 5419
rect 2099 5278 2100 5289
rect 2102 5288 2103 5419
rect 2170 5278 2171 5289
rect 2106 5290 2107 5419
rect 2218 5278 2219 5291
rect 2113 5292 2114 5419
rect 2134 5292 2135 5419
rect 2116 5278 2117 5295
rect 2196 5294 2197 5419
rect 2119 5296 2120 5419
rect 2151 5278 2152 5297
rect 2122 5298 2123 5419
rect 2128 5278 2129 5299
rect 2128 5300 2129 5419
rect 2131 5278 2132 5301
rect 2131 5302 2132 5419
rect 2141 5278 2142 5303
rect 2138 5304 2139 5419
rect 2226 5304 2227 5419
rect 2148 5306 2149 5419
rect 2163 5306 2164 5419
rect 2155 5278 2156 5309
rect 2221 5278 2222 5309
rect 2157 5310 2158 5419
rect 2272 5278 2273 5311
rect 2167 5278 2168 5313
rect 2175 5312 2176 5419
rect 2169 5314 2170 5419
rect 2209 5278 2210 5315
rect 2203 5278 2204 5317
rect 2208 5316 2209 5419
rect 2206 5278 2207 5319
rect 2211 5318 2212 5419
rect 2215 5278 2216 5319
rect 2223 5318 2224 5419
rect 2200 5278 2201 5321
rect 2214 5320 2215 5419
rect 2191 5278 2192 5323
rect 2199 5322 2200 5419
rect 2217 5322 2218 5419
rect 2247 5322 2248 5419
rect 2229 5324 2230 5419
rect 2278 5278 2279 5325
rect 2233 5278 2234 5327
rect 2244 5326 2245 5419
rect 2238 5328 2239 5419
rect 2275 5278 2276 5329
rect 2241 5330 2242 5419
rect 2281 5278 2282 5331
rect 2254 5278 2255 5333
rect 2286 5332 2287 5419
rect 2257 5278 2258 5335
rect 2508 5278 2509 5335
rect 2260 5278 2261 5337
rect 2410 5278 2411 5337
rect 2259 5338 2260 5419
rect 2374 5278 2375 5339
rect 2266 5278 2267 5341
rect 2277 5340 2278 5419
rect 2265 5342 2266 5419
rect 2350 5278 2351 5343
rect 2271 5344 2272 5419
rect 2402 5344 2403 5419
rect 2296 5278 2297 5347
rect 2331 5346 2332 5419
rect 2302 5278 2303 5349
rect 2546 5278 2547 5349
rect 2308 5278 2309 5351
rect 2334 5350 2335 5419
rect 2290 5278 2291 5353
rect 2307 5352 2308 5419
rect 2289 5354 2290 5419
rect 2511 5278 2512 5355
rect 2314 5278 2315 5357
rect 2522 5278 2523 5357
rect 2319 5358 2320 5419
rect 2398 5358 2399 5419
rect 2322 5360 2323 5419
rect 2347 5278 2348 5361
rect 2325 5362 2326 5419
rect 2362 5278 2363 5363
rect 2338 5278 2339 5365
rect 2340 5364 2341 5419
rect 2344 5278 2345 5365
rect 2352 5364 2353 5419
rect 2359 5278 2360 5365
rect 2515 5278 2516 5365
rect 2368 5278 2369 5367
rect 2417 5278 2418 5367
rect 2367 5368 2368 5419
rect 2460 5278 2461 5369
rect 2371 5278 2372 5371
rect 2379 5370 2380 5419
rect 2370 5372 2371 5419
rect 2445 5278 2446 5373
rect 2386 5278 2387 5375
rect 2525 5278 2526 5375
rect 2383 5278 2384 5377
rect 2385 5376 2386 5419
rect 2382 5378 2383 5419
rect 2395 5378 2396 5419
rect 2388 5380 2389 5419
rect 2442 5278 2443 5381
rect 2392 5278 2393 5383
rect 2529 5278 2530 5383
rect 2414 5384 2415 5419
rect 2430 5278 2431 5385
rect 2417 5386 2418 5419
rect 2433 5278 2434 5387
rect 2420 5278 2421 5389
rect 2476 5278 2477 5389
rect 2313 5390 2314 5419
rect 2420 5390 2421 5419
rect 2427 5390 2428 5419
rect 2442 5390 2443 5419
rect 2430 5392 2431 5419
rect 2482 5278 2483 5393
rect 2329 5278 2330 5395
rect 2482 5394 2483 5419
rect 2328 5396 2329 5419
rect 2485 5278 2486 5397
rect 2433 5398 2434 5419
rect 2470 5278 2471 5399
rect 2436 5400 2437 5419
rect 2501 5278 2502 5401
rect 2445 5402 2446 5419
rect 2488 5278 2489 5403
rect 2448 5404 2449 5419
rect 2491 5278 2492 5405
rect 2454 5278 2455 5407
rect 2465 5406 2466 5419
rect 2473 5278 2474 5407
rect 2536 5278 2537 5407
rect 2284 5278 2285 5409
rect 2472 5408 2473 5419
rect 2283 5410 2284 5419
rect 2424 5278 2425 5411
rect 2377 5278 2378 5413
rect 2423 5412 2424 5419
rect 2479 5278 2480 5413
rect 2532 5278 2533 5413
rect 2491 5414 2492 5419
rect 2500 5414 2501 5419
rect 2494 5416 2495 5419
rect 2497 5416 2498 5419
rect 2065 5423 2066 5426
rect 2072 5423 2073 5426
rect 2079 5423 2080 5426
rect 2128 5423 2129 5426
rect 2099 5423 2100 5428
rect 2113 5423 2114 5428
rect 2106 5423 2107 5430
rect 2172 5429 2173 5552
rect 2111 5431 2112 5552
rect 2178 5431 2179 5552
rect 2115 5433 2116 5552
rect 2214 5423 2215 5434
rect 2119 5423 2120 5436
rect 2181 5435 2182 5552
rect 2125 5423 2126 5438
rect 2251 5437 2252 5552
rect 2127 5439 2128 5552
rect 2208 5423 2209 5440
rect 2131 5423 2132 5442
rect 2220 5423 2221 5442
rect 2130 5443 2131 5552
rect 2211 5423 2212 5444
rect 2141 5445 2142 5552
rect 2232 5423 2233 5446
rect 2145 5423 2146 5448
rect 2157 5423 2158 5448
rect 2138 5423 2139 5450
rect 2144 5449 2145 5552
rect 2148 5449 2149 5552
rect 2241 5423 2242 5450
rect 2151 5451 2152 5552
rect 2257 5451 2258 5552
rect 2163 5423 2164 5454
rect 2166 5453 2167 5552
rect 2175 5423 2176 5454
rect 2205 5453 2206 5552
rect 2196 5423 2197 5456
rect 2221 5455 2222 5552
rect 2118 5457 2119 5552
rect 2196 5457 2197 5552
rect 2223 5423 2224 5458
rect 2254 5457 2255 5552
rect 2199 5423 2200 5460
rect 2224 5459 2225 5552
rect 2184 5423 2185 5462
rect 2199 5461 2200 5552
rect 2169 5423 2170 5464
rect 2184 5463 2185 5552
rect 2226 5423 2227 5464
rect 2227 5463 2228 5552
rect 2229 5423 2230 5464
rect 2305 5463 2306 5552
rect 2238 5423 2239 5466
rect 2275 5465 2276 5552
rect 2247 5423 2248 5468
rect 2265 5423 2266 5468
rect 2248 5469 2249 5552
rect 2322 5423 2323 5470
rect 2134 5423 2135 5472
rect 2323 5471 2324 5552
rect 2259 5423 2260 5474
rect 2468 5423 2469 5474
rect 2260 5475 2261 5552
rect 2382 5423 2383 5476
rect 2218 5477 2219 5552
rect 2383 5477 2384 5552
rect 2277 5423 2278 5480
rect 2338 5479 2339 5552
rect 2215 5481 2216 5552
rect 2278 5481 2279 5552
rect 2283 5423 2284 5482
rect 2391 5423 2392 5482
rect 2284 5483 2285 5552
rect 2359 5483 2360 5552
rect 2286 5423 2287 5486
rect 2296 5485 2297 5552
rect 2287 5487 2288 5552
rect 2313 5423 2314 5488
rect 2289 5423 2290 5490
rect 2419 5489 2420 5552
rect 2307 5423 2308 5492
rect 2454 5423 2455 5492
rect 2244 5423 2245 5494
rect 2308 5493 2309 5552
rect 2245 5495 2246 5552
rect 2319 5423 2320 5496
rect 2317 5497 2318 5552
rect 2389 5497 2390 5552
rect 2328 5423 2329 5500
rect 2410 5499 2411 5552
rect 2271 5423 2272 5502
rect 2329 5501 2330 5552
rect 2235 5423 2236 5504
rect 2272 5503 2273 5552
rect 2334 5423 2335 5504
rect 2335 5503 2336 5552
rect 2347 5503 2348 5552
rect 2423 5423 2424 5504
rect 2352 5423 2353 5506
rect 2404 5505 2405 5552
rect 2370 5423 2371 5508
rect 2402 5423 2403 5508
rect 2374 5509 2375 5552
rect 2417 5423 2418 5510
rect 2379 5423 2380 5512
rect 2395 5423 2396 5512
rect 2380 5513 2381 5552
rect 2438 5513 2439 5552
rect 2385 5423 2386 5516
rect 2483 5515 2484 5552
rect 2365 5517 2366 5552
rect 2386 5517 2387 5552
rect 2407 5517 2408 5552
rect 2430 5423 2431 5518
rect 2340 5423 2341 5520
rect 2431 5519 2432 5552
rect 2341 5521 2342 5552
rect 2422 5521 2423 5552
rect 2414 5423 2415 5524
rect 2455 5523 2456 5552
rect 2413 5525 2414 5552
rect 2433 5423 2434 5526
rect 2353 5527 2354 5552
rect 2434 5527 2435 5552
rect 2416 5529 2417 5552
rect 2436 5423 2437 5530
rect 2425 5531 2426 5552
rect 2452 5531 2453 5552
rect 2428 5533 2429 5552
rect 2445 5423 2446 5534
rect 2367 5423 2368 5536
rect 2445 5535 2446 5552
rect 2441 5537 2442 5552
rect 2448 5423 2449 5538
rect 2325 5423 2326 5540
rect 2448 5539 2449 5552
rect 2326 5541 2327 5552
rect 2398 5423 2399 5542
rect 2331 5423 2332 5544
rect 2398 5543 2399 5552
rect 2476 5543 2477 5552
rect 2494 5423 2495 5544
rect 2487 5545 2488 5552
rect 2494 5545 2495 5552
rect 2491 5423 2492 5548
rect 2514 5423 2515 5548
rect 2500 5423 2501 5550
rect 2504 5423 2505 5550
rect 2089 5556 2090 5559
rect 2192 5558 2193 5669
rect 2092 5560 2093 5669
rect 2189 5560 2190 5669
rect 2101 5556 2102 5563
rect 2205 5556 2206 5563
rect 2111 5556 2112 5565
rect 2172 5556 2173 5565
rect 2104 5566 2105 5669
rect 2111 5566 2112 5669
rect 2118 5566 2119 5669
rect 2196 5556 2197 5567
rect 2132 5568 2133 5669
rect 2153 5568 2154 5669
rect 2134 5556 2135 5571
rect 2248 5556 2249 5571
rect 2137 5556 2138 5573
rect 2221 5556 2222 5573
rect 2141 5556 2142 5575
rect 2278 5556 2279 5575
rect 2148 5556 2149 5577
rect 2272 5556 2273 5577
rect 2159 5578 2160 5669
rect 2199 5556 2200 5579
rect 2162 5580 2163 5669
rect 2184 5556 2185 5581
rect 2166 5556 2167 5583
rect 2222 5582 2223 5669
rect 2171 5584 2172 5669
rect 2178 5556 2179 5585
rect 2174 5586 2175 5669
rect 2181 5556 2182 5587
rect 2183 5586 2184 5669
rect 2257 5556 2258 5587
rect 2195 5588 2196 5669
rect 2211 5556 2212 5589
rect 2198 5590 2199 5669
rect 2438 5556 2439 5591
rect 2204 5592 2205 5669
rect 2224 5556 2225 5593
rect 2208 5556 2209 5595
rect 2326 5556 2327 5595
rect 2144 5556 2145 5597
rect 2207 5596 2208 5669
rect 2216 5596 2217 5669
rect 2227 5556 2228 5597
rect 2225 5598 2226 5669
rect 2275 5556 2276 5599
rect 2228 5600 2229 5669
rect 2254 5556 2255 5601
rect 2231 5602 2232 5669
rect 2241 5602 2242 5669
rect 2233 5556 2234 5605
rect 2289 5604 2290 5669
rect 2234 5606 2235 5669
rect 2251 5556 2252 5607
rect 2236 5556 2237 5609
rect 2292 5608 2293 5669
rect 2237 5610 2238 5669
rect 2262 5610 2263 5669
rect 2247 5612 2248 5669
rect 2305 5556 2306 5613
rect 2245 5556 2246 5615
rect 2304 5614 2305 5669
rect 2284 5556 2285 5617
rect 2323 5556 2324 5617
rect 2283 5618 2284 5669
rect 2338 5556 2339 5619
rect 2287 5556 2288 5621
rect 2317 5556 2318 5621
rect 2286 5622 2287 5669
rect 2329 5556 2330 5623
rect 2296 5556 2297 5625
rect 2298 5624 2299 5669
rect 2260 5556 2261 5627
rect 2295 5626 2296 5669
rect 2259 5628 2260 5669
rect 2308 5556 2309 5629
rect 2307 5630 2308 5669
rect 2365 5556 2366 5631
rect 2310 5632 2311 5669
rect 2419 5556 2420 5633
rect 2322 5634 2323 5669
rect 2448 5556 2449 5635
rect 2325 5636 2326 5669
rect 2341 5556 2342 5637
rect 2335 5556 2336 5639
rect 2365 5638 2366 5669
rect 2340 5640 2341 5669
rect 2344 5640 2345 5669
rect 2347 5556 2348 5641
rect 2393 5640 2394 5669
rect 2350 5642 2351 5669
rect 2416 5556 2417 5643
rect 2353 5556 2354 5645
rect 2400 5644 2401 5669
rect 2356 5646 2357 5669
rect 2383 5556 2384 5647
rect 2359 5556 2360 5649
rect 2378 5648 2379 5669
rect 2359 5650 2360 5669
rect 2374 5556 2375 5651
rect 2369 5652 2370 5669
rect 2380 5556 2381 5653
rect 2372 5654 2373 5669
rect 2387 5654 2388 5669
rect 2375 5656 2376 5669
rect 2407 5556 2408 5657
rect 2390 5658 2391 5669
rect 2413 5556 2414 5659
rect 2404 5556 2405 5661
rect 2487 5556 2488 5661
rect 2406 5662 2407 5669
rect 2425 5556 2426 5663
rect 2410 5556 2411 5665
rect 2445 5556 2446 5665
rect 2428 5556 2429 5667
rect 2441 5556 2442 5667
rect 2473 5556 2474 5667
rect 2483 5556 2484 5667
rect 2089 5673 2090 5676
rect 2192 5673 2193 5676
rect 2092 5673 2093 5678
rect 2099 5677 2100 5756
rect 2104 5673 2105 5678
rect 2171 5673 2172 5678
rect 2096 5679 2097 5756
rect 2103 5679 2104 5756
rect 2106 5679 2107 5756
rect 2216 5673 2217 5680
rect 2108 5673 2109 5682
rect 2174 5673 2175 5682
rect 2109 5683 2110 5756
rect 2189 5673 2190 5684
rect 2115 5685 2116 5756
rect 2122 5685 2123 5756
rect 2118 5673 2119 5688
rect 2195 5673 2196 5688
rect 2125 5673 2126 5690
rect 2153 5673 2154 5690
rect 2126 5691 2127 5756
rect 2204 5673 2205 5692
rect 2129 5673 2130 5694
rect 2207 5673 2208 5694
rect 2138 5695 2139 5756
rect 2198 5673 2199 5696
rect 2141 5673 2142 5698
rect 2183 5673 2184 5698
rect 2132 5673 2133 5700
rect 2141 5699 2142 5756
rect 2144 5673 2145 5700
rect 2231 5673 2232 5700
rect 2144 5701 2145 5756
rect 2228 5673 2229 5702
rect 2151 5703 2152 5756
rect 2190 5703 2191 5756
rect 2154 5705 2155 5756
rect 2225 5673 2226 5706
rect 2157 5707 2158 5756
rect 2259 5673 2260 5708
rect 2163 5709 2164 5756
rect 2262 5673 2263 5710
rect 2172 5711 2173 5756
rect 2289 5673 2290 5712
rect 2181 5713 2182 5756
rect 2295 5673 2296 5714
rect 2184 5715 2185 5756
rect 2298 5673 2299 5716
rect 2193 5717 2194 5756
rect 2362 5673 2363 5718
rect 2196 5719 2197 5756
rect 2283 5673 2284 5720
rect 2205 5721 2206 5756
rect 2292 5673 2293 5722
rect 2208 5723 2209 5756
rect 2247 5673 2248 5724
rect 2211 5725 2212 5756
rect 2359 5673 2360 5726
rect 2222 5673 2223 5728
rect 2400 5673 2401 5728
rect 2221 5729 2222 5756
rect 2322 5673 2323 5730
rect 2228 5731 2229 5756
rect 2325 5673 2326 5732
rect 2234 5733 2235 5756
rect 2375 5673 2376 5734
rect 2237 5735 2238 5756
rect 2378 5673 2379 5736
rect 2244 5673 2245 5738
rect 2304 5673 2305 5738
rect 2246 5739 2247 5756
rect 2396 5673 2397 5740
rect 2249 5741 2250 5756
rect 2387 5673 2388 5742
rect 2255 5743 2256 5756
rect 2310 5673 2311 5744
rect 2262 5745 2263 5756
rect 2390 5673 2391 5746
rect 2286 5673 2287 5748
rect 2340 5673 2341 5748
rect 2307 5673 2308 5750
rect 2413 5673 2414 5750
rect 2350 5673 2351 5752
rect 2393 5673 2394 5752
rect 2356 5673 2357 5754
rect 2369 5673 2370 5754
rect 2065 5760 2066 5763
rect 2072 5760 2073 5763
rect 2089 5760 2090 5763
rect 2109 5760 2110 5763
rect 2119 5760 2120 5763
rect 2141 5760 2142 5763
rect 2122 5760 2123 5765
rect 2157 5760 2158 5765
rect 2126 5760 2127 5767
rect 2138 5760 2139 5767
rect 2147 5760 2148 5767
rect 2151 5760 2152 5767
rect 2153 5766 2154 5787
rect 2156 5766 2157 5787
rect 2159 5766 2160 5787
rect 2234 5760 2235 5767
rect 2166 5768 2167 5787
rect 2181 5760 2182 5769
rect 2169 5770 2170 5787
rect 2214 5760 2215 5771
rect 2172 5760 2173 5773
rect 2190 5760 2191 5773
rect 2184 5760 2185 5775
rect 2221 5760 2222 5775
rect 2193 5760 2194 5777
rect 2208 5760 2209 5777
rect 2196 5760 2197 5779
rect 2224 5760 2225 5779
rect 2211 5760 2212 5781
rect 2231 5760 2232 5781
rect 2237 5760 2238 5781
rect 2255 5760 2256 5781
rect 2246 5760 2247 5783
rect 2262 5760 2263 5783
rect 2249 5760 2250 5785
rect 2259 5760 2260 5785
rect 2146 5791 2147 5794
rect 2150 5791 2151 5794
rect 2153 5793 2154 5796
rect 2153 5791 2154 5794
rect 2156 5791 2157 5794
rect 2159 5791 2160 5794
rect 2143 5800 2144 5803
rect 2153 5800 2154 5803
<< via >>
rect 2134 1007 2135 1008
rect 2137 1007 2138 1008
rect 2077 1017 2078 1018
rect 2147 1017 2148 1018
rect 2087 1019 2088 1020
rect 2120 1019 2121 1020
rect 2101 1021 2102 1022
rect 2129 1021 2130 1022
rect 2108 1023 2109 1024
rect 2111 1023 2112 1024
rect 2131 1023 2132 1024
rect 2174 1023 2175 1024
rect 2091 1025 2092 1026
rect 2132 1025 2133 1026
rect 2134 1025 2135 1026
rect 2198 1025 2199 1026
rect 2135 1027 2136 1028
rect 2207 1027 2208 1028
rect 2137 1029 2138 1030
rect 2183 1029 2184 1030
rect 2138 1031 2139 1032
rect 2159 1031 2160 1032
rect 2140 1033 2141 1034
rect 2211 1033 2212 1034
rect 2143 1035 2144 1036
rect 2180 1035 2181 1036
rect 2150 1037 2151 1038
rect 2171 1037 2172 1038
rect 2155 1039 2156 1040
rect 2201 1039 2202 1040
rect 2156 1041 2157 1042
rect 2227 1041 2228 1042
rect 2162 1043 2163 1044
rect 2214 1043 2215 1044
rect 2195 1045 2196 1046
rect 2221 1045 2222 1046
rect 2224 1045 2225 1046
rect 2243 1045 2244 1046
rect 2233 1047 2234 1048
rect 2236 1047 2237 1048
rect 2246 1047 2247 1048
rect 2274 1047 2275 1048
rect 2255 1049 2256 1050
rect 2264 1049 2265 1050
rect 2258 1051 2259 1052
rect 2261 1051 2262 1052
rect 2084 1060 2085 1061
rect 2230 1060 2231 1061
rect 2084 1062 2085 1063
rect 2143 1062 2144 1063
rect 2087 1064 2088 1065
rect 2159 1064 2160 1065
rect 2077 1066 2078 1067
rect 2158 1066 2159 1067
rect 2078 1068 2079 1069
rect 2389 1068 2390 1069
rect 2098 1070 2099 1071
rect 2311 1070 2312 1071
rect 2114 1072 2115 1073
rect 2251 1072 2252 1073
rect 2124 1074 2125 1075
rect 2156 1074 2157 1075
rect 2129 1076 2130 1077
rect 2176 1076 2177 1077
rect 2138 1078 2139 1079
rect 2155 1078 2156 1079
rect 2152 1080 2153 1081
rect 2162 1080 2163 1081
rect 2120 1082 2121 1083
rect 2161 1082 2162 1083
rect 2111 1084 2112 1085
rect 2121 1084 2122 1085
rect 2165 1084 2166 1085
rect 2218 1084 2219 1085
rect 2168 1086 2169 1087
rect 2266 1086 2267 1087
rect 2174 1088 2175 1089
rect 2218 1088 2219 1089
rect 2180 1090 2181 1091
rect 2278 1090 2279 1091
rect 2095 1092 2096 1093
rect 2179 1092 2180 1093
rect 2201 1092 2202 1093
rect 2227 1092 2228 1093
rect 2207 1094 2208 1095
rect 2281 1094 2282 1095
rect 2185 1096 2186 1097
rect 2206 1096 2207 1097
rect 2221 1096 2222 1097
rect 2290 1096 2291 1097
rect 2224 1098 2225 1099
rect 2323 1098 2324 1099
rect 2233 1100 2234 1101
rect 2317 1100 2318 1101
rect 2091 1102 2092 1103
rect 2233 1102 2234 1103
rect 2236 1102 2237 1103
rect 2353 1102 2354 1103
rect 2147 1104 2148 1105
rect 2236 1104 2237 1105
rect 2239 1104 2240 1105
rect 2350 1104 2351 1105
rect 2167 1106 2168 1107
rect 2239 1106 2240 1107
rect 2243 1106 2244 1107
rect 2341 1106 2342 1107
rect 2171 1108 2172 1109
rect 2242 1108 2243 1109
rect 2132 1110 2133 1111
rect 2170 1110 2171 1111
rect 2246 1110 2247 1111
rect 2338 1110 2339 1111
rect 2183 1112 2184 1113
rect 2245 1112 2246 1113
rect 2182 1114 2183 1115
rect 2195 1114 2196 1115
rect 2080 1116 2081 1117
rect 2194 1116 2195 1117
rect 2081 1118 2082 1119
rect 2127 1118 2128 1119
rect 2255 1118 2256 1119
rect 2380 1118 2381 1119
rect 2211 1120 2212 1121
rect 2254 1120 2255 1121
rect 2198 1122 2199 1123
rect 2212 1122 2213 1123
rect 2258 1122 2259 1123
rect 2383 1122 2384 1123
rect 2268 1124 2269 1125
rect 2362 1124 2363 1125
rect 2088 1126 2089 1127
rect 2269 1126 2270 1127
rect 2271 1126 2272 1127
rect 2386 1126 2387 1127
rect 2274 1128 2275 1129
rect 2406 1128 2407 1129
rect 2299 1130 2300 1131
rect 2430 1130 2431 1131
rect 2335 1132 2336 1133
rect 2393 1132 2394 1133
rect 2371 1134 2372 1135
rect 2440 1134 2441 1135
rect 2409 1136 2410 1137
rect 2416 1136 2417 1137
rect 2068 1145 2069 1146
rect 2248 1145 2249 1146
rect 2072 1147 2073 1148
rect 2275 1147 2276 1148
rect 2078 1149 2079 1150
rect 2093 1149 2094 1150
rect 2084 1151 2085 1152
rect 2272 1151 2273 1152
rect 2087 1153 2088 1154
rect 2302 1153 2303 1154
rect 2098 1155 2099 1156
rect 2293 1155 2294 1156
rect 2099 1157 2100 1158
rect 2230 1157 2231 1158
rect 2108 1159 2109 1160
rect 2179 1159 2180 1160
rect 2117 1161 2118 1162
rect 2145 1161 2146 1162
rect 2121 1163 2122 1164
rect 2404 1163 2405 1164
rect 2124 1165 2125 1166
rect 2278 1165 2279 1166
rect 2135 1167 2136 1168
rect 2266 1167 2267 1168
rect 2137 1169 2138 1170
rect 2284 1169 2285 1170
rect 2143 1171 2144 1172
rect 2172 1171 2173 1172
rect 2152 1173 2153 1174
rect 2199 1173 2200 1174
rect 2155 1175 2156 1176
rect 2287 1175 2288 1176
rect 2081 1177 2082 1178
rect 2154 1177 2155 1178
rect 2161 1177 2162 1178
rect 2278 1177 2279 1178
rect 2127 1179 2128 1180
rect 2160 1179 2161 1180
rect 2128 1181 2129 1182
rect 2314 1181 2315 1182
rect 2167 1183 2168 1184
rect 2245 1183 2246 1184
rect 2065 1185 2066 1186
rect 2245 1185 2246 1186
rect 2062 1187 2063 1188
rect 2066 1187 2067 1188
rect 2176 1187 2177 1188
rect 2220 1187 2221 1188
rect 2178 1189 2179 1190
rect 2389 1189 2390 1190
rect 2182 1191 2183 1192
rect 2194 1191 2195 1192
rect 2206 1191 2207 1192
rect 2263 1191 2264 1192
rect 2212 1193 2213 1194
rect 2296 1193 2297 1194
rect 2170 1195 2171 1196
rect 2211 1195 2212 1196
rect 2233 1195 2234 1196
rect 2308 1195 2309 1196
rect 2236 1197 2237 1198
rect 2257 1197 2258 1198
rect 2239 1199 2240 1200
rect 2329 1199 2330 1200
rect 2242 1201 2243 1202
rect 2332 1201 2333 1202
rect 2251 1203 2252 1204
rect 2326 1203 2327 1204
rect 2269 1205 2270 1206
rect 2356 1205 2357 1206
rect 2080 1207 2081 1208
rect 2269 1207 2270 1208
rect 2281 1207 2282 1208
rect 2359 1207 2360 1208
rect 2281 1209 2282 1210
rect 2443 1209 2444 1210
rect 2290 1211 2291 1212
rect 2374 1211 2375 1212
rect 2114 1213 2115 1214
rect 2290 1213 2291 1214
rect 2114 1215 2115 1216
rect 2181 1215 2182 1216
rect 2299 1215 2300 1216
rect 2386 1215 2387 1216
rect 2311 1217 2312 1218
rect 2398 1217 2399 1218
rect 2117 1219 2118 1220
rect 2311 1219 2312 1220
rect 2317 1219 2318 1220
rect 2446 1219 2447 1220
rect 2131 1221 2132 1222
rect 2317 1221 2318 1222
rect 2335 1221 2336 1222
rect 2443 1221 2444 1222
rect 2218 1223 2219 1224
rect 2335 1223 2336 1224
rect 2158 1225 2159 1226
rect 2217 1225 2218 1226
rect 2338 1225 2339 1226
rect 2518 1225 2519 1226
rect 2341 1227 2342 1228
rect 2428 1227 2429 1228
rect 2254 1229 2255 1230
rect 2341 1229 2342 1230
rect 2350 1229 2351 1230
rect 2458 1229 2459 1230
rect 2353 1231 2354 1232
rect 2461 1231 2462 1232
rect 2142 1233 2143 1234
rect 2353 1233 2354 1234
rect 2362 1233 2363 1234
rect 2464 1233 2465 1234
rect 2371 1235 2372 1236
rect 2486 1235 2487 1236
rect 2380 1237 2381 1238
rect 2502 1237 2503 1238
rect 2383 1239 2384 1240
rect 2489 1239 2490 1240
rect 2377 1241 2378 1242
rect 2383 1241 2384 1242
rect 2396 1241 2397 1242
rect 2440 1241 2441 1242
rect 2406 1243 2407 1244
rect 2409 1243 2410 1244
rect 2410 1245 2411 1246
rect 2470 1245 2471 1246
rect 2430 1247 2431 1248
rect 2492 1247 2493 1248
rect 2323 1249 2324 1250
rect 2431 1249 2432 1250
rect 2433 1249 2434 1250
rect 2467 1249 2468 1250
rect 2483 1249 2484 1250
rect 2563 1249 2564 1250
rect 2515 1251 2516 1252
rect 2521 1251 2522 1252
rect 2059 1260 2060 1261
rect 2281 1260 2282 1261
rect 2068 1262 2069 1263
rect 2108 1262 2109 1263
rect 2073 1264 2074 1265
rect 2345 1264 2346 1265
rect 2072 1266 2073 1267
rect 2245 1266 2246 1267
rect 2080 1268 2081 1269
rect 2204 1268 2205 1269
rect 2086 1270 2087 1271
rect 2201 1270 2202 1271
rect 2093 1272 2094 1273
rect 2112 1272 2113 1273
rect 2096 1274 2097 1275
rect 2369 1274 2370 1275
rect 2118 1276 2119 1277
rect 2302 1276 2303 1277
rect 2124 1278 2125 1279
rect 2408 1278 2409 1279
rect 2125 1280 2126 1281
rect 2311 1280 2312 1281
rect 2128 1282 2129 1283
rect 2351 1282 2352 1283
rect 2142 1284 2143 1285
rect 2326 1284 2327 1285
rect 2131 1286 2132 1287
rect 2141 1286 2142 1287
rect 2160 1286 2161 1287
rect 2231 1286 2232 1287
rect 2165 1288 2166 1289
rect 2172 1288 2173 1289
rect 2181 1288 2182 1289
rect 2207 1288 2208 1289
rect 2189 1290 2190 1291
rect 2199 1290 2200 1291
rect 2211 1290 2212 1291
rect 2240 1290 2241 1291
rect 2220 1292 2221 1293
rect 2252 1292 2253 1293
rect 2226 1294 2227 1295
rect 2329 1294 2330 1295
rect 2178 1296 2179 1297
rect 2225 1296 2226 1297
rect 2154 1298 2155 1299
rect 2177 1298 2178 1299
rect 2233 1298 2234 1299
rect 2353 1298 2354 1299
rect 2217 1300 2218 1301
rect 2234 1300 2235 1301
rect 2272 1300 2273 1301
rect 2312 1300 2313 1301
rect 2138 1302 2139 1303
rect 2273 1302 2274 1303
rect 2275 1302 2276 1303
rect 2321 1302 2322 1303
rect 2248 1304 2249 1305
rect 2276 1304 2277 1305
rect 2278 1304 2279 1305
rect 2348 1304 2349 1305
rect 2284 1306 2285 1307
rect 2392 1306 2393 1307
rect 2287 1308 2288 1309
rect 2390 1308 2391 1309
rect 2290 1310 2291 1311
rect 2327 1310 2328 1311
rect 2079 1312 2080 1313
rect 2291 1312 2292 1313
rect 2293 1312 2294 1313
rect 2372 1312 2373 1313
rect 2296 1314 2297 1315
rect 2363 1314 2364 1315
rect 2257 1316 2258 1317
rect 2297 1316 2298 1317
rect 2096 1318 2097 1319
rect 2258 1318 2259 1319
rect 2314 1318 2315 1319
rect 2339 1318 2340 1319
rect 2263 1320 2264 1321
rect 2315 1320 2316 1321
rect 2093 1322 2094 1323
rect 2264 1322 2265 1323
rect 2317 1322 2318 1323
rect 2354 1322 2355 1323
rect 2335 1324 2336 1325
rect 2381 1324 2382 1325
rect 2236 1326 2237 1327
rect 2336 1326 2337 1327
rect 2341 1326 2342 1327
rect 2393 1326 2394 1327
rect 2356 1328 2357 1329
rect 2396 1328 2397 1329
rect 2308 1330 2309 1331
rect 2357 1330 2358 1331
rect 2269 1332 2270 1333
rect 2309 1332 2310 1333
rect 2100 1334 2101 1335
rect 2270 1334 2271 1335
rect 2359 1334 2360 1335
rect 2417 1334 2418 1335
rect 2114 1336 2115 1337
rect 2360 1336 2361 1337
rect 2374 1336 2375 1337
rect 2438 1336 2439 1337
rect 2332 1338 2333 1339
rect 2375 1338 2376 1339
rect 2121 1340 2122 1341
rect 2333 1340 2334 1341
rect 2377 1340 2378 1341
rect 2426 1340 2427 1341
rect 2410 1342 2411 1343
rect 2471 1342 2472 1343
rect 2435 1344 2436 1345
rect 2589 1344 2590 1345
rect 2440 1346 2441 1347
rect 2534 1346 2535 1347
rect 2386 1348 2387 1349
rect 2441 1348 2442 1349
rect 2090 1350 2091 1351
rect 2387 1350 2388 1351
rect 2443 1350 2444 1351
rect 2495 1350 2496 1351
rect 2446 1352 2447 1353
rect 2507 1352 2508 1353
rect 2447 1354 2448 1355
rect 2555 1354 2556 1355
rect 2458 1356 2459 1357
rect 2519 1356 2520 1357
rect 2398 1358 2399 1359
rect 2459 1358 2460 1359
rect 2145 1360 2146 1361
rect 2399 1360 2400 1361
rect 2461 1360 2462 1361
rect 2522 1360 2523 1361
rect 2464 1362 2465 1363
rect 2525 1362 2526 1363
rect 2404 1364 2405 1365
rect 2465 1364 2466 1365
rect 2229 1366 2230 1367
rect 2405 1366 2406 1367
rect 2467 1366 2468 1367
rect 2528 1366 2529 1367
rect 2483 1368 2484 1369
rect 2543 1368 2544 1369
rect 2486 1370 2487 1371
rect 2546 1370 2547 1371
rect 2489 1372 2490 1373
rect 2576 1372 2577 1373
rect 2428 1374 2429 1375
rect 2489 1374 2490 1375
rect 2492 1374 2493 1375
rect 2564 1374 2565 1375
rect 2431 1376 2432 1377
rect 2492 1376 2493 1377
rect 2365 1378 2366 1379
rect 2432 1378 2433 1379
rect 2502 1378 2503 1379
rect 2549 1378 2550 1379
rect 2515 1380 2516 1381
rect 2607 1380 2608 1381
rect 2531 1382 2532 1383
rect 2586 1382 2587 1383
rect 2567 1384 2568 1385
rect 2621 1384 2622 1385
rect 2645 1384 2646 1385
rect 2648 1384 2649 1385
rect 2065 1393 2066 1394
rect 2324 1393 2325 1394
rect 2072 1395 2073 1396
rect 2342 1395 2343 1396
rect 2082 1397 2083 1398
rect 2318 1397 2319 1398
rect 2086 1399 2087 1400
rect 2201 1399 2202 1400
rect 2093 1401 2094 1402
rect 2327 1401 2328 1402
rect 2096 1403 2097 1404
rect 2252 1403 2253 1404
rect 2096 1405 2097 1406
rect 2240 1405 2241 1406
rect 2105 1407 2106 1408
rect 2112 1407 2113 1408
rect 2108 1409 2109 1410
rect 2147 1409 2148 1410
rect 2111 1411 2112 1412
rect 2201 1411 2202 1412
rect 2115 1413 2116 1414
rect 2252 1413 2253 1414
rect 2115 1415 2116 1416
rect 2402 1415 2403 1416
rect 2118 1417 2119 1418
rect 2504 1417 2505 1418
rect 2118 1419 2119 1420
rect 2384 1419 2385 1420
rect 2122 1421 2123 1422
rect 2366 1421 2367 1422
rect 2132 1423 2133 1424
rect 2336 1423 2337 1424
rect 2134 1425 2135 1426
rect 2141 1425 2142 1426
rect 2140 1427 2141 1428
rect 2189 1427 2190 1428
rect 2143 1429 2144 1430
rect 2390 1429 2391 1430
rect 2159 1431 2160 1432
rect 2165 1431 2166 1432
rect 2177 1431 2178 1432
rect 2189 1431 2190 1432
rect 2177 1433 2178 1434
rect 2474 1433 2475 1434
rect 2195 1435 2196 1436
rect 2207 1435 2208 1436
rect 2204 1437 2205 1438
rect 2222 1437 2223 1438
rect 2219 1439 2220 1440
rect 2399 1439 2400 1440
rect 2089 1441 2090 1442
rect 2219 1441 2220 1442
rect 2225 1441 2226 1442
rect 2243 1441 2244 1442
rect 2225 1443 2226 1444
rect 2408 1443 2409 1444
rect 2228 1445 2229 1446
rect 2393 1445 2394 1446
rect 2231 1447 2232 1448
rect 2246 1447 2247 1448
rect 2234 1449 2235 1450
rect 2237 1449 2238 1450
rect 2258 1449 2259 1450
rect 2282 1449 2283 1450
rect 2068 1451 2069 1452
rect 2258 1451 2259 1452
rect 2068 1453 2069 1454
rect 2291 1453 2292 1454
rect 2264 1455 2265 1456
rect 2288 1455 2289 1456
rect 2264 1457 2265 1458
rect 2270 1457 2271 1458
rect 2276 1457 2277 1458
rect 2327 1457 2328 1458
rect 2279 1459 2280 1460
rect 2393 1459 2394 1460
rect 2297 1461 2298 1462
rect 2330 1461 2331 1462
rect 2321 1463 2322 1464
rect 2336 1463 2337 1464
rect 2333 1465 2334 1466
rect 2390 1465 2391 1466
rect 2339 1467 2340 1468
rect 2408 1467 2409 1468
rect 2354 1469 2355 1470
rect 2411 1469 2412 1470
rect 2345 1471 2346 1472
rect 2354 1471 2355 1472
rect 2369 1471 2370 1472
rect 2378 1471 2379 1472
rect 2375 1473 2376 1474
rect 2444 1473 2445 1474
rect 2405 1475 2406 1476
rect 2456 1475 2457 1476
rect 2273 1477 2274 1478
rect 2405 1477 2406 1478
rect 2414 1477 2415 1478
rect 2498 1477 2499 1478
rect 2363 1479 2364 1480
rect 2414 1479 2415 1480
rect 2417 1479 2418 1480
rect 2486 1479 2487 1480
rect 2426 1481 2427 1482
rect 2450 1481 2451 1482
rect 2156 1483 2157 1484
rect 2426 1483 2427 1484
rect 2435 1483 2436 1484
rect 2585 1483 2586 1484
rect 2396 1485 2397 1486
rect 2435 1485 2436 1486
rect 2351 1487 2352 1488
rect 2396 1487 2397 1488
rect 2312 1489 2313 1490
rect 2351 1489 2352 1490
rect 2312 1491 2313 1492
rect 2432 1491 2433 1492
rect 2381 1493 2382 1494
rect 2432 1493 2433 1494
rect 2372 1495 2373 1496
rect 2381 1495 2382 1496
rect 2357 1497 2358 1498
rect 2372 1497 2373 1498
rect 2348 1499 2349 1500
rect 2357 1499 2358 1500
rect 2309 1501 2310 1502
rect 2348 1501 2349 1502
rect 2438 1501 2439 1502
rect 2667 1501 2668 1502
rect 2125 1503 2126 1504
rect 2438 1503 2439 1504
rect 2441 1503 2442 1504
rect 2468 1503 2469 1504
rect 2387 1505 2388 1506
rect 2441 1505 2442 1506
rect 2360 1507 2361 1508
rect 2387 1507 2388 1508
rect 2315 1509 2316 1510
rect 2360 1509 2361 1510
rect 2447 1509 2448 1510
rect 2462 1509 2463 1510
rect 2453 1511 2454 1512
rect 2582 1511 2583 1512
rect 2459 1513 2460 1514
rect 2516 1513 2517 1514
rect 2459 1515 2460 1516
rect 2552 1515 2553 1516
rect 2471 1517 2472 1518
rect 2594 1517 2595 1518
rect 2501 1519 2502 1520
rect 2573 1519 2574 1520
rect 2507 1521 2508 1522
rect 2600 1521 2601 1522
rect 2510 1523 2511 1524
rect 2728 1523 2729 1524
rect 2519 1525 2520 1526
rect 2636 1525 2637 1526
rect 2522 1527 2523 1528
rect 2639 1527 2640 1528
rect 2522 1529 2523 1530
rect 2725 1529 2726 1530
rect 2525 1531 2526 1532
rect 2606 1531 2607 1532
rect 2528 1533 2529 1534
rect 2609 1533 2610 1534
rect 2465 1535 2466 1536
rect 2528 1535 2529 1536
rect 2531 1535 2532 1536
rect 2654 1535 2655 1536
rect 2534 1537 2535 1538
rect 2657 1537 2658 1538
rect 2537 1539 2538 1540
rect 2660 1539 2661 1540
rect 2540 1541 2541 1542
rect 2591 1541 2592 1542
rect 2543 1543 2544 1544
rect 2612 1543 2613 1544
rect 2276 1545 2277 1546
rect 2543 1545 2544 1546
rect 2546 1545 2547 1546
rect 2627 1545 2628 1546
rect 2546 1547 2547 1548
rect 2663 1547 2664 1548
rect 2549 1549 2550 1550
rect 2633 1549 2634 1550
rect 2564 1551 2565 1552
rect 2624 1551 2625 1552
rect 2495 1553 2496 1554
rect 2564 1553 2565 1554
rect 2306 1555 2307 1556
rect 2495 1555 2496 1556
rect 2306 1557 2307 1558
rect 2690 1557 2691 1558
rect 2567 1559 2568 1560
rect 2651 1559 2652 1560
rect 2576 1561 2577 1562
rect 2674 1561 2675 1562
rect 2489 1563 2490 1564
rect 2576 1563 2577 1564
rect 2579 1563 2580 1564
rect 2680 1563 2681 1564
rect 2492 1565 2493 1566
rect 2579 1565 2580 1566
rect 2261 1567 2262 1568
rect 2492 1567 2493 1568
rect 2630 1567 2631 1568
rect 2735 1567 2736 1568
rect 2648 1569 2649 1570
rect 2745 1569 2746 1570
rect 2621 1571 2622 1572
rect 2648 1571 2649 1572
rect 2057 1580 2058 1581
rect 2122 1580 2123 1581
rect 2072 1582 2073 1583
rect 2094 1582 2095 1583
rect 2075 1584 2076 1585
rect 2096 1584 2097 1585
rect 2075 1586 2076 1587
rect 2306 1586 2307 1587
rect 2089 1588 2090 1589
rect 2222 1588 2223 1589
rect 2101 1590 2102 1591
rect 2219 1590 2220 1591
rect 2105 1592 2106 1593
rect 2131 1592 2132 1593
rect 2111 1594 2112 1595
rect 2195 1594 2196 1595
rect 2116 1596 2117 1597
rect 2327 1596 2328 1597
rect 2119 1598 2120 1599
rect 2360 1598 2361 1599
rect 2128 1600 2129 1601
rect 2159 1600 2160 1601
rect 2134 1602 2135 1603
rect 2153 1602 2154 1603
rect 2134 1604 2135 1605
rect 2303 1604 2304 1605
rect 2140 1606 2141 1607
rect 2183 1606 2184 1607
rect 2143 1608 2144 1609
rect 2465 1608 2466 1609
rect 2171 1610 2172 1611
rect 2564 1610 2565 1611
rect 2189 1612 2190 1613
rect 2219 1612 2220 1613
rect 2201 1614 2202 1615
rect 2234 1614 2235 1615
rect 2225 1616 2226 1617
rect 2240 1616 2241 1617
rect 2231 1618 2232 1619
rect 2683 1618 2684 1619
rect 2237 1620 2238 1621
rect 2267 1620 2268 1621
rect 2258 1622 2259 1623
rect 2414 1622 2415 1623
rect 2243 1624 2244 1625
rect 2258 1624 2259 1625
rect 2261 1624 2262 1625
rect 2480 1624 2481 1625
rect 2252 1626 2253 1627
rect 2261 1626 2262 1627
rect 2246 1628 2247 1629
rect 2252 1628 2253 1629
rect 2264 1628 2265 1629
rect 2273 1628 2274 1629
rect 2276 1628 2277 1629
rect 2639 1628 2640 1629
rect 2282 1630 2283 1631
rect 2291 1630 2292 1631
rect 2285 1632 2286 1633
rect 2357 1632 2358 1633
rect 2288 1634 2289 1635
rect 2297 1634 2298 1635
rect 2315 1634 2316 1635
rect 2704 1634 2705 1635
rect 2318 1636 2319 1637
rect 2321 1636 2322 1637
rect 2324 1636 2325 1637
rect 2327 1636 2328 1637
rect 2351 1636 2352 1637
rect 2369 1636 2370 1637
rect 2098 1638 2099 1639
rect 2351 1638 2352 1639
rect 2363 1638 2364 1639
rect 2504 1638 2505 1639
rect 2396 1640 2397 1641
rect 2414 1640 2415 1641
rect 2396 1642 2397 1643
rect 2402 1642 2403 1643
rect 2390 1644 2391 1645
rect 2402 1644 2403 1645
rect 2384 1646 2385 1647
rect 2390 1646 2391 1647
rect 2372 1648 2373 1649
rect 2384 1648 2385 1649
rect 2366 1650 2367 1651
rect 2372 1650 2373 1651
rect 2082 1652 2083 1653
rect 2366 1652 2367 1653
rect 2068 1654 2069 1655
rect 2081 1654 2082 1655
rect 2068 1656 2069 1657
rect 2165 1656 2166 1657
rect 2399 1656 2400 1657
rect 2405 1656 2406 1657
rect 2393 1658 2394 1659
rect 2405 1658 2406 1659
rect 2387 1660 2388 1661
rect 2393 1660 2394 1661
rect 2408 1660 2409 1661
rect 2420 1660 2421 1661
rect 2408 1662 2409 1663
rect 2426 1662 2427 1663
rect 2411 1664 2412 1665
rect 2423 1664 2424 1665
rect 2432 1664 2433 1665
rect 2552 1664 2553 1665
rect 2432 1666 2433 1667
rect 2441 1666 2442 1667
rect 2435 1668 2436 1669
rect 2555 1668 2556 1669
rect 2459 1670 2460 1671
rect 2489 1670 2490 1671
rect 2462 1672 2463 1673
rect 2726 1672 2727 1673
rect 2438 1674 2439 1675
rect 2462 1674 2463 1675
rect 2438 1676 2439 1677
rect 2670 1676 2671 1677
rect 2468 1678 2469 1679
rect 2667 1678 2668 1679
rect 2456 1680 2457 1681
rect 2468 1680 2469 1681
rect 2456 1682 2457 1683
rect 2669 1682 2670 1683
rect 2474 1684 2475 1685
rect 2588 1684 2589 1685
rect 2150 1686 2151 1687
rect 2474 1686 2475 1687
rect 2486 1686 2487 1687
rect 2531 1686 2532 1687
rect 2444 1688 2445 1689
rect 2486 1688 2487 1689
rect 2162 1690 2163 1691
rect 2444 1690 2445 1691
rect 2492 1690 2493 1691
rect 2558 1690 2559 1691
rect 2495 1692 2496 1693
rect 2561 1692 2562 1693
rect 2504 1694 2505 1695
rect 2510 1694 2511 1695
rect 2501 1696 2502 1697
rect 2510 1696 2511 1697
rect 2516 1696 2517 1697
rect 2525 1696 2526 1697
rect 2498 1698 2499 1699
rect 2516 1698 2517 1699
rect 2519 1698 2520 1699
rect 2784 1698 2785 1699
rect 2522 1700 2523 1701
rect 2537 1700 2538 1701
rect 2543 1700 2544 1701
rect 2570 1700 2571 1701
rect 2543 1702 2544 1703
rect 2609 1702 2610 1703
rect 2546 1704 2547 1705
rect 2591 1704 2592 1705
rect 2528 1706 2529 1707
rect 2546 1706 2547 1707
rect 2564 1706 2565 1707
rect 2791 1706 2792 1707
rect 2582 1708 2583 1709
rect 2666 1708 2667 1709
rect 2582 1710 2583 1711
rect 2674 1710 2675 1711
rect 2585 1712 2586 1713
rect 2663 1712 2664 1713
rect 2594 1714 2595 1715
rect 2684 1714 2685 1715
rect 2540 1716 2541 1717
rect 2594 1716 2595 1717
rect 2600 1716 2601 1717
rect 2711 1716 2712 1717
rect 2579 1718 2580 1719
rect 2600 1718 2601 1719
rect 2606 1718 2607 1719
rect 2697 1718 2698 1719
rect 2624 1720 2625 1721
rect 2794 1720 2795 1721
rect 2627 1722 2628 1723
rect 2675 1722 2676 1723
rect 2576 1724 2577 1725
rect 2627 1724 2628 1725
rect 2360 1726 2361 1727
rect 2576 1726 2577 1727
rect 2630 1726 2631 1727
rect 2787 1726 2788 1727
rect 2633 1728 2634 1729
rect 2678 1728 2679 1729
rect 2636 1730 2637 1731
rect 2708 1730 2709 1731
rect 2636 1732 2637 1733
rect 2766 1732 2767 1733
rect 2639 1734 2640 1735
rect 2763 1734 2764 1735
rect 2642 1736 2643 1737
rect 2756 1736 2757 1737
rect 2648 1738 2649 1739
rect 2696 1738 2697 1739
rect 2651 1740 2652 1741
rect 2699 1740 2700 1741
rect 2654 1742 2655 1743
rect 2720 1742 2721 1743
rect 2612 1744 2613 1745
rect 2654 1744 2655 1745
rect 2657 1744 2658 1745
rect 2723 1744 2724 1745
rect 2312 1746 2313 1747
rect 2657 1746 2658 1747
rect 2159 1748 2160 1749
rect 2312 1748 2313 1749
rect 2660 1748 2661 1749
rect 2714 1748 2715 1749
rect 2279 1750 2280 1751
rect 2660 1750 2661 1751
rect 2137 1752 2138 1753
rect 2279 1752 2280 1753
rect 2680 1752 2681 1753
rect 2739 1752 2740 1753
rect 2681 1754 2682 1755
rect 2718 1754 2719 1755
rect 2513 1756 2514 1757
rect 2717 1756 2718 1757
rect 2745 1756 2746 1757
rect 2818 1756 2819 1757
rect 2808 1758 2809 1759
rect 2812 1758 2813 1759
rect 2047 1767 2048 1768
rect 2122 1767 2123 1768
rect 2054 1769 2055 1770
rect 2075 1769 2076 1770
rect 2059 1771 2060 1772
rect 2075 1771 2076 1772
rect 2061 1773 2062 1774
rect 2081 1773 2082 1774
rect 2071 1775 2072 1776
rect 2454 1775 2455 1776
rect 2064 1777 2065 1778
rect 2072 1777 2073 1778
rect 2078 1777 2079 1778
rect 2165 1777 2166 1778
rect 2087 1779 2088 1780
rect 2348 1779 2349 1780
rect 2089 1781 2090 1782
rect 2234 1781 2235 1782
rect 2082 1783 2083 1784
rect 2235 1783 2236 1784
rect 2092 1785 2093 1786
rect 2376 1785 2377 1786
rect 2113 1787 2114 1788
rect 2354 1787 2355 1788
rect 2116 1789 2117 1790
rect 2384 1789 2385 1790
rect 2119 1791 2120 1792
rect 2390 1791 2391 1792
rect 2119 1793 2120 1794
rect 2131 1793 2132 1794
rect 2125 1795 2126 1796
rect 2423 1795 2424 1796
rect 2128 1797 2129 1798
rect 2460 1797 2461 1798
rect 2129 1799 2130 1800
rect 2153 1799 2154 1800
rect 2134 1801 2135 1802
rect 2256 1801 2257 1802
rect 2137 1803 2138 1804
rect 2273 1803 2274 1804
rect 2144 1805 2145 1806
rect 2444 1805 2445 1806
rect 2125 1807 2126 1808
rect 2144 1807 2145 1808
rect 2148 1807 2149 1808
rect 2499 1807 2500 1808
rect 2171 1809 2172 1810
rect 2378 1809 2379 1810
rect 2174 1811 2175 1812
rect 2279 1811 2280 1812
rect 2181 1813 2182 1814
rect 2489 1813 2490 1814
rect 2202 1815 2203 1816
rect 2231 1815 2232 1816
rect 2205 1817 2206 1818
rect 2219 1817 2220 1818
rect 2207 1819 2208 1820
rect 2486 1819 2487 1820
rect 2210 1821 2211 1822
rect 2673 1821 2674 1822
rect 2223 1823 2224 1824
rect 2252 1823 2253 1824
rect 2229 1825 2230 1826
rect 2393 1825 2394 1826
rect 2240 1827 2241 1828
rect 2472 1827 2473 1828
rect 2241 1829 2242 1830
rect 2258 1829 2259 1830
rect 2244 1831 2245 1832
rect 2309 1831 2310 1832
rect 2250 1833 2251 1834
rect 2267 1833 2268 1834
rect 2268 1835 2269 1836
rect 2291 1835 2292 1836
rect 2274 1837 2275 1838
rect 2297 1837 2298 1838
rect 2280 1839 2281 1840
rect 2303 1839 2304 1840
rect 2289 1841 2290 1842
rect 2627 1841 2628 1842
rect 2292 1843 2293 1844
rect 2315 1843 2316 1844
rect 2310 1845 2311 1846
rect 2321 1845 2322 1846
rect 2312 1847 2313 1848
rect 2715 1847 2716 1848
rect 2316 1849 2317 1850
rect 2330 1849 2331 1850
rect 2322 1851 2323 1852
rect 2372 1851 2373 1852
rect 2327 1853 2328 1854
rect 2391 1853 2392 1854
rect 2328 1855 2329 1856
rect 2402 1855 2403 1856
rect 2151 1857 2152 1858
rect 2403 1857 2404 1858
rect 2331 1859 2332 1860
rect 2405 1859 2406 1860
rect 2334 1861 2335 1862
rect 2570 1861 2571 1862
rect 2346 1863 2347 1864
rect 2438 1863 2439 1864
rect 2351 1865 2352 1866
rect 2436 1865 2437 1866
rect 2352 1867 2353 1868
rect 2552 1867 2553 1868
rect 2355 1869 2356 1870
rect 2555 1869 2556 1870
rect 2360 1871 2361 1872
rect 2588 1871 2589 1872
rect 2363 1873 2364 1874
rect 2594 1873 2595 1874
rect 2364 1875 2365 1876
rect 2561 1875 2562 1876
rect 2379 1877 2380 1878
rect 2657 1877 2658 1878
rect 2385 1879 2386 1880
rect 2462 1879 2463 1880
rect 2366 1881 2367 1882
rect 2463 1881 2464 1882
rect 2396 1883 2397 1884
rect 2487 1883 2488 1884
rect 2101 1885 2102 1886
rect 2397 1885 2398 1886
rect 2399 1885 2400 1886
rect 2490 1885 2491 1886
rect 2381 1887 2382 1888
rect 2400 1887 2401 1888
rect 2420 1887 2421 1888
rect 2445 1887 2446 1888
rect 2068 1889 2069 1890
rect 2421 1889 2422 1890
rect 2069 1891 2070 1892
rect 2319 1891 2320 1892
rect 2427 1891 2428 1892
rect 2808 1891 2809 1892
rect 2432 1893 2433 1894
rect 2493 1893 2494 1894
rect 2342 1895 2343 1896
rect 2433 1895 2434 1896
rect 2439 1895 2440 1896
rect 2468 1895 2469 1896
rect 2098 1897 2099 1898
rect 2469 1897 2470 1898
rect 2465 1899 2466 1900
rect 2508 1899 2509 1900
rect 2369 1901 2370 1902
rect 2466 1901 2467 1902
rect 2370 1903 2371 1904
rect 2531 1903 2532 1904
rect 2474 1905 2475 1906
rect 2733 1905 2734 1906
rect 2475 1907 2476 1908
rect 2564 1907 2565 1908
rect 2484 1909 2485 1910
rect 2558 1909 2559 1910
rect 2504 1911 2505 1912
rect 2589 1911 2590 1912
rect 2408 1913 2409 1914
rect 2505 1913 2506 1914
rect 2159 1915 2160 1916
rect 2409 1915 2410 1916
rect 2160 1917 2161 1918
rect 2183 1917 2184 1918
rect 2510 1917 2511 1918
rect 2586 1917 2587 1918
rect 2511 1919 2512 1920
rect 2729 1919 2730 1920
rect 2516 1921 2517 1922
rect 2541 1921 2542 1922
rect 2141 1923 2142 1924
rect 2517 1923 2518 1924
rect 2141 1925 2142 1926
rect 2298 1925 2299 1926
rect 2523 1925 2524 1926
rect 2546 1925 2547 1926
rect 2525 1927 2526 1928
rect 2553 1927 2554 1928
rect 2529 1929 2530 1930
rect 2537 1929 2538 1930
rect 2547 1929 2548 1930
rect 2642 1929 2643 1930
rect 2550 1931 2551 1932
rect 2660 1931 2661 1932
rect 2559 1933 2560 1934
rect 2582 1933 2583 1934
rect 2571 1935 2572 1936
rect 2749 1935 2750 1936
rect 2580 1937 2581 1938
rect 2775 1937 2776 1938
rect 2613 1939 2614 1940
rect 2663 1939 2664 1940
rect 2616 1941 2617 1942
rect 2666 1941 2667 1942
rect 2619 1943 2620 1944
rect 2850 1943 2851 1944
rect 2624 1945 2625 1946
rect 2634 1945 2635 1946
rect 2628 1947 2629 1948
rect 2723 1947 2724 1948
rect 2636 1949 2637 1950
rect 2661 1949 2662 1950
rect 2600 1951 2601 1952
rect 2637 1951 2638 1952
rect 2519 1953 2520 1954
rect 2601 1953 2602 1954
rect 2639 1953 2640 1954
rect 2649 1953 2650 1954
rect 2640 1955 2641 1956
rect 2839 1955 2840 1956
rect 2667 1957 2668 1958
rect 2763 1957 2764 1958
rect 2576 1959 2577 1960
rect 2763 1959 2764 1960
rect 2543 1961 2544 1962
rect 2577 1961 2578 1962
rect 2513 1963 2514 1964
rect 2544 1963 2545 1964
rect 2675 1963 2676 1964
rect 2703 1963 2704 1964
rect 2678 1965 2679 1966
rect 2724 1965 2725 1966
rect 2654 1967 2655 1968
rect 2679 1967 2680 1968
rect 2681 1967 2682 1968
rect 2752 1967 2753 1968
rect 2682 1969 2683 1970
rect 2843 1969 2844 1970
rect 2696 1971 2697 1972
rect 2760 1971 2761 1972
rect 2697 1973 2698 1974
rect 2708 1973 2709 1974
rect 2699 1975 2700 1976
rect 2727 1975 2728 1976
rect 2700 1977 2701 1978
rect 2711 1977 2712 1978
rect 2706 1979 2707 1980
rect 2791 1979 2792 1980
rect 2720 1981 2721 1982
rect 2784 1981 2785 1982
rect 2736 1983 2737 1984
rect 2742 1983 2743 1984
rect 2739 1985 2740 1986
rect 2769 1985 2770 1986
rect 2739 1987 2740 1988
rect 2801 1987 2802 1988
rect 2742 1989 2743 1990
rect 2766 1989 2767 1990
rect 2450 1991 2451 1992
rect 2766 1991 2767 1992
rect 2084 1993 2085 1994
rect 2451 1993 2452 1994
rect 2085 1995 2086 1996
rect 2261 1995 2262 1996
rect 2262 1997 2263 1998
rect 2285 1997 2286 1998
rect 2286 1999 2287 2000
rect 2456 1999 2457 2000
rect 2414 2001 2415 2002
rect 2457 2001 2458 2002
rect 2336 2003 2337 2004
rect 2415 2003 2416 2004
rect 2757 2003 2758 2004
rect 2829 2003 2830 2004
rect 2772 2005 2773 2006
rect 2778 2005 2779 2006
rect 2781 2005 2782 2006
rect 2790 2005 2791 2006
rect 2797 2005 2798 2006
rect 2808 2005 2809 2006
rect 2812 2005 2813 2006
rect 2821 2005 2822 2006
rect 2811 2007 2812 2008
rect 2825 2007 2826 2008
rect 2818 2009 2819 2010
rect 2856 2009 2857 2010
rect 2721 2011 2722 2012
rect 2818 2011 2819 2012
rect 2822 2011 2823 2012
rect 2846 2011 2847 2012
rect 2011 2020 2012 2021
rect 2447 2020 2448 2021
rect 2066 2022 2067 2023
rect 2463 2022 2464 2023
rect 2069 2024 2070 2025
rect 2451 2024 2452 2025
rect 2072 2026 2073 2027
rect 2381 2026 2382 2027
rect 2078 2028 2079 2029
rect 2171 2028 2172 2029
rect 2092 2030 2093 2031
rect 2122 2030 2123 2031
rect 2104 2032 2105 2033
rect 2160 2032 2161 2033
rect 2110 2034 2111 2035
rect 2436 2034 2437 2035
rect 2113 2036 2114 2037
rect 2409 2036 2410 2037
rect 2119 2038 2120 2039
rect 2135 2038 2136 2039
rect 2129 2040 2130 2041
rect 2490 2040 2491 2041
rect 2141 2042 2142 2043
rect 2501 2042 2502 2043
rect 2141 2044 2142 2045
rect 2415 2044 2416 2045
rect 2144 2046 2145 2047
rect 2439 2046 2440 2047
rect 2148 2048 2149 2049
rect 2385 2048 2386 2049
rect 2148 2050 2149 2051
rect 2229 2050 2230 2051
rect 2152 2052 2153 2053
rect 2310 2052 2311 2053
rect 2155 2054 2156 2055
rect 2493 2054 2494 2055
rect 2159 2056 2160 2057
rect 2489 2056 2490 2057
rect 2178 2058 2179 2059
rect 2207 2058 2208 2059
rect 2075 2060 2076 2061
rect 2177 2060 2178 2061
rect 2181 2060 2182 2061
rect 2492 2060 2493 2061
rect 2190 2062 2191 2063
rect 2715 2062 2716 2063
rect 2202 2064 2203 2065
rect 2450 2064 2451 2065
rect 2205 2066 2206 2067
rect 2231 2066 2232 2067
rect 2243 2068 2244 2069
rect 2472 2068 2473 2069
rect 2256 2070 2257 2071
rect 2324 2070 2325 2071
rect 2219 2072 2220 2073
rect 2255 2072 2256 2073
rect 2262 2072 2263 2073
rect 2306 2072 2307 2073
rect 2264 2074 2265 2075
rect 2603 2074 2604 2075
rect 2268 2076 2269 2077
rect 2312 2076 2313 2077
rect 2082 2078 2083 2079
rect 2267 2078 2268 2079
rect 2276 2078 2277 2079
rect 2466 2078 2467 2079
rect 2280 2080 2281 2081
rect 2849 2080 2850 2081
rect 2250 2082 2251 2083
rect 2279 2082 2280 2083
rect 2289 2082 2290 2083
rect 2697 2082 2698 2083
rect 2292 2084 2293 2085
rect 2342 2084 2343 2085
rect 2241 2086 2242 2087
rect 2291 2086 2292 2087
rect 2298 2086 2299 2087
rect 2348 2086 2349 2087
rect 2316 2088 2317 2089
rect 2360 2088 2361 2089
rect 2322 2090 2323 2091
rect 2366 2090 2367 2091
rect 2328 2092 2329 2093
rect 2372 2092 2373 2093
rect 2346 2094 2347 2095
rect 2384 2094 2385 2095
rect 2352 2096 2353 2097
rect 2408 2096 2409 2097
rect 2364 2098 2365 2099
rect 2414 2098 2415 2099
rect 2319 2100 2320 2101
rect 2363 2100 2364 2101
rect 2274 2102 2275 2103
rect 2318 2102 2319 2103
rect 2235 2104 2236 2105
rect 2273 2104 2274 2105
rect 2370 2104 2371 2105
rect 2429 2104 2430 2105
rect 2397 2106 2398 2107
rect 2465 2106 2466 2107
rect 2379 2108 2380 2109
rect 2396 2108 2397 2109
rect 2059 2110 2060 2111
rect 2378 2110 2379 2111
rect 2427 2110 2428 2111
rect 2471 2110 2472 2111
rect 2376 2112 2377 2113
rect 2426 2112 2427 2113
rect 2331 2114 2332 2115
rect 2375 2114 2376 2115
rect 2125 2116 2126 2117
rect 2330 2116 2331 2117
rect 2125 2118 2126 2119
rect 2195 2118 2196 2119
rect 2433 2118 2434 2119
rect 2495 2118 2496 2119
rect 2445 2120 2446 2121
rect 2519 2120 2520 2121
rect 2444 2122 2445 2123
rect 2484 2122 2485 2123
rect 2421 2124 2422 2125
rect 2483 2124 2484 2125
rect 2193 2126 2194 2127
rect 2420 2126 2421 2127
rect 2457 2126 2458 2127
rect 2525 2126 2526 2127
rect 2469 2128 2470 2129
rect 2477 2128 2478 2129
rect 2475 2130 2476 2131
rect 2513 2130 2514 2131
rect 2481 2132 2482 2133
rect 2531 2132 2532 2133
rect 2499 2134 2500 2135
rect 2537 2134 2538 2135
rect 2076 2136 2077 2137
rect 2498 2136 2499 2137
rect 2505 2136 2506 2137
rect 2561 2136 2562 2137
rect 2400 2138 2401 2139
rect 2504 2138 2505 2139
rect 2508 2138 2509 2139
rect 2564 2138 2565 2139
rect 2116 2140 2117 2141
rect 2507 2140 2508 2141
rect 2511 2140 2512 2141
rect 2789 2140 2790 2141
rect 2355 2142 2356 2143
rect 2510 2142 2511 2143
rect 2334 2144 2335 2145
rect 2354 2144 2355 2145
rect 2517 2144 2518 2145
rect 2852 2144 2853 2145
rect 2523 2146 2524 2147
rect 2573 2146 2574 2147
rect 2541 2148 2542 2149
rect 2597 2148 2598 2149
rect 2544 2150 2545 2151
rect 2801 2150 2802 2151
rect 2487 2152 2488 2153
rect 2543 2152 2544 2153
rect 2069 2154 2070 2155
rect 2486 2154 2487 2155
rect 2547 2154 2548 2155
rect 2567 2154 2568 2155
rect 2286 2156 2287 2157
rect 2546 2156 2547 2157
rect 2555 2156 2556 2157
rect 2559 2156 2560 2157
rect 2586 2156 2587 2157
rect 2642 2156 2643 2157
rect 2261 2158 2262 2159
rect 2585 2158 2586 2159
rect 2609 2158 2610 2159
rect 2775 2158 2776 2159
rect 2619 2160 2620 2161
rect 2832 2160 2833 2161
rect 2621 2162 2622 2163
rect 2772 2162 2773 2163
rect 2640 2164 2641 2165
rect 2708 2164 2709 2165
rect 2577 2166 2578 2167
rect 2639 2166 2640 2167
rect 2649 2166 2650 2167
rect 2750 2166 2751 2167
rect 2589 2168 2590 2169
rect 2648 2168 2649 2169
rect 2247 2170 2248 2171
rect 2588 2170 2589 2171
rect 2667 2170 2668 2171
rect 2762 2170 2763 2171
rect 2637 2172 2638 2173
rect 2666 2172 2667 2173
rect 2673 2172 2674 2173
rect 2865 2172 2866 2173
rect 2672 2174 2673 2175
rect 2942 2174 2943 2175
rect 2676 2176 2677 2177
rect 2706 2176 2707 2177
rect 2682 2178 2683 2179
rect 2771 2178 2772 2179
rect 2685 2180 2686 2181
rect 2859 2180 2860 2181
rect 2628 2182 2629 2183
rect 2684 2182 2685 2183
rect 2571 2184 2572 2185
rect 2627 2184 2628 2185
rect 2550 2186 2551 2187
rect 2570 2186 2571 2187
rect 2690 2186 2691 2187
rect 2907 2186 2908 2187
rect 2693 2188 2694 2189
rect 2889 2188 2890 2189
rect 2696 2190 2697 2191
rect 2900 2190 2901 2191
rect 2703 2192 2704 2193
rect 2804 2192 2805 2193
rect 2711 2194 2712 2195
rect 2754 2194 2755 2195
rect 2718 2196 2719 2197
rect 2798 2196 2799 2197
rect 2721 2198 2722 2199
rect 2819 2198 2820 2199
rect 2724 2200 2725 2201
rect 2822 2200 2823 2201
rect 2729 2202 2730 2203
rect 2935 2202 2936 2203
rect 2739 2204 2740 2205
rect 2837 2204 2838 2205
rect 2616 2206 2617 2207
rect 2738 2206 2739 2207
rect 2553 2208 2554 2209
rect 2615 2208 2616 2209
rect 2742 2208 2743 2209
rect 2840 2208 2841 2209
rect 2747 2210 2748 2211
rect 2954 2210 2955 2211
rect 2757 2212 2758 2213
rect 2825 2212 2826 2213
rect 2661 2214 2662 2215
rect 2756 2214 2757 2215
rect 2601 2216 2602 2217
rect 2660 2216 2661 2217
rect 2727 2216 2728 2217
rect 2825 2216 2826 2217
rect 2760 2218 2761 2219
rect 2877 2218 2878 2219
rect 2766 2220 2767 2221
rect 2896 2220 2897 2221
rect 2769 2222 2770 2223
rect 2862 2222 2863 2223
rect 2679 2224 2680 2225
rect 2768 2224 2769 2225
rect 2781 2224 2782 2225
rect 2880 2224 2881 2225
rect 2613 2226 2614 2227
rect 2780 2226 2781 2227
rect 2784 2226 2785 2227
rect 2883 2226 2884 2227
rect 2735 2228 2736 2229
rect 2783 2228 2784 2229
rect 2787 2228 2788 2229
rect 2794 2228 2795 2229
rect 2634 2230 2635 2231
rect 2795 2230 2796 2231
rect 2580 2232 2581 2233
rect 2633 2232 2634 2233
rect 2529 2234 2530 2235
rect 2579 2234 2580 2235
rect 2460 2236 2461 2237
rect 2528 2236 2529 2237
rect 2391 2238 2392 2239
rect 2459 2238 2460 2239
rect 2390 2240 2391 2241
rect 2454 2240 2455 2241
rect 2403 2242 2404 2243
rect 2453 2242 2454 2243
rect 2145 2244 2146 2245
rect 2402 2244 2403 2245
rect 2700 2244 2701 2245
rect 2786 2244 2787 2245
rect 2792 2244 2793 2245
rect 2868 2244 2869 2245
rect 2856 2246 2857 2247
rect 2948 2246 2949 2247
rect 2702 2248 2703 2249
rect 2856 2248 2857 2249
rect 2874 2248 2875 2249
rect 2921 2248 2922 2249
rect 2045 2257 2046 2258
rect 2049 2257 2050 2258
rect 2062 2257 2063 2258
rect 2483 2257 2484 2258
rect 2066 2259 2067 2260
rect 2390 2259 2391 2260
rect 2070 2261 2071 2262
rect 2486 2261 2487 2262
rect 2080 2263 2081 2264
rect 2110 2263 2111 2264
rect 2088 2265 2089 2266
rect 2229 2265 2230 2266
rect 2089 2267 2090 2268
rect 2498 2267 2499 2268
rect 2097 2269 2098 2270
rect 2400 2269 2401 2270
rect 2098 2271 2099 2272
rect 2322 2271 2323 2272
rect 2107 2273 2108 2274
rect 2171 2273 2172 2274
rect 2107 2275 2108 2276
rect 2231 2275 2232 2276
rect 2117 2277 2118 2278
rect 2418 2277 2419 2278
rect 2125 2279 2126 2280
rect 2363 2279 2364 2280
rect 2126 2281 2127 2282
rect 2366 2281 2367 2282
rect 2129 2283 2130 2284
rect 2525 2283 2526 2284
rect 2138 2285 2139 2286
rect 2154 2285 2155 2286
rect 2141 2287 2142 2288
rect 2465 2287 2466 2288
rect 2143 2289 2144 2290
rect 2495 2289 2496 2290
rect 2157 2291 2158 2292
rect 2469 2291 2470 2292
rect 2159 2293 2160 2294
rect 2288 2293 2289 2294
rect 2135 2295 2136 2296
rect 2160 2295 2161 2296
rect 2162 2295 2163 2296
rect 2477 2295 2478 2296
rect 2152 2297 2153 2298
rect 2163 2297 2164 2298
rect 2177 2297 2178 2298
rect 2193 2297 2194 2298
rect 2187 2299 2188 2300
rect 2564 2299 2565 2300
rect 2195 2301 2196 2302
rect 2211 2301 2212 2302
rect 2199 2303 2200 2304
rect 2207 2303 2208 2304
rect 2217 2303 2218 2304
rect 2528 2303 2529 2304
rect 2219 2305 2220 2306
rect 2510 2305 2511 2306
rect 2222 2307 2223 2308
rect 2607 2307 2608 2308
rect 2243 2309 2244 2310
rect 2289 2309 2290 2310
rect 2250 2311 2251 2312
rect 2496 2311 2497 2312
rect 2255 2313 2256 2314
rect 2346 2313 2347 2314
rect 2259 2315 2260 2316
rect 2279 2315 2280 2316
rect 2267 2317 2268 2318
rect 2271 2317 2272 2318
rect 2276 2317 2277 2318
rect 2280 2317 2281 2318
rect 2273 2319 2274 2320
rect 2277 2319 2278 2320
rect 2291 2319 2292 2320
rect 2295 2319 2296 2320
rect 2304 2319 2305 2320
rect 2312 2319 2313 2320
rect 2076 2321 2077 2322
rect 2313 2321 2314 2322
rect 2306 2323 2307 2324
rect 2310 2323 2311 2324
rect 2316 2323 2317 2324
rect 2318 2323 2319 2324
rect 2324 2323 2325 2324
rect 2328 2323 2329 2324
rect 2330 2323 2331 2324
rect 2334 2323 2335 2324
rect 2340 2323 2341 2324
rect 2342 2323 2343 2324
rect 2348 2323 2349 2324
rect 2364 2323 2365 2324
rect 2352 2325 2353 2326
rect 2447 2325 2448 2326
rect 2166 2327 2167 2328
rect 2448 2327 2449 2328
rect 2358 2329 2359 2330
rect 2378 2329 2379 2330
rect 2360 2331 2361 2332
rect 2370 2331 2371 2332
rect 2361 2333 2362 2334
rect 2381 2333 2382 2334
rect 2372 2335 2373 2336
rect 2394 2335 2395 2336
rect 2122 2337 2123 2338
rect 2373 2337 2374 2338
rect 2382 2337 2383 2338
rect 2459 2337 2460 2338
rect 2148 2339 2149 2340
rect 2460 2339 2461 2340
rect 2147 2341 2148 2342
rect 2265 2341 2266 2342
rect 2391 2341 2392 2342
rect 2426 2341 2427 2342
rect 2247 2343 2248 2344
rect 2427 2343 2428 2344
rect 2402 2345 2403 2346
rect 2478 2345 2479 2346
rect 2406 2347 2407 2348
rect 2501 2347 2502 2348
rect 2412 2349 2413 2350
rect 2745 2349 2746 2350
rect 2424 2351 2425 2352
rect 2519 2351 2520 2352
rect 2429 2353 2430 2354
rect 2592 2353 2593 2354
rect 2436 2355 2437 2356
rect 2453 2355 2454 2356
rect 2442 2357 2443 2358
rect 2543 2357 2544 2358
rect 2136 2359 2137 2360
rect 2544 2359 2545 2360
rect 2454 2361 2455 2362
rect 2561 2361 2562 2362
rect 2466 2363 2467 2364
rect 2871 2363 2872 2364
rect 2475 2365 2476 2366
rect 2492 2365 2493 2366
rect 2484 2367 2485 2368
rect 2585 2367 2586 2368
rect 2502 2369 2503 2370
rect 2507 2369 2508 2370
rect 2420 2371 2421 2372
rect 2508 2371 2509 2372
rect 2421 2373 2422 2374
rect 2504 2373 2505 2374
rect 2520 2373 2521 2374
rect 2573 2373 2574 2374
rect 2526 2375 2527 2376
rect 2889 2375 2890 2376
rect 2550 2377 2551 2378
rect 2648 2377 2649 2378
rect 2574 2379 2575 2380
rect 2945 2379 2946 2380
rect 2609 2381 2610 2382
rect 2655 2381 2656 2382
rect 2619 2383 2620 2384
rect 2693 2383 2694 2384
rect 2621 2385 2622 2386
rect 2649 2385 2650 2386
rect 2627 2387 2628 2388
rect 2903 2387 2904 2388
rect 2628 2389 2629 2390
rect 2708 2389 2709 2390
rect 2537 2391 2538 2392
rect 2709 2391 2710 2392
rect 2414 2393 2415 2394
rect 2538 2393 2539 2394
rect 2415 2395 2416 2396
rect 2622 2395 2623 2396
rect 2631 2395 2632 2396
rect 2633 2395 2634 2396
rect 2637 2395 2638 2396
rect 2702 2395 2703 2396
rect 2555 2397 2556 2398
rect 2703 2397 2704 2398
rect 2556 2399 2557 2400
rect 2642 2399 2643 2400
rect 2639 2401 2640 2402
rect 2844 2401 2845 2402
rect 2679 2403 2680 2404
rect 2747 2403 2748 2404
rect 2588 2405 2589 2406
rect 2748 2405 2749 2406
rect 2684 2407 2685 2408
rect 2900 2407 2901 2408
rect 2471 2409 2472 2410
rect 2685 2409 2686 2410
rect 2472 2411 2473 2412
rect 2489 2411 2490 2412
rect 2490 2413 2491 2414
rect 2531 2413 2532 2414
rect 2532 2415 2533 2416
rect 2579 2415 2580 2416
rect 2580 2417 2581 2418
rect 2660 2417 2661 2418
rect 2444 2419 2445 2420
rect 2661 2419 2662 2420
rect 2445 2421 2446 2422
rect 2546 2421 2547 2422
rect 2696 2421 2697 2422
rect 2935 2421 2936 2422
rect 2697 2423 2698 2424
rect 2958 2423 2959 2424
rect 2241 2425 2242 2426
rect 2959 2425 2960 2426
rect 2700 2427 2701 2428
rect 2966 2427 2967 2428
rect 2715 2429 2716 2430
rect 2914 2429 2915 2430
rect 2729 2431 2730 2432
rect 2733 2431 2734 2432
rect 2735 2431 2736 2432
rect 2829 2431 2830 2432
rect 2738 2433 2739 2434
rect 2832 2433 2833 2434
rect 2750 2435 2751 2436
rect 2931 2435 2932 2436
rect 2396 2437 2397 2438
rect 2751 2437 2752 2438
rect 2375 2439 2376 2440
rect 2397 2439 2398 2440
rect 2100 2441 2101 2442
rect 2376 2441 2377 2442
rect 2756 2441 2757 2442
rect 2938 2441 2939 2442
rect 2757 2443 2758 2444
rect 2762 2443 2763 2444
rect 2666 2445 2667 2446
rect 2763 2445 2764 2446
rect 2667 2447 2668 2448
rect 2945 2447 2946 2448
rect 2760 2449 2761 2450
rect 2795 2449 2796 2450
rect 2771 2451 2772 2452
rect 2775 2451 2776 2452
rect 2768 2453 2769 2454
rect 2772 2453 2773 2454
rect 2784 2453 2785 2454
rect 2813 2453 2814 2454
rect 2786 2455 2787 2456
rect 2847 2455 2848 2456
rect 2597 2457 2598 2458
rect 2787 2457 2788 2458
rect 2513 2459 2514 2460
rect 2598 2459 2599 2460
rect 2789 2459 2790 2460
rect 2850 2459 2851 2460
rect 2570 2461 2571 2462
rect 2790 2461 2791 2462
rect 2796 2461 2797 2462
rect 2804 2461 2805 2462
rect 2567 2463 2568 2464
rect 2805 2463 2806 2464
rect 2568 2465 2569 2466
rect 2672 2465 2673 2466
rect 2673 2467 2674 2468
rect 2711 2467 2712 2468
rect 2798 2467 2799 2468
rect 2870 2467 2871 2468
rect 2801 2469 2802 2470
rect 2816 2469 2817 2470
rect 2811 2471 2812 2472
rect 2819 2471 2820 2472
rect 2814 2473 2815 2474
rect 2822 2473 2823 2474
rect 2817 2475 2818 2476
rect 2825 2475 2826 2476
rect 2823 2477 2824 2478
rect 2877 2477 2878 2478
rect 2837 2479 2838 2480
rect 2891 2479 2892 2480
rect 2840 2481 2841 2482
rect 2868 2481 2869 2482
rect 2792 2483 2793 2484
rect 2867 2483 2868 2484
rect 2354 2485 2355 2486
rect 2793 2485 2794 2486
rect 2355 2487 2356 2488
rect 2450 2487 2451 2488
rect 2841 2487 2842 2488
rect 2893 2487 2894 2488
rect 2852 2489 2853 2490
rect 2856 2489 2857 2490
rect 2603 2491 2604 2492
rect 2856 2491 2857 2492
rect 2408 2493 2409 2494
rect 2604 2493 2605 2494
rect 2865 2493 2866 2494
rect 2888 2493 2889 2494
rect 2874 2495 2875 2496
rect 2918 2495 2919 2496
rect 2873 2497 2874 2498
rect 2952 2497 2953 2498
rect 2880 2499 2881 2500
rect 2897 2499 2898 2500
rect 2879 2501 2880 2502
rect 2938 2501 2939 2502
rect 2883 2503 2884 2504
rect 2886 2503 2887 2504
rect 2862 2505 2863 2506
rect 2885 2505 2886 2506
rect 2615 2507 2616 2508
rect 2863 2507 2864 2508
rect 2616 2509 2617 2510
rect 2690 2509 2691 2510
rect 2915 2509 2916 2510
rect 2921 2509 2922 2510
rect 2948 2509 2949 2510
rect 2969 2509 2970 2510
rect 2035 2518 2036 2519
rect 2361 2518 2362 2519
rect 2038 2520 2039 2521
rect 2042 2520 2043 2521
rect 2049 2520 2050 2521
rect 2056 2520 2057 2521
rect 2063 2520 2064 2521
rect 2358 2520 2359 2521
rect 2080 2522 2081 2523
rect 2104 2522 2105 2523
rect 2084 2524 2085 2525
rect 2089 2524 2090 2525
rect 2093 2524 2094 2525
rect 2336 2524 2337 2525
rect 2095 2526 2096 2527
rect 2538 2526 2539 2527
rect 2098 2528 2099 2529
rect 2793 2528 2794 2529
rect 2100 2530 2101 2531
rect 2418 2530 2419 2531
rect 2110 2532 2111 2533
rect 2480 2532 2481 2533
rect 2077 2534 2078 2535
rect 2110 2534 2111 2535
rect 2114 2534 2115 2535
rect 2187 2534 2188 2535
rect 2129 2536 2130 2537
rect 2508 2536 2509 2537
rect 2133 2538 2134 2539
rect 2424 2538 2425 2539
rect 2139 2540 2140 2541
rect 2237 2540 2238 2541
rect 2142 2542 2143 2543
rect 2160 2542 2161 2543
rect 2145 2544 2146 2545
rect 2394 2544 2395 2545
rect 2147 2546 2148 2547
rect 2259 2546 2260 2547
rect 2148 2548 2149 2549
rect 2402 2548 2403 2549
rect 2176 2550 2177 2551
rect 2199 2550 2200 2551
rect 2188 2552 2189 2553
rect 2211 2552 2212 2553
rect 2206 2554 2207 2555
rect 2229 2554 2230 2555
rect 2224 2556 2225 2557
rect 2478 2556 2479 2557
rect 2227 2558 2228 2559
rect 2265 2558 2266 2559
rect 2231 2560 2232 2561
rect 2552 2560 2553 2561
rect 2243 2562 2244 2563
rect 2289 2562 2290 2563
rect 2247 2564 2248 2565
rect 2502 2564 2503 2565
rect 2255 2566 2256 2567
rect 2561 2566 2562 2567
rect 2261 2568 2262 2569
rect 2271 2568 2272 2569
rect 2267 2570 2268 2571
rect 2277 2570 2278 2571
rect 2291 2570 2292 2571
rect 2328 2570 2329 2571
rect 2297 2572 2298 2573
rect 2322 2572 2323 2573
rect 2304 2574 2305 2575
rect 2318 2574 2319 2575
rect 2303 2576 2304 2577
rect 2385 2576 2386 2577
rect 2310 2578 2311 2579
rect 2330 2578 2331 2579
rect 2316 2580 2317 2581
rect 2324 2580 2325 2581
rect 2295 2582 2296 2583
rect 2315 2582 2316 2583
rect 2340 2582 2341 2583
rect 2360 2582 2361 2583
rect 2342 2584 2343 2585
rect 2751 2584 2752 2585
rect 2352 2586 2353 2587
rect 2498 2586 2499 2587
rect 2355 2588 2356 2589
rect 2501 2588 2502 2589
rect 2334 2590 2335 2591
rect 2354 2590 2355 2591
rect 2313 2592 2314 2593
rect 2333 2592 2334 2593
rect 2366 2592 2367 2593
rect 2604 2592 2605 2593
rect 2373 2594 2374 2595
rect 2486 2594 2487 2595
rect 2364 2596 2365 2597
rect 2372 2596 2373 2597
rect 2376 2596 2377 2597
rect 2384 2596 2385 2597
rect 2375 2598 2376 2599
rect 2427 2598 2428 2599
rect 2066 2600 2067 2601
rect 2426 2600 2427 2601
rect 2391 2602 2392 2603
rect 2477 2602 2478 2603
rect 2390 2604 2391 2605
rect 2745 2604 2746 2605
rect 2406 2606 2407 2607
rect 2528 2606 2529 2607
rect 2408 2608 2409 2609
rect 2860 2608 2861 2609
rect 2412 2610 2413 2611
rect 2429 2610 2430 2611
rect 2397 2612 2398 2613
rect 2411 2612 2412 2613
rect 2370 2614 2371 2615
rect 2396 2614 2397 2615
rect 2415 2614 2416 2615
rect 2661 2614 2662 2615
rect 2400 2616 2401 2617
rect 2414 2616 2415 2617
rect 2436 2616 2437 2617
rect 2585 2616 2586 2617
rect 2435 2618 2436 2619
rect 2622 2618 2623 2619
rect 2442 2620 2443 2621
rect 2594 2620 2595 2621
rect 2166 2622 2167 2623
rect 2441 2622 2442 2623
rect 2167 2624 2168 2625
rect 2454 2624 2455 2625
rect 2448 2626 2449 2627
rect 2453 2626 2454 2627
rect 2163 2628 2164 2629
rect 2447 2628 2448 2629
rect 2164 2630 2165 2631
rect 2624 2630 2625 2631
rect 2460 2632 2461 2633
rect 2576 2632 2577 2633
rect 2466 2634 2467 2635
rect 2582 2634 2583 2635
rect 2097 2636 2098 2637
rect 2465 2636 2466 2637
rect 2472 2636 2473 2637
rect 2534 2636 2535 2637
rect 2475 2638 2476 2639
rect 2537 2638 2538 2639
rect 2474 2640 2475 2641
rect 2832 2640 2833 2641
rect 2490 2642 2491 2643
rect 2546 2642 2547 2643
rect 2489 2644 2490 2645
rect 2685 2644 2686 2645
rect 2496 2646 2497 2647
rect 2935 2646 2936 2647
rect 2382 2648 2383 2649
rect 2495 2648 2496 2649
rect 2510 2648 2511 2649
rect 2709 2648 2710 2649
rect 2516 2650 2517 2651
rect 2835 2650 2836 2651
rect 2520 2652 2521 2653
rect 2735 2652 2736 2653
rect 2522 2654 2523 2655
rect 2598 2654 2599 2655
rect 2445 2656 2446 2657
rect 2597 2656 2598 2657
rect 2544 2658 2545 2659
rect 2558 2658 2559 2659
rect 2568 2658 2569 2659
rect 2720 2658 2721 2659
rect 2567 2660 2568 2661
rect 2784 2660 2785 2661
rect 2570 2662 2571 2663
rect 2703 2662 2704 2663
rect 2550 2664 2551 2665
rect 2702 2664 2703 2665
rect 2574 2666 2575 2667
rect 2726 2666 2727 2667
rect 2592 2668 2593 2669
rect 2877 2668 2878 2669
rect 2607 2670 2608 2671
rect 2805 2670 2806 2671
rect 2532 2672 2533 2673
rect 2606 2672 2607 2673
rect 2421 2674 2422 2675
rect 2531 2674 2532 2675
rect 2420 2676 2421 2677
rect 2715 2676 2716 2677
rect 2580 2678 2581 2679
rect 2714 2678 2715 2679
rect 2612 2680 2613 2681
rect 2655 2680 2656 2681
rect 2616 2682 2617 2683
rect 2711 2682 2712 2683
rect 2619 2684 2620 2685
rect 2690 2684 2691 2685
rect 2618 2686 2619 2687
rect 2856 2686 2857 2687
rect 2628 2688 2629 2689
rect 2750 2688 2751 2689
rect 2346 2690 2347 2691
rect 2627 2690 2628 2691
rect 2639 2690 2640 2691
rect 2748 2690 2749 2691
rect 2654 2692 2655 2693
rect 2891 2692 2892 2693
rect 2657 2694 2658 2695
rect 2760 2694 2761 2695
rect 2621 2696 2622 2697
rect 2759 2696 2760 2697
rect 2667 2698 2668 2699
rect 2906 2698 2907 2699
rect 2673 2700 2674 2701
rect 2945 2700 2946 2701
rect 2526 2702 2527 2703
rect 2672 2702 2673 2703
rect 2525 2704 2526 2705
rect 2829 2704 2830 2705
rect 2679 2706 2680 2707
rect 2938 2706 2939 2707
rect 2469 2708 2470 2709
rect 2678 2708 2679 2709
rect 2280 2710 2281 2711
rect 2468 2710 2469 2711
rect 2129 2712 2130 2713
rect 2279 2712 2280 2713
rect 2684 2712 2685 2713
rect 2733 2712 2734 2713
rect 2697 2714 2698 2715
rect 2982 2714 2983 2715
rect 2556 2716 2557 2717
rect 2696 2716 2697 2717
rect 2700 2716 2701 2717
rect 2979 2716 2980 2717
rect 2708 2718 2709 2719
rect 2891 2718 2892 2719
rect 2732 2720 2733 2721
rect 2847 2720 2848 2721
rect 2738 2722 2739 2723
rect 2972 2722 2973 2723
rect 2744 2724 2745 2725
rect 2912 2724 2913 2725
rect 2757 2726 2758 2727
rect 2863 2726 2864 2727
rect 2763 2728 2764 2729
rect 2894 2728 2895 2729
rect 2631 2730 2632 2731
rect 2894 2730 2895 2731
rect 2630 2732 2631 2733
rect 2649 2732 2650 2733
rect 2648 2734 2649 2735
rect 2900 2734 2901 2735
rect 2637 2736 2638 2737
rect 2901 2736 2902 2737
rect 2484 2738 2485 2739
rect 2636 2738 2637 2739
rect 2126 2740 2127 2741
rect 2483 2740 2484 2741
rect 2125 2742 2126 2743
rect 2193 2742 2194 2743
rect 2194 2744 2195 2745
rect 2217 2744 2218 2745
rect 2218 2746 2219 2747
rect 2241 2746 2242 2747
rect 2772 2746 2773 2747
rect 2777 2746 2778 2747
rect 2783 2746 2784 2747
rect 2796 2746 2797 2747
rect 2787 2748 2788 2749
rect 2853 2748 2854 2749
rect 2786 2750 2787 2751
rect 2966 2750 2967 2751
rect 2792 2752 2793 2753
rect 2844 2752 2845 2753
rect 2122 2754 2123 2755
rect 2844 2754 2845 2755
rect 2795 2756 2796 2757
rect 2811 2756 2812 2757
rect 2154 2758 2155 2759
rect 2810 2758 2811 2759
rect 2798 2760 2799 2761
rect 2814 2760 2815 2761
rect 2790 2762 2791 2763
rect 2814 2762 2815 2763
rect 2789 2764 2790 2765
rect 2841 2764 2842 2765
rect 2801 2766 2802 2767
rect 2823 2766 2824 2767
rect 2808 2768 2809 2769
rect 2838 2768 2839 2769
rect 2807 2770 2808 2771
rect 2850 2770 2851 2771
rect 2817 2772 2818 2773
rect 2963 2772 2964 2773
rect 2820 2774 2821 2775
rect 2885 2774 2886 2775
rect 2823 2776 2824 2777
rect 2888 2776 2889 2777
rect 2826 2778 2827 2779
rect 2908 2778 2909 2779
rect 2829 2780 2830 2781
rect 2873 2780 2874 2781
rect 2841 2782 2842 2783
rect 2897 2782 2898 2783
rect 2859 2784 2860 2785
rect 2942 2784 2943 2785
rect 2862 2786 2863 2787
rect 2928 2786 2929 2787
rect 2871 2788 2872 2789
rect 2915 2788 2916 2789
rect 2775 2790 2776 2791
rect 2915 2790 2916 2791
rect 2874 2792 2875 2793
rect 2918 2792 2919 2793
rect 2879 2794 2880 2795
rect 2949 2794 2950 2795
rect 2918 2796 2919 2797
rect 2969 2796 2970 2797
rect 2935 2798 2936 2799
rect 2942 2798 2943 2799
rect 2059 2807 2060 2808
rect 2154 2807 2155 2808
rect 2065 2809 2066 2810
rect 2480 2809 2481 2810
rect 2068 2811 2069 2812
rect 2084 2811 2085 2812
rect 2069 2813 2070 2814
rect 2110 2813 2111 2814
rect 2075 2815 2076 2816
rect 2261 2815 2262 2816
rect 2076 2817 2077 2818
rect 2495 2817 2496 2818
rect 2083 2819 2084 2820
rect 2465 2819 2466 2820
rect 2087 2821 2088 2822
rect 2426 2821 2427 2822
rect 2093 2823 2094 2824
rect 2627 2823 2628 2824
rect 2094 2825 2095 2826
rect 2188 2825 2189 2826
rect 2097 2827 2098 2828
rect 2477 2827 2478 2828
rect 2104 2829 2105 2830
rect 2525 2829 2526 2830
rect 2119 2831 2120 2832
rect 2372 2831 2373 2832
rect 2122 2833 2123 2834
rect 2333 2833 2334 2834
rect 2125 2835 2126 2836
rect 2396 2835 2397 2836
rect 2080 2837 2081 2838
rect 2125 2837 2126 2838
rect 2129 2837 2130 2838
rect 2468 2837 2469 2838
rect 2112 2839 2113 2840
rect 2469 2839 2470 2840
rect 2131 2841 2132 2842
rect 2447 2841 2448 2842
rect 2136 2843 2137 2844
rect 2384 2843 2385 2844
rect 2135 2845 2136 2846
rect 2214 2845 2215 2846
rect 2142 2847 2143 2848
rect 2157 2847 2158 2848
rect 2142 2849 2143 2850
rect 2534 2849 2535 2850
rect 2145 2851 2146 2852
rect 2334 2851 2335 2852
rect 2145 2853 2146 2854
rect 2582 2853 2583 2854
rect 2160 2855 2161 2856
rect 2486 2855 2487 2856
rect 2163 2857 2164 2858
rect 2194 2857 2195 2858
rect 2167 2859 2168 2860
rect 2594 2859 2595 2860
rect 2176 2861 2177 2862
rect 2190 2861 2191 2862
rect 2178 2863 2179 2864
rect 2218 2863 2219 2864
rect 2196 2865 2197 2866
rect 2366 2865 2367 2866
rect 2199 2867 2200 2868
rect 2624 2867 2625 2868
rect 2202 2869 2203 2870
rect 2243 2869 2244 2870
rect 2206 2871 2207 2872
rect 2289 2871 2290 2872
rect 2208 2873 2209 2874
rect 2237 2873 2238 2874
rect 2220 2875 2221 2876
rect 2406 2875 2407 2876
rect 2224 2877 2225 2878
rect 2706 2877 2707 2878
rect 2223 2879 2224 2880
rect 2639 2879 2640 2880
rect 2227 2881 2228 2882
rect 2328 2881 2329 2882
rect 2231 2883 2232 2884
rect 2435 2883 2436 2884
rect 2152 2885 2153 2886
rect 2436 2885 2437 2886
rect 2232 2887 2233 2888
rect 2267 2887 2268 2888
rect 2244 2889 2245 2890
rect 2279 2889 2280 2890
rect 2262 2891 2263 2892
rect 2291 2891 2292 2892
rect 2268 2893 2269 2894
rect 2315 2893 2316 2894
rect 2271 2895 2272 2896
rect 2318 2895 2319 2896
rect 2277 2897 2278 2898
rect 2324 2897 2325 2898
rect 2283 2899 2284 2900
rect 2330 2899 2331 2900
rect 2286 2901 2287 2902
rect 2336 2901 2337 2902
rect 2297 2903 2298 2904
rect 2394 2903 2395 2904
rect 2303 2905 2304 2906
rect 2331 2905 2332 2906
rect 2304 2907 2305 2908
rect 2354 2907 2355 2908
rect 2310 2909 2311 2910
rect 2360 2909 2361 2910
rect 2313 2911 2314 2912
rect 2375 2911 2376 2912
rect 2072 2913 2073 2914
rect 2376 2913 2377 2914
rect 2322 2915 2323 2916
rect 2342 2915 2343 2916
rect 2340 2917 2341 2918
rect 2498 2917 2499 2918
rect 2343 2919 2344 2920
rect 2501 2919 2502 2920
rect 2346 2921 2347 2922
rect 2402 2921 2403 2922
rect 2352 2923 2353 2924
rect 2414 2923 2415 2924
rect 2355 2925 2356 2926
rect 2597 2925 2598 2926
rect 2358 2927 2359 2928
rect 2408 2927 2409 2928
rect 2364 2929 2365 2930
rect 2420 2929 2421 2930
rect 2370 2931 2371 2932
rect 2429 2931 2430 2932
rect 2379 2933 2380 2934
rect 2453 2933 2454 2934
rect 2382 2935 2383 2936
rect 2537 2935 2538 2936
rect 2385 2937 2386 2938
rect 2390 2937 2391 2938
rect 2391 2939 2392 2940
rect 2483 2939 2484 2940
rect 2397 2941 2398 2942
rect 2528 2941 2529 2942
rect 2400 2943 2401 2944
rect 2531 2943 2532 2944
rect 2403 2945 2404 2946
rect 2762 2945 2763 2946
rect 2411 2947 2412 2948
rect 2439 2947 2440 2948
rect 2424 2949 2425 2950
rect 2489 2949 2490 2950
rect 2430 2951 2431 2952
rect 2516 2951 2517 2952
rect 2441 2953 2442 2954
rect 2484 2953 2485 2954
rect 2442 2955 2443 2956
rect 2576 2955 2577 2956
rect 2445 2957 2446 2958
rect 2585 2957 2586 2958
rect 2448 2959 2449 2960
rect 2522 2959 2523 2960
rect 2454 2961 2455 2962
rect 2552 2961 2553 2962
rect 2460 2963 2461 2964
rect 2546 2963 2547 2964
rect 2466 2965 2467 2966
rect 2636 2965 2637 2966
rect 2472 2967 2473 2968
rect 2558 2967 2559 2968
rect 2474 2969 2475 2970
rect 2481 2969 2482 2970
rect 2475 2971 2476 2972
rect 2561 2971 2562 2972
rect 2478 2973 2479 2974
rect 2510 2973 2511 2974
rect 2490 2975 2491 2976
rect 2735 2975 2736 2976
rect 2496 2977 2497 2978
rect 2810 2977 2811 2978
rect 2508 2979 2509 2980
rect 2630 2979 2631 2980
rect 2514 2981 2515 2982
rect 2730 2981 2731 2982
rect 2526 2983 2527 2984
rect 2877 2983 2878 2984
rect 2532 2985 2533 2986
rect 2696 2985 2697 2986
rect 2544 2987 2545 2988
rect 2702 2987 2703 2988
rect 2550 2989 2551 2990
rect 2894 2989 2895 2990
rect 2553 2991 2554 2992
rect 2708 2991 2709 2992
rect 2556 2993 2557 2994
rect 2612 2993 2613 2994
rect 2562 2995 2563 2996
rect 2720 2995 2721 2996
rect 2567 2997 2568 2998
rect 2688 2997 2689 2998
rect 2241 2999 2242 3000
rect 2568 2999 2569 3000
rect 2570 2999 2571 3000
rect 2759 2999 2760 3000
rect 2574 3001 2575 3002
rect 2838 3001 2839 3002
rect 2580 3003 2581 3004
rect 2648 3003 2649 3004
rect 2592 3005 2593 3006
rect 2853 3005 2854 3006
rect 2595 3007 2596 3008
rect 2846 3007 2847 3008
rect 2598 3009 2599 3010
rect 2901 3009 2902 3010
rect 2604 3011 2605 3012
rect 2744 3011 2745 3012
rect 2606 3013 2607 3014
rect 2718 3013 2719 3014
rect 2610 3015 2611 3016
rect 2750 3015 2751 3016
rect 2613 3017 2614 3018
rect 2823 3017 2824 3018
rect 2618 3019 2619 3020
rect 2817 3019 2818 3020
rect 2631 3021 2632 3022
rect 2654 3021 2655 3022
rect 2634 3023 2635 3024
rect 2657 3023 2658 3024
rect 2637 3025 2638 3026
rect 2850 3025 2851 3026
rect 2643 3027 2644 3028
rect 2697 3027 2698 3028
rect 2672 3029 2673 3030
rect 2835 3029 2836 3030
rect 2673 3031 2674 3032
rect 2798 3031 2799 3032
rect 2676 3033 2677 3034
rect 2684 3033 2685 3034
rect 2621 3035 2622 3036
rect 2685 3035 2686 3036
rect 2678 3037 2679 3038
rect 2757 3037 2758 3038
rect 2679 3039 2680 3040
rect 2783 3039 2784 3040
rect 2682 3041 2683 3042
rect 2786 3041 2787 3042
rect 2502 3043 2503 3044
rect 2785 3043 2786 3044
rect 2690 3045 2691 3046
rect 2891 3045 2892 3046
rect 2691 3047 2692 3048
rect 2844 3047 2845 3048
rect 2703 3049 2704 3050
rect 2732 3049 2733 3050
rect 2709 3051 2710 3052
rect 2789 3051 2790 3052
rect 2711 3053 2712 3054
rect 2788 3053 2789 3054
rect 2712 3055 2713 3056
rect 2792 3055 2793 3056
rect 2733 3057 2734 3058
rect 2820 3057 2821 3058
rect 2736 3059 2737 3060
rect 2748 3059 2749 3060
rect 2738 3061 2739 3062
rect 2912 3061 2913 3062
rect 2739 3063 2740 3064
rect 2826 3063 2827 3064
rect 2754 3065 2755 3066
rect 2841 3065 2842 3066
rect 2760 3067 2761 3068
rect 2862 3067 2863 3068
rect 2763 3069 2764 3070
rect 2777 3069 2778 3070
rect 2772 3071 2773 3072
rect 2871 3071 2872 3072
rect 2775 3073 2776 3074
rect 2874 3073 2875 3074
rect 2781 3075 2782 3076
rect 2795 3075 2796 3076
rect 2801 3075 2802 3076
rect 2884 3075 2885 3076
rect 2826 3077 2827 3078
rect 2918 3077 2919 3078
rect 2829 3079 2830 3080
rect 2938 3079 2939 3080
rect 2726 3081 2727 3082
rect 2829 3081 2830 3082
rect 2714 3083 2715 3084
rect 2727 3083 2728 3084
rect 2859 3083 2860 3084
rect 2931 3083 2932 3084
rect 2062 3092 2063 3093
rect 2190 3092 2191 3093
rect 2065 3094 2066 3095
rect 2374 3094 2375 3095
rect 2087 3096 2088 3097
rect 2277 3096 2278 3097
rect 2097 3098 2098 3099
rect 2289 3098 2290 3099
rect 2079 3100 2080 3101
rect 2098 3100 2099 3101
rect 2101 3100 2102 3101
rect 2304 3100 2305 3101
rect 2104 3102 2105 3103
rect 2125 3102 2126 3103
rect 2110 3104 2111 3105
rect 2400 3104 2401 3105
rect 2115 3106 2116 3107
rect 2394 3106 2395 3107
rect 2073 3108 2074 3109
rect 2395 3108 2396 3109
rect 2114 3110 2115 3111
rect 2313 3110 2314 3111
rect 2120 3112 2121 3113
rect 2154 3112 2155 3113
rect 2123 3114 2124 3115
rect 2157 3114 2158 3115
rect 2126 3116 2127 3117
rect 2346 3116 2347 3117
rect 2135 3118 2136 3119
rect 2176 3118 2177 3119
rect 2138 3120 2139 3121
rect 2208 3120 2209 3121
rect 2142 3122 2143 3123
rect 2262 3122 2263 3123
rect 2141 3124 2142 3125
rect 2305 3124 2306 3125
rect 2145 3126 2146 3127
rect 2442 3126 2443 3127
rect 2157 3128 2158 3129
rect 2178 3128 2179 3129
rect 2173 3130 2174 3131
rect 2281 3130 2282 3131
rect 2182 3132 2183 3133
rect 2214 3132 2215 3133
rect 2202 3134 2203 3135
rect 2368 3134 2369 3135
rect 2218 3136 2219 3137
rect 2244 3136 2245 3137
rect 2224 3138 2225 3139
rect 2355 3138 2356 3139
rect 2232 3140 2233 3141
rect 2362 3140 2363 3141
rect 2236 3142 2237 3143
rect 2385 3142 2386 3143
rect 2238 3144 2239 3145
rect 2382 3144 2383 3145
rect 2241 3146 2242 3147
rect 2472 3146 2473 3147
rect 2242 3148 2243 3149
rect 2268 3148 2269 3149
rect 2263 3150 2264 3151
rect 2286 3150 2287 3151
rect 2269 3152 2270 3153
rect 2310 3152 2311 3153
rect 2138 3154 2139 3155
rect 2311 3154 2312 3155
rect 2283 3156 2284 3157
rect 2410 3156 2411 3157
rect 2293 3158 2294 3159
rect 2328 3158 2329 3159
rect 2296 3160 2297 3161
rect 2331 3160 2332 3161
rect 2317 3162 2318 3163
rect 2358 3162 2359 3163
rect 2083 3164 2084 3165
rect 2359 3164 2360 3165
rect 2329 3166 2330 3167
rect 2334 3166 2335 3167
rect 2335 3168 2336 3169
rect 2340 3168 2341 3169
rect 2338 3170 2339 3171
rect 2343 3170 2344 3171
rect 2341 3172 2342 3173
rect 2370 3172 2371 3173
rect 2347 3174 2348 3175
rect 2364 3174 2365 3175
rect 2365 3176 2366 3177
rect 2379 3176 2380 3177
rect 2371 3178 2372 3179
rect 2376 3178 2377 3179
rect 2383 3178 2384 3179
rect 2406 3178 2407 3179
rect 2072 3180 2073 3181
rect 2407 3180 2408 3181
rect 2389 3182 2390 3183
rect 2391 3182 2392 3183
rect 2112 3184 2113 3185
rect 2392 3184 2393 3185
rect 2397 3184 2398 3185
rect 2401 3184 2402 3185
rect 2076 3186 2077 3187
rect 2398 3186 2399 3187
rect 2075 3188 2076 3189
rect 2271 3188 2272 3189
rect 2403 3188 2404 3189
rect 2413 3188 2414 3189
rect 2094 3190 2095 3191
rect 2404 3190 2405 3191
rect 2094 3192 2095 3193
rect 2272 3192 2273 3193
rect 2422 3192 2423 3193
rect 2478 3192 2479 3193
rect 2428 3194 2429 3195
rect 2445 3194 2446 3195
rect 2436 3196 2437 3197
rect 2443 3196 2444 3197
rect 2424 3198 2425 3199
rect 2437 3198 2438 3199
rect 2439 3198 2440 3199
rect 2446 3198 2447 3199
rect 2448 3198 2449 3199
rect 2650 3198 2651 3199
rect 2160 3200 2161 3201
rect 2449 3200 2450 3201
rect 2466 3200 2467 3201
rect 2473 3200 2474 3201
rect 2460 3202 2461 3203
rect 2467 3202 2468 3203
rect 2454 3204 2455 3205
rect 2461 3204 2462 3205
rect 2430 3206 2431 3207
rect 2455 3206 2456 3207
rect 2131 3208 2132 3209
rect 2431 3208 2432 3209
rect 2479 3208 2480 3209
rect 2653 3208 2654 3209
rect 2490 3210 2491 3211
rect 2718 3210 2719 3211
rect 2287 3212 2288 3213
rect 2491 3212 2492 3213
rect 2496 3212 2497 3213
rect 2730 3212 2731 3213
rect 2484 3214 2485 3215
rect 2497 3214 2498 3215
rect 2502 3214 2503 3215
rect 2696 3214 2697 3215
rect 2503 3216 2504 3217
rect 2508 3216 2509 3217
rect 2521 3216 2522 3217
rect 2712 3216 2713 3217
rect 2524 3218 2525 3219
rect 2568 3218 2569 3219
rect 2532 3220 2533 3221
rect 2539 3220 2540 3221
rect 2536 3222 2537 3223
rect 2550 3222 2551 3223
rect 2542 3224 2543 3225
rect 2544 3224 2545 3225
rect 2553 3224 2554 3225
rect 2820 3224 2821 3225
rect 2554 3226 2555 3227
rect 2580 3226 2581 3227
rect 2556 3228 2557 3229
rect 2711 3228 2712 3229
rect 2560 3230 2561 3231
rect 2562 3230 2563 3231
rect 2572 3230 2573 3231
rect 2631 3230 2632 3231
rect 2574 3232 2575 3233
rect 2660 3232 2661 3233
rect 2575 3234 2576 3235
rect 2634 3234 2635 3235
rect 2578 3236 2579 3237
rect 2669 3236 2670 3237
rect 2590 3238 2591 3239
rect 2800 3238 2801 3239
rect 2592 3240 2593 3241
rect 2846 3240 2847 3241
rect 2593 3242 2594 3243
rect 2610 3242 2611 3243
rect 2595 3244 2596 3245
rect 2839 3244 2840 3245
rect 2475 3246 2476 3247
rect 2596 3246 2597 3247
rect 2469 3248 2470 3249
rect 2476 3248 2477 3249
rect 2598 3248 2599 3249
rect 2836 3248 2837 3249
rect 2322 3250 2323 3251
rect 2599 3250 2600 3251
rect 2323 3252 2324 3253
rect 2352 3252 2353 3253
rect 2128 3254 2129 3255
rect 2353 3254 2354 3255
rect 2129 3256 2130 3257
rect 2434 3256 2435 3257
rect 2602 3256 2603 3257
rect 2832 3256 2833 3257
rect 2604 3258 2605 3259
rect 2803 3258 2804 3259
rect 2613 3260 2614 3261
rect 2720 3260 2721 3261
rect 2620 3262 2621 3263
rect 2685 3262 2686 3263
rect 2623 3264 2624 3265
rect 2643 3264 2644 3265
rect 2632 3266 2633 3267
rect 2806 3266 2807 3267
rect 2635 3268 2636 3269
rect 2823 3268 2824 3269
rect 2641 3270 2642 3271
rect 2682 3270 2683 3271
rect 2644 3272 2645 3273
rect 2741 3272 2742 3273
rect 2663 3274 2664 3275
rect 2703 3274 2704 3275
rect 2666 3276 2667 3277
rect 2706 3276 2707 3277
rect 2673 3278 2674 3279
rect 2777 3278 2778 3279
rect 2676 3280 2677 3281
rect 2809 3280 2810 3281
rect 2675 3282 2676 3283
rect 2787 3282 2788 3283
rect 2681 3284 2682 3285
rect 2817 3284 2818 3285
rect 2684 3286 2685 3287
rect 2813 3286 2814 3287
rect 2688 3288 2689 3289
rect 2700 3288 2701 3289
rect 2702 3288 2703 3289
rect 2791 3288 2792 3289
rect 2709 3290 2710 3291
rect 2784 3290 2785 3291
rect 2708 3292 2709 3293
rect 2733 3292 2734 3293
rect 2723 3294 2724 3295
rect 2748 3294 2749 3295
rect 2726 3296 2727 3297
rect 2754 3296 2755 3297
rect 2729 3298 2730 3299
rect 2757 3298 2758 3299
rect 2732 3300 2733 3301
rect 2760 3300 2761 3301
rect 2514 3302 2515 3303
rect 2759 3302 2760 3303
rect 2515 3304 2516 3305
rect 2637 3304 2638 3305
rect 2638 3306 2639 3307
rect 2679 3306 2680 3307
rect 2736 3306 2737 3307
rect 2751 3306 2752 3307
rect 2735 3308 2736 3309
rect 2763 3308 2764 3309
rect 2739 3310 2740 3311
rect 2766 3310 2767 3311
rect 2691 3312 2692 3313
rect 2738 3312 2739 3313
rect 2690 3314 2691 3315
rect 2780 3314 2781 3315
rect 2750 3316 2751 3317
rect 2772 3316 2773 3317
rect 2526 3318 2527 3319
rect 2773 3318 2774 3319
rect 2753 3320 2754 3321
rect 2775 3320 2776 3321
rect 2797 3320 2798 3321
rect 2826 3320 2827 3321
rect 2011 3329 2012 3330
rect 2338 3329 2339 3330
rect 2065 3331 2066 3332
rect 2395 3331 2396 3332
rect 2068 3333 2069 3334
rect 2267 3333 2268 3334
rect 2068 3335 2069 3336
rect 2398 3335 2399 3336
rect 2072 3337 2073 3338
rect 2138 3337 2139 3338
rect 2079 3339 2080 3340
rect 2389 3339 2390 3340
rect 2082 3341 2083 3342
rect 2387 3341 2388 3342
rect 2094 3343 2095 3344
rect 2263 3343 2264 3344
rect 2098 3345 2099 3346
rect 2252 3345 2253 3346
rect 2108 3347 2109 3348
rect 2120 3347 2121 3348
rect 2114 3349 2115 3350
rect 2261 3349 2262 3350
rect 2041 3351 2042 3352
rect 2114 3351 2115 3352
rect 2117 3351 2118 3352
rect 2272 3351 2273 3352
rect 2117 3353 2118 3354
rect 2123 3353 2124 3354
rect 2120 3355 2121 3356
rect 2309 3355 2310 3356
rect 2126 3357 2127 3358
rect 2323 3357 2324 3358
rect 2127 3359 2128 3360
rect 2218 3359 2219 3360
rect 2129 3361 2130 3362
rect 2148 3361 2149 3362
rect 2141 3363 2142 3364
rect 2285 3363 2286 3364
rect 2166 3365 2167 3366
rect 2392 3365 2393 3366
rect 2153 3367 2154 3368
rect 2393 3367 2394 3368
rect 2157 3369 2158 3370
rect 2165 3369 2166 3370
rect 2156 3371 2157 3372
rect 2585 3371 2586 3372
rect 2171 3373 2172 3374
rect 2368 3373 2369 3374
rect 2173 3375 2174 3376
rect 2296 3375 2297 3376
rect 2174 3377 2175 3378
rect 2663 3377 2664 3378
rect 2176 3379 2177 3380
rect 2287 3379 2288 3380
rect 2177 3381 2178 3382
rect 2182 3381 2183 3382
rect 2207 3381 2208 3382
rect 2449 3381 2450 3382
rect 2224 3383 2225 3384
rect 2234 3383 2235 3384
rect 2225 3385 2226 3386
rect 2242 3385 2243 3386
rect 2228 3387 2229 3388
rect 2410 3387 2411 3388
rect 2210 3389 2211 3390
rect 2411 3389 2412 3390
rect 2239 3391 2240 3392
rect 2357 3391 2358 3392
rect 2243 3393 2244 3394
rect 2365 3393 2366 3394
rect 2258 3395 2259 3396
rect 2269 3395 2270 3396
rect 2104 3397 2105 3398
rect 2270 3397 2271 3398
rect 2279 3397 2280 3398
rect 2293 3397 2294 3398
rect 2291 3399 2292 3400
rect 2305 3399 2306 3400
rect 2297 3401 2298 3402
rect 2311 3401 2312 3402
rect 2303 3403 2304 3404
rect 2317 3403 2318 3404
rect 2312 3405 2313 3406
rect 2329 3405 2330 3406
rect 2324 3407 2325 3408
rect 2341 3407 2342 3408
rect 2330 3409 2331 3410
rect 2347 3409 2348 3410
rect 2339 3411 2340 3412
rect 2353 3411 2354 3412
rect 2345 3413 2346 3414
rect 2359 3413 2360 3414
rect 2351 3415 2352 3416
rect 2383 3415 2384 3416
rect 2362 3417 2363 3418
rect 2390 3417 2391 3418
rect 2363 3419 2364 3420
rect 2437 3419 2438 3420
rect 2369 3421 2370 3422
rect 2371 3421 2372 3422
rect 2372 3423 2373 3424
rect 2374 3423 2375 3424
rect 2375 3425 2376 3426
rect 2401 3425 2402 3426
rect 2087 3427 2088 3428
rect 2402 3427 2403 3428
rect 2378 3429 2379 3430
rect 2404 3429 2405 3430
rect 2396 3431 2397 3432
rect 2428 3431 2429 3432
rect 2399 3433 2400 3434
rect 2413 3433 2414 3434
rect 2405 3435 2406 3436
rect 2407 3435 2408 3436
rect 2075 3437 2076 3438
rect 2408 3437 2409 3438
rect 2429 3437 2430 3438
rect 2431 3437 2432 3438
rect 2432 3439 2433 3440
rect 2434 3439 2435 3440
rect 2435 3441 2436 3442
rect 2461 3441 2462 3442
rect 2441 3443 2442 3444
rect 2491 3443 2492 3444
rect 2446 3445 2447 3446
rect 2450 3445 2451 3446
rect 2443 3447 2444 3448
rect 2447 3447 2448 3448
rect 2453 3447 2454 3448
rect 2467 3447 2468 3448
rect 2455 3449 2456 3450
rect 2650 3449 2651 3450
rect 2465 3451 2466 3452
rect 2669 3451 2670 3452
rect 2471 3453 2472 3454
rect 2473 3453 2474 3454
rect 2474 3455 2475 3456
rect 2476 3455 2477 3456
rect 2240 3457 2241 3458
rect 2477 3457 2478 3458
rect 2482 3457 2483 3458
rect 2501 3457 2502 3458
rect 2483 3459 2484 3460
rect 2696 3459 2697 3460
rect 2489 3461 2490 3462
rect 2596 3461 2597 3462
rect 2492 3463 2493 3464
rect 2599 3463 2600 3464
rect 2495 3465 2496 3466
rect 2711 3465 2712 3466
rect 2497 3467 2498 3468
rect 2612 3467 2613 3468
rect 2507 3469 2508 3470
rect 2723 3469 2724 3470
rect 2515 3471 2516 3472
rect 2660 3471 2661 3472
rect 2521 3473 2522 3474
rect 2528 3473 2529 3474
rect 2542 3473 2543 3474
rect 2549 3473 2550 3474
rect 2543 3475 2544 3476
rect 2572 3475 2573 3476
rect 2546 3477 2547 3478
rect 2575 3477 2576 3478
rect 2554 3479 2555 3480
rect 2737 3479 2738 3480
rect 2539 3481 2540 3482
rect 2555 3481 2556 3482
rect 2560 3481 2561 3482
rect 2567 3481 2568 3482
rect 2578 3481 2579 3482
rect 2657 3481 2658 3482
rect 2593 3483 2594 3484
rect 2606 3483 2607 3484
rect 2609 3483 2610 3484
rect 2666 3483 2667 3484
rect 2503 3485 2504 3486
rect 2667 3485 2668 3486
rect 2422 3487 2423 3488
rect 2504 3487 2505 3488
rect 2423 3489 2424 3490
rect 2479 3489 2480 3490
rect 2620 3489 2621 3490
rect 2657 3489 2658 3490
rect 2623 3491 2624 3492
rect 2648 3491 2649 3492
rect 2627 3493 2628 3494
rect 2780 3493 2781 3494
rect 2519 3495 2520 3496
rect 2780 3495 2781 3496
rect 2630 3497 2631 3498
rect 2635 3497 2636 3498
rect 2632 3499 2633 3500
rect 2777 3499 2778 3500
rect 2633 3501 2634 3502
rect 2638 3501 2639 3502
rect 2636 3503 2637 3504
rect 2641 3503 2642 3504
rect 2639 3505 2640 3506
rect 2740 3505 2741 3506
rect 2644 3507 2645 3508
rect 2832 3507 2833 3508
rect 2645 3509 2646 3510
rect 2660 3509 2661 3510
rect 2675 3509 2676 3510
rect 2695 3509 2696 3510
rect 2702 3509 2703 3510
rect 2713 3509 2714 3510
rect 2701 3511 2702 3512
rect 2811 3511 2812 3512
rect 2720 3513 2721 3514
rect 2804 3513 2805 3514
rect 2726 3515 2727 3516
rect 2743 3515 2744 3516
rect 2725 3517 2726 3518
rect 2759 3517 2760 3518
rect 2729 3519 2730 3520
rect 2746 3519 2747 3520
rect 2708 3521 2709 3522
rect 2728 3521 2729 3522
rect 2690 3523 2691 3524
rect 2707 3523 2708 3524
rect 2750 3523 2751 3524
rect 2761 3523 2762 3524
rect 2732 3525 2733 3526
rect 2749 3525 2750 3526
rect 2753 3525 2754 3526
rect 2764 3525 2765 3526
rect 2735 3527 2736 3528
rect 2752 3527 2753 3528
rect 2734 3529 2735 3530
rect 2787 3529 2788 3530
rect 2767 3531 2768 3532
rect 2807 3531 2808 3532
rect 2684 3533 2685 3534
rect 2808 3533 2809 3534
rect 2773 3535 2774 3536
rect 2784 3535 2785 3536
rect 2264 3537 2265 3538
rect 2773 3537 2774 3538
rect 2674 3539 2675 3540
rect 2783 3539 2784 3540
rect 2797 3539 2798 3540
rect 2838 3539 2839 3540
rect 2677 3541 2678 3542
rect 2797 3541 2798 3542
rect 2817 3541 2818 3542
rect 2825 3541 2826 3542
rect 2814 3543 2815 3544
rect 2818 3543 2819 3544
rect 2731 3545 2732 3546
rect 2815 3545 2816 3546
rect 2038 3554 2039 3555
rect 2225 3554 2226 3555
rect 2044 3556 2045 3557
rect 2108 3556 2109 3557
rect 2052 3558 2053 3559
rect 2059 3558 2060 3559
rect 2056 3560 2057 3561
rect 2345 3560 2346 3561
rect 2066 3562 2067 3563
rect 2270 3562 2271 3563
rect 2072 3564 2073 3565
rect 2429 3564 2430 3565
rect 2068 3566 2069 3567
rect 2073 3566 2074 3567
rect 2084 3566 2085 3567
rect 2390 3566 2391 3567
rect 2084 3568 2085 3569
rect 2199 3568 2200 3569
rect 2094 3570 2095 3571
rect 2402 3570 2403 3571
rect 2102 3572 2103 3573
rect 2378 3572 2379 3573
rect 2105 3574 2106 3575
rect 2220 3574 2221 3575
rect 2106 3576 2107 3577
rect 2375 3576 2376 3577
rect 2110 3578 2111 3579
rect 2252 3578 2253 3579
rect 2114 3580 2115 3581
rect 2123 3580 2124 3581
rect 2117 3582 2118 3583
rect 2126 3582 2127 3583
rect 2117 3584 2118 3585
rect 2277 3584 2278 3585
rect 2130 3586 2131 3587
rect 2289 3586 2290 3587
rect 2129 3588 2130 3589
rect 2655 3588 2656 3589
rect 2132 3590 2133 3591
rect 2234 3590 2235 3591
rect 2134 3592 2135 3593
rect 2253 3592 2254 3593
rect 2137 3594 2138 3595
rect 2483 3594 2484 3595
rect 2139 3596 2140 3597
rect 2291 3596 2292 3597
rect 2146 3598 2147 3599
rect 2376 3598 2377 3599
rect 2184 3600 2185 3601
rect 2282 3600 2283 3601
rect 2087 3602 2088 3603
rect 2283 3602 2284 3603
rect 2190 3604 2191 3605
rect 2228 3604 2229 3605
rect 2192 3606 2193 3607
rect 2435 3606 2436 3607
rect 2196 3608 2197 3609
rect 2267 3608 2268 3609
rect 2205 3610 2206 3611
rect 2336 3610 2337 3611
rect 2207 3612 2208 3613
rect 2367 3612 2368 3613
rect 2165 3614 2166 3615
rect 2208 3614 2209 3615
rect 2217 3614 2218 3615
rect 2355 3614 2356 3615
rect 2223 3616 2224 3617
rect 2258 3616 2259 3617
rect 2229 3618 2230 3619
rect 2339 3618 2340 3619
rect 2235 3620 2236 3621
rect 2369 3620 2370 3621
rect 2238 3622 2239 3623
rect 2372 3622 2373 3623
rect 2177 3624 2178 3625
rect 2373 3624 2374 3625
rect 2178 3626 2179 3627
rect 2450 3626 2451 3627
rect 2241 3628 2242 3629
rect 2432 3628 2433 3629
rect 2243 3630 2244 3631
rect 2453 3630 2454 3631
rect 2250 3632 2251 3633
rect 2387 3632 2388 3633
rect 2256 3634 2257 3635
rect 2309 3634 2310 3635
rect 2261 3636 2262 3637
rect 2292 3636 2293 3637
rect 2262 3638 2263 3639
rect 2405 3638 2406 3639
rect 2268 3640 2269 3641
rect 2399 3640 2400 3641
rect 2279 3642 2280 3643
rect 2454 3642 2455 3643
rect 2285 3644 2286 3645
rect 2343 3644 2344 3645
rect 2120 3646 2121 3647
rect 2286 3646 2287 3647
rect 2120 3648 2121 3649
rect 2301 3648 2302 3649
rect 2295 3650 2296 3651
rect 2297 3650 2298 3651
rect 2307 3650 2308 3651
rect 2447 3650 2448 3651
rect 2312 3652 2313 3653
rect 2319 3652 2320 3653
rect 2303 3654 2304 3655
rect 2313 3654 2314 3655
rect 2324 3654 2325 3655
rect 2535 3654 2536 3655
rect 2330 3656 2331 3657
rect 2523 3656 2524 3657
rect 2331 3658 2332 3659
rect 2396 3658 2397 3659
rect 2334 3660 2335 3661
rect 2393 3660 2394 3661
rect 2337 3662 2338 3663
rect 2471 3662 2472 3663
rect 2349 3664 2350 3665
rect 2477 3664 2478 3665
rect 2351 3666 2352 3667
rect 2457 3666 2458 3667
rect 2357 3668 2358 3669
rect 2541 3668 2542 3669
rect 2361 3670 2362 3671
rect 2411 3670 2412 3671
rect 2379 3672 2380 3673
rect 2667 3672 2668 3673
rect 2385 3674 2386 3675
rect 2519 3674 2520 3675
rect 2397 3676 2398 3677
rect 2537 3676 2538 3677
rect 2403 3678 2404 3679
rect 2423 3678 2424 3679
rect 2424 3680 2425 3681
rect 2528 3680 2529 3681
rect 2439 3682 2440 3683
rect 2495 3682 2496 3683
rect 2174 3684 2175 3685
rect 2496 3684 2497 3685
rect 2175 3686 2176 3687
rect 2451 3686 2452 3687
rect 2463 3686 2464 3687
rect 2737 3686 2738 3687
rect 2465 3688 2466 3689
rect 2585 3688 2586 3689
rect 2474 3690 2475 3691
rect 2559 3690 2560 3691
rect 2487 3692 2488 3693
rect 2612 3692 2613 3693
rect 2499 3694 2500 3695
rect 2603 3694 2604 3695
rect 2501 3696 2502 3697
rect 2598 3696 2599 3697
rect 2502 3698 2503 3699
rect 2606 3698 2607 3699
rect 2504 3700 2505 3701
rect 2601 3700 2602 3701
rect 2363 3702 2364 3703
rect 2505 3702 2506 3703
rect 2507 3702 2508 3703
rect 2511 3702 2512 3703
rect 2529 3702 2530 3703
rect 2670 3702 2671 3703
rect 2543 3704 2544 3705
rect 2689 3704 2690 3705
rect 2546 3706 2547 3707
rect 2589 3706 2590 3707
rect 2549 3708 2550 3709
rect 2776 3708 2777 3709
rect 2553 3710 2554 3711
rect 2752 3710 2753 3711
rect 2555 3712 2556 3713
rect 2686 3712 2687 3713
rect 2571 3714 2572 3715
rect 2591 3714 2592 3715
rect 2583 3716 2584 3717
rect 2633 3716 2634 3717
rect 2586 3718 2587 3719
rect 2692 3718 2693 3719
rect 2604 3720 2605 3721
rect 2639 3720 2640 3721
rect 2627 3722 2628 3723
rect 2661 3722 2662 3723
rect 2628 3724 2629 3725
rect 2664 3724 2665 3725
rect 2630 3726 2631 3727
rect 2778 3726 2779 3727
rect 2631 3728 2632 3729
rect 2657 3728 2658 3729
rect 2636 3730 2637 3731
rect 2818 3730 2819 3731
rect 2427 3732 2428 3733
rect 2818 3732 2819 3733
rect 2640 3734 2641 3735
rect 2645 3734 2646 3735
rect 2489 3736 2490 3737
rect 2646 3736 2647 3737
rect 2441 3738 2442 3739
rect 2490 3738 2491 3739
rect 2643 3738 2644 3739
rect 2648 3738 2649 3739
rect 2492 3740 2493 3741
rect 2649 3740 2650 3741
rect 2264 3742 2265 3743
rect 2493 3742 2494 3743
rect 2265 3744 2266 3745
rect 2408 3744 2409 3745
rect 2409 3746 2410 3747
rect 2752 3746 2753 3747
rect 2658 3748 2659 3749
rect 2808 3748 2809 3749
rect 2673 3750 2674 3751
rect 2716 3750 2717 3751
rect 2677 3752 2678 3753
rect 2683 3752 2684 3753
rect 2609 3754 2610 3755
rect 2677 3754 2678 3755
rect 2610 3756 2611 3757
rect 2734 3756 2735 3757
rect 2680 3758 2681 3759
rect 2801 3758 2802 3759
rect 2695 3760 2696 3761
rect 2758 3760 2759 3761
rect 2701 3762 2702 3763
rect 2815 3762 2816 3763
rect 2707 3764 2708 3765
rect 2811 3764 2812 3765
rect 2707 3766 2708 3767
rect 2773 3766 2774 3767
rect 2710 3768 2711 3769
rect 2713 3768 2714 3769
rect 2713 3770 2714 3771
rect 2728 3770 2729 3771
rect 2722 3772 2723 3773
rect 2725 3772 2726 3773
rect 2734 3772 2735 3773
rect 2790 3772 2791 3773
rect 2737 3774 2738 3775
rect 2746 3774 2747 3775
rect 2743 3776 2744 3777
rect 2787 3776 2788 3777
rect 2421 3778 2422 3779
rect 2787 3778 2788 3779
rect 2743 3780 2744 3781
rect 2767 3780 2768 3781
rect 2481 3782 2482 3783
rect 2768 3782 2769 3783
rect 2746 3784 2747 3785
rect 2770 3784 2771 3785
rect 2755 3786 2756 3787
rect 2761 3786 2762 3787
rect 2567 3788 2568 3789
rect 2761 3788 2762 3789
rect 2764 3788 2765 3789
rect 2783 3788 2784 3789
rect 2680 3790 2681 3791
rect 2764 3790 2765 3791
rect 2749 3792 2750 3793
rect 2784 3792 2785 3793
rect 2525 3794 2526 3795
rect 2749 3794 2750 3795
rect 2781 3794 2782 3795
rect 2811 3794 2812 3795
rect 2815 3794 2816 3795
rect 2832 3794 2833 3795
rect 2038 3803 2039 3804
rect 2123 3803 2124 3804
rect 2042 3805 2043 3806
rect 2126 3805 2127 3806
rect 2059 3807 2060 3808
rect 2235 3807 2236 3808
rect 2068 3809 2069 3810
rect 2225 3809 2226 3810
rect 2077 3811 2078 3812
rect 2229 3811 2230 3812
rect 2087 3813 2088 3814
rect 2250 3813 2251 3814
rect 2089 3815 2090 3816
rect 2216 3815 2217 3816
rect 2091 3817 2092 3818
rect 2112 3817 2113 3818
rect 2100 3819 2101 3820
rect 2283 3819 2284 3820
rect 2124 3821 2125 3822
rect 2339 3821 2340 3822
rect 2129 3823 2130 3824
rect 2241 3823 2242 3824
rect 2072 3825 2073 3826
rect 2240 3825 2241 3826
rect 2132 3827 2133 3828
rect 2258 3827 2259 3828
rect 2139 3829 2140 3830
rect 2313 3829 2314 3830
rect 2120 3831 2121 3832
rect 2312 3831 2313 3832
rect 2141 3833 2142 3834
rect 2355 3833 2356 3834
rect 2172 3835 2173 3836
rect 2598 3835 2599 3836
rect 2175 3837 2176 3838
rect 2334 3837 2335 3838
rect 2174 3839 2175 3840
rect 2178 3839 2179 3840
rect 2180 3839 2181 3840
rect 2238 3839 2239 3840
rect 2184 3841 2185 3842
rect 2337 3841 2338 3842
rect 2187 3843 2188 3844
rect 2262 3843 2263 3844
rect 2192 3845 2193 3846
rect 2496 3845 2497 3846
rect 2196 3847 2197 3848
rect 2234 3847 2235 3848
rect 2075 3849 2076 3850
rect 2195 3849 2196 3850
rect 2199 3849 2200 3850
rect 2210 3849 2211 3850
rect 2198 3851 2199 3852
rect 2208 3851 2209 3852
rect 2205 3853 2206 3854
rect 2237 3853 2238 3854
rect 2190 3855 2191 3856
rect 2204 3855 2205 3856
rect 2214 3855 2215 3856
rect 2529 3855 2530 3856
rect 2228 3857 2229 3858
rect 2454 3857 2455 3858
rect 2246 3859 2247 3860
rect 2373 3859 2374 3860
rect 2268 3861 2269 3862
rect 2297 3861 2298 3862
rect 2080 3863 2081 3864
rect 2267 3863 2268 3864
rect 2079 3865 2080 3866
rect 2220 3865 2221 3866
rect 2271 3865 2272 3866
rect 2559 3865 2560 3866
rect 2265 3867 2266 3868
rect 2270 3867 2271 3868
rect 2274 3867 2275 3868
rect 2516 3867 2517 3868
rect 2273 3869 2274 3870
rect 2343 3869 2344 3870
rect 2277 3871 2278 3872
rect 2309 3871 2310 3872
rect 2279 3873 2280 3874
rect 2286 3873 2287 3874
rect 2256 3875 2257 3876
rect 2285 3875 2286 3876
rect 2289 3875 2290 3876
rect 2315 3875 2316 3876
rect 2295 3877 2296 3878
rect 2303 3877 2304 3878
rect 2253 3879 2254 3880
rect 2294 3879 2295 3880
rect 2223 3881 2224 3882
rect 2252 3881 2253 3882
rect 2301 3881 2302 3882
rect 2345 3881 2346 3882
rect 2094 3883 2095 3884
rect 2300 3883 2301 3884
rect 2093 3885 2094 3886
rect 2222 3885 2223 3886
rect 2307 3885 2308 3886
rect 2333 3885 2334 3886
rect 2319 3887 2320 3888
rect 2321 3887 2322 3888
rect 2292 3889 2293 3890
rect 2318 3889 2319 3890
rect 2117 3891 2118 3892
rect 2291 3891 2292 3892
rect 2327 3891 2328 3892
rect 2349 3891 2350 3892
rect 2348 3893 2349 3894
rect 2376 3893 2377 3894
rect 2351 3895 2352 3896
rect 2535 3895 2536 3896
rect 2354 3897 2355 3898
rect 2493 3897 2494 3898
rect 2357 3899 2358 3900
rect 2451 3899 2452 3900
rect 2372 3901 2373 3902
rect 2457 3901 2458 3902
rect 2385 3903 2386 3904
rect 2727 3903 2728 3904
rect 2390 3905 2391 3906
rect 2764 3905 2765 3906
rect 2397 3907 2398 3908
rect 2815 3907 2816 3908
rect 2396 3909 2397 3910
rect 2403 3909 2404 3910
rect 2379 3911 2380 3912
rect 2402 3911 2403 3912
rect 2409 3911 2410 3912
rect 2617 3911 2618 3912
rect 2414 3913 2415 3914
rect 2601 3913 2602 3914
rect 2417 3915 2418 3916
rect 2505 3915 2506 3916
rect 2424 3917 2425 3918
rect 2749 3917 2750 3918
rect 2429 3919 2430 3920
rect 2752 3919 2753 3920
rect 2432 3921 2433 3922
rect 2686 3921 2687 3922
rect 2427 3923 2428 3924
rect 2686 3923 2687 3924
rect 2421 3925 2422 3926
rect 2426 3925 2427 3926
rect 2439 3925 2440 3926
rect 2771 3925 2772 3926
rect 2438 3927 2439 3928
rect 2463 3927 2464 3928
rect 2456 3929 2457 3930
rect 2490 3929 2491 3930
rect 2462 3931 2463 3932
rect 2655 3931 2656 3932
rect 2474 3933 2475 3934
rect 2502 3933 2503 3934
rect 2492 3935 2493 3936
rect 2511 3935 2512 3936
rect 2499 3937 2500 3938
rect 2513 3937 2514 3938
rect 2481 3939 2482 3940
rect 2498 3939 2499 3940
rect 2480 3941 2481 3942
rect 2523 3941 2524 3942
rect 2510 3943 2511 3944
rect 2801 3943 2802 3944
rect 2528 3945 2529 3946
rect 2628 3945 2629 3946
rect 2531 3947 2532 3948
rect 2631 3947 2632 3948
rect 2534 3949 2535 3950
rect 2586 3949 2587 3950
rect 2537 3951 2538 3952
rect 2571 3951 2572 3952
rect 2487 3953 2488 3954
rect 2570 3953 2571 3954
rect 2486 3955 2487 3956
rect 2541 3955 2542 3956
rect 2543 3955 2544 3956
rect 2640 3955 2641 3956
rect 2546 3957 2547 3958
rect 2601 3957 2602 3958
rect 2549 3959 2550 3960
rect 2553 3959 2554 3960
rect 2567 3959 2568 3960
rect 2677 3959 2678 3960
rect 2573 3961 2574 3962
rect 2604 3961 2605 3962
rect 2583 3963 2584 3964
rect 2692 3963 2693 3964
rect 2585 3965 2586 3966
rect 2646 3965 2647 3966
rect 2589 3967 2590 3968
rect 2689 3967 2690 3968
rect 2588 3969 2589 3970
rect 2649 3969 2650 3970
rect 2604 3971 2605 3972
rect 2811 3971 2812 3972
rect 2610 3973 2611 3974
rect 2668 3973 2669 3974
rect 2610 3975 2611 3976
rect 2734 3975 2735 3976
rect 2331 3977 2332 3978
rect 2734 3977 2735 3978
rect 2623 3979 2624 3980
rect 2658 3979 2659 3980
rect 2626 3981 2627 3982
rect 2661 3981 2662 3982
rect 2643 3983 2644 3984
rect 2673 3983 2674 3984
rect 2647 3985 2648 3986
rect 2707 3985 2708 3986
rect 2650 3987 2651 3988
rect 2710 3987 2711 3988
rect 2653 3989 2654 3990
rect 2720 3989 2721 3990
rect 2665 3991 2666 3992
rect 2731 3991 2732 3992
rect 2450 3993 2451 3994
rect 2730 3993 2731 3994
rect 2683 3995 2684 3996
rect 2808 3995 2809 3996
rect 2683 3997 2684 3998
rect 2743 3997 2744 3998
rect 2689 3999 2690 4000
rect 2794 3999 2795 4000
rect 2695 4001 2696 4002
rect 2775 4001 2776 4002
rect 2701 4003 2702 4004
rect 2755 4003 2756 4004
rect 2704 4005 2705 4006
rect 2758 4005 2759 4006
rect 2707 4007 2708 4008
rect 2713 4007 2714 4008
rect 2710 4009 2711 4010
rect 2716 4009 2717 4010
rect 2635 4011 2636 4012
rect 2716 4011 2717 4012
rect 2737 4011 2738 4012
rect 2763 4011 2764 4012
rect 2740 4013 2741 4014
rect 2781 4013 2782 4014
rect 2743 4015 2744 4016
rect 2784 4015 2785 4016
rect 2746 4017 2747 4018
rect 2787 4017 2788 4018
rect 2698 4019 2699 4020
rect 2746 4019 2747 4020
rect 2056 4028 2057 4029
rect 2267 4028 2268 4029
rect 2082 4030 2083 4031
rect 2285 4030 2286 4031
rect 2083 4032 2084 4033
rect 2291 4032 2292 4033
rect 2087 4034 2088 4035
rect 2163 4034 2164 4035
rect 2089 4036 2090 4037
rect 2300 4036 2301 4037
rect 2097 4038 2098 4039
rect 2127 4038 2128 4039
rect 2100 4040 2101 4041
rect 2385 4040 2386 4041
rect 2103 4042 2104 4043
rect 2318 4042 2319 4043
rect 2104 4044 2105 4045
rect 2312 4044 2313 4045
rect 2079 4046 2080 4047
rect 2313 4046 2314 4047
rect 2080 4048 2081 4049
rect 2094 4048 2095 4049
rect 2112 4048 2113 4049
rect 2370 4048 2371 4049
rect 2119 4050 2120 4051
rect 2315 4050 2316 4051
rect 2122 4052 2123 4053
rect 2343 4052 2344 4053
rect 2129 4054 2130 4055
rect 2222 4054 2223 4055
rect 2131 4056 2132 4057
rect 2303 4056 2304 4057
rect 2133 4058 2134 4059
rect 2246 4058 2247 4059
rect 2138 4060 2139 4061
rect 2339 4060 2340 4061
rect 2141 4062 2142 4063
rect 2345 4062 2346 4063
rect 2148 4064 2149 4065
rect 2340 4064 2341 4065
rect 2157 4066 2158 4067
rect 2193 4066 2194 4067
rect 2189 4068 2190 4069
rect 2265 4068 2266 4069
rect 2068 4070 2069 4071
rect 2190 4070 2191 4071
rect 2198 4070 2199 4071
rect 2202 4070 2203 4071
rect 2195 4072 2196 4073
rect 2199 4072 2200 4073
rect 2204 4072 2205 4073
rect 2208 4072 2209 4073
rect 2210 4072 2211 4073
rect 2214 4072 2215 4073
rect 2216 4072 2217 4073
rect 2220 4072 2221 4073
rect 2225 4072 2226 4073
rect 2388 4072 2389 4073
rect 2226 4074 2227 4075
rect 2546 4074 2547 4075
rect 2228 4076 2229 4077
rect 2304 4076 2305 4077
rect 2231 4078 2232 4079
rect 2357 4078 2358 4079
rect 2234 4080 2235 4081
rect 2268 4080 2269 4081
rect 2237 4082 2238 4083
rect 2301 4082 2302 4083
rect 2240 4084 2241 4085
rect 2244 4084 2245 4085
rect 2252 4084 2253 4085
rect 2346 4084 2347 4085
rect 2256 4086 2257 4087
rect 2421 4086 2422 4087
rect 2258 4088 2259 4089
rect 2406 4088 2407 4089
rect 2261 4090 2262 4091
rect 2480 4090 2481 4091
rect 2262 4092 2263 4093
rect 2354 4092 2355 4093
rect 2076 4094 2077 4095
rect 2355 4094 2356 4095
rect 2270 4096 2271 4097
rect 2358 4096 2359 4097
rect 2271 4098 2272 4099
rect 2273 4098 2274 4099
rect 2277 4098 2278 4099
rect 2321 4098 2322 4099
rect 2279 4100 2280 4101
rect 2376 4100 2377 4101
rect 2294 4102 2295 4103
rect 2316 4102 2317 4103
rect 2295 4104 2296 4105
rect 2486 4104 2487 4105
rect 2319 4106 2320 4107
rect 2372 4106 2373 4107
rect 2309 4108 2310 4109
rect 2373 4108 2374 4109
rect 2325 4110 2326 4111
rect 2516 4110 2517 4111
rect 2330 4112 2331 4113
rect 2583 4112 2584 4113
rect 2331 4114 2332 4115
rect 2417 4114 2418 4115
rect 2337 4116 2338 4117
rect 2351 4116 2352 4117
rect 2348 4118 2349 4119
rect 2418 4118 2419 4119
rect 2360 4120 2361 4121
rect 2379 4120 2380 4121
rect 2366 4122 2367 4123
rect 2594 4122 2595 4123
rect 2297 4124 2298 4125
rect 2367 4124 2368 4125
rect 2390 4124 2391 4125
rect 2478 4124 2479 4125
rect 2391 4126 2392 4127
rect 2528 4126 2529 4127
rect 2394 4128 2395 4129
rect 2531 4128 2532 4129
rect 2396 4130 2397 4131
rect 2409 4130 2410 4131
rect 2402 4132 2403 4133
rect 2490 4132 2491 4133
rect 2126 4134 2127 4135
rect 2403 4134 2404 4135
rect 2429 4134 2430 4135
rect 2502 4134 2503 4135
rect 2438 4136 2439 4137
rect 2610 4136 2611 4137
rect 2450 4138 2451 4139
rect 2520 4138 2521 4139
rect 2451 4140 2452 4141
rect 2543 4140 2544 4141
rect 2454 4142 2455 4143
rect 2534 4142 2535 4143
rect 2460 4144 2461 4145
rect 2567 4144 2568 4145
rect 2466 4146 2467 4147
rect 2585 4146 2586 4147
rect 2414 4148 2415 4149
rect 2586 4148 2587 4149
rect 2333 4150 2334 4151
rect 2415 4150 2416 4151
rect 2469 4150 2470 4151
rect 2588 4150 2589 4151
rect 2492 4152 2493 4153
rect 2718 4152 2719 4153
rect 2508 4154 2509 4155
rect 2730 4154 2731 4155
rect 2505 4156 2506 4157
rect 2731 4156 2732 4157
rect 2510 4158 2511 4159
rect 2568 4158 2569 4159
rect 2513 4160 2514 4161
rect 2773 4160 2774 4161
rect 2432 4162 2433 4163
rect 2514 4162 2515 4163
rect 2433 4164 2434 4165
rect 2637 4164 2638 4165
rect 2537 4166 2538 4167
rect 2544 4166 2545 4167
rect 2462 4168 2463 4169
rect 2538 4168 2539 4169
rect 2463 4170 2464 4171
rect 2570 4170 2571 4171
rect 2474 4172 2475 4173
rect 2571 4172 2572 4173
rect 2549 4174 2550 4175
rect 2595 4174 2596 4175
rect 2550 4176 2551 4177
rect 2573 4176 2574 4177
rect 2498 4178 2499 4179
rect 2574 4178 2575 4179
rect 2426 4180 2427 4181
rect 2499 4180 2500 4181
rect 2427 4182 2428 4183
rect 2456 4182 2457 4183
rect 2457 4184 2458 4185
rect 2617 4184 2618 4185
rect 2562 4186 2563 4187
rect 2668 4186 2669 4187
rect 2580 4188 2581 4189
rect 2692 4188 2693 4189
rect 2598 4190 2599 4191
rect 2613 4190 2614 4191
rect 2238 4192 2239 4193
rect 2613 4192 2614 4193
rect 2601 4194 2602 4195
rect 2781 4194 2782 4195
rect 2623 4196 2624 4197
rect 2755 4196 2756 4197
rect 2445 4198 2446 4199
rect 2622 4198 2623 4199
rect 2643 4198 2644 4199
rect 2753 4198 2754 4199
rect 2647 4200 2648 4201
rect 2673 4200 2674 4201
rect 2646 4202 2647 4203
rect 2767 4202 2768 4203
rect 2650 4204 2651 4205
rect 2727 4204 2728 4205
rect 2653 4206 2654 4207
rect 2713 4206 2714 4207
rect 2652 4208 2653 4209
rect 2676 4208 2677 4209
rect 2655 4210 2656 4211
rect 2724 4210 2725 4211
rect 2679 4212 2680 4213
rect 2743 4212 2744 4213
rect 2689 4214 2690 4215
rect 2760 4214 2761 4215
rect 2691 4216 2692 4217
rect 2707 4216 2708 4217
rect 2695 4218 2696 4219
rect 2749 4218 2750 4219
rect 2526 4220 2527 4221
rect 2748 4220 2749 4221
rect 2635 4222 2636 4223
rect 2694 4222 2695 4223
rect 2701 4222 2702 4223
rect 2721 4222 2722 4223
rect 2686 4224 2687 4225
rect 2700 4224 2701 4225
rect 2704 4224 2705 4225
rect 2777 4224 2778 4225
rect 2665 4226 2666 4227
rect 2703 4226 2704 4227
rect 2710 4226 2711 4227
rect 2716 4226 2717 4227
rect 2484 4228 2485 4229
rect 2715 4228 2716 4229
rect 2698 4230 2699 4231
rect 2709 4230 2710 4231
rect 2683 4232 2684 4233
rect 2697 4232 2698 4233
rect 2604 4234 2605 4235
rect 2682 4234 2683 4235
rect 2712 4234 2713 4235
rect 2734 4234 2735 4235
rect 2626 4236 2627 4237
rect 2734 4236 2735 4237
rect 2740 4236 2741 4237
rect 2780 4236 2781 4237
rect 2706 4238 2707 4239
rect 2741 4238 2742 4239
rect 2044 4247 2045 4248
rect 2190 4247 2191 4248
rect 2059 4249 2060 4250
rect 2087 4249 2088 4250
rect 2063 4251 2064 4252
rect 2268 4251 2269 4252
rect 2067 4253 2068 4254
rect 2199 4253 2200 4254
rect 2069 4255 2070 4256
rect 2206 4255 2207 4256
rect 2074 4257 2075 4258
rect 2233 4257 2234 4258
rect 2076 4259 2077 4260
rect 2083 4259 2084 4260
rect 2084 4261 2085 4262
rect 2293 4261 2294 4262
rect 2095 4263 2096 4264
rect 2365 4263 2366 4264
rect 2097 4265 2098 4266
rect 2388 4265 2389 4266
rect 2098 4267 2099 4268
rect 2403 4267 2404 4268
rect 2104 4269 2105 4270
rect 2311 4269 2312 4270
rect 2107 4271 2108 4272
rect 2116 4271 2117 4272
rect 2113 4273 2114 4274
rect 2373 4273 2374 4274
rect 2129 4275 2130 4276
rect 2353 4275 2354 4276
rect 2133 4277 2134 4278
rect 2415 4277 2416 4278
rect 2135 4279 2136 4280
rect 2275 4279 2276 4280
rect 2142 4281 2143 4282
rect 2202 4281 2203 4282
rect 2070 4283 2071 4284
rect 2203 4283 2204 4284
rect 2148 4285 2149 4286
rect 2271 4285 2272 4286
rect 2157 4287 2158 4288
rect 2316 4287 2317 4288
rect 2160 4289 2161 4290
rect 2265 4289 2266 4290
rect 2163 4291 2164 4292
rect 2317 4291 2318 4292
rect 2166 4293 2167 4294
rect 2284 4293 2285 4294
rect 2181 4295 2182 4296
rect 2188 4295 2189 4296
rect 2193 4295 2194 4296
rect 2226 4295 2227 4296
rect 2214 4297 2215 4298
rect 2227 4297 2228 4298
rect 2215 4299 2216 4300
rect 2220 4299 2221 4300
rect 2208 4301 2209 4302
rect 2221 4301 2222 4302
rect 2238 4301 2239 4302
rect 2325 4301 2326 4302
rect 2244 4303 2245 4304
rect 2254 4303 2255 4304
rect 2245 4305 2246 4306
rect 2301 4305 2302 4306
rect 2248 4307 2249 4308
rect 2626 4307 2627 4308
rect 2256 4309 2257 4310
rect 2370 4309 2371 4310
rect 2241 4311 2242 4312
rect 2371 4311 2372 4312
rect 2119 4313 2120 4314
rect 2242 4313 2243 4314
rect 2272 4313 2273 4314
rect 2406 4313 2407 4314
rect 2290 4315 2291 4316
rect 2313 4315 2314 4316
rect 2299 4317 2300 4318
rect 2418 4317 2419 4318
rect 2302 4319 2303 4320
rect 2355 4319 2356 4320
rect 2308 4321 2309 4322
rect 2376 4321 2377 4322
rect 2314 4323 2315 4324
rect 2367 4323 2368 4324
rect 2326 4325 2327 4326
rect 2385 4325 2386 4326
rect 2323 4327 2324 4328
rect 2386 4327 2387 4328
rect 2335 4329 2336 4330
rect 2343 4329 2344 4330
rect 2340 4331 2341 4332
rect 2356 4331 2357 4332
rect 2304 4333 2305 4334
rect 2341 4333 2342 4334
rect 2305 4335 2306 4336
rect 2358 4335 2359 4336
rect 2319 4337 2320 4338
rect 2359 4337 2360 4338
rect 2262 4339 2263 4340
rect 2320 4339 2321 4340
rect 2368 4339 2369 4340
rect 2718 4339 2719 4340
rect 2377 4341 2378 4342
rect 2445 4341 2446 4342
rect 2389 4343 2390 4344
rect 2409 4343 2410 4344
rect 2401 4345 2402 4346
rect 2586 4345 2587 4346
rect 2413 4347 2414 4348
rect 2478 4347 2479 4348
rect 2419 4349 2420 4350
rect 2484 4349 2485 4350
rect 2425 4351 2426 4352
rect 2490 4351 2491 4352
rect 2427 4353 2428 4354
rect 2637 4353 2638 4354
rect 2433 4355 2434 4356
rect 2437 4355 2438 4356
rect 2449 4355 2450 4356
rect 2514 4355 2515 4356
rect 2451 4357 2452 4358
rect 2530 4357 2531 4358
rect 2457 4359 2458 4360
rect 2619 4359 2620 4360
rect 2229 4361 2230 4362
rect 2620 4361 2621 4362
rect 2463 4363 2464 4364
rect 2640 4363 2641 4364
rect 2466 4365 2467 4366
rect 2617 4365 2618 4366
rect 2469 4367 2470 4368
rect 2518 4367 2519 4368
rect 2491 4369 2492 4370
rect 2796 4369 2797 4370
rect 2497 4371 2498 4372
rect 2684 4371 2685 4372
rect 2508 4373 2509 4374
rect 2512 4373 2513 4374
rect 2509 4375 2510 4376
rect 2571 4375 2572 4376
rect 2520 4377 2521 4378
rect 2745 4377 2746 4378
rect 2421 4379 2422 4380
rect 2745 4379 2746 4380
rect 2533 4381 2534 4382
rect 2574 4381 2575 4382
rect 2542 4383 2543 4384
rect 2652 4383 2653 4384
rect 2550 4385 2551 4386
rect 2605 4385 2606 4386
rect 2544 4387 2545 4388
rect 2551 4387 2552 4388
rect 2545 4389 2546 4390
rect 2649 4389 2650 4390
rect 2460 4391 2461 4392
rect 2650 4391 2651 4392
rect 2295 4393 2296 4394
rect 2461 4393 2462 4394
rect 2277 4395 2278 4396
rect 2296 4395 2297 4396
rect 2562 4395 2563 4396
rect 2599 4395 2600 4396
rect 2563 4397 2564 4398
rect 2595 4397 2596 4398
rect 2568 4399 2569 4400
rect 2773 4399 2774 4400
rect 2569 4401 2570 4402
rect 2580 4401 2581 4402
rect 2394 4403 2395 4404
rect 2581 4403 2582 4404
rect 2331 4405 2332 4406
rect 2395 4405 2396 4406
rect 2575 4405 2576 4406
rect 2601 4405 2602 4406
rect 2587 4407 2588 4408
rect 2687 4407 2688 4408
rect 2593 4409 2594 4410
rect 2738 4409 2739 4410
rect 2610 4411 2611 4412
rect 2622 4411 2623 4412
rect 2583 4413 2584 4414
rect 2623 4413 2624 4414
rect 2391 4415 2392 4416
rect 2584 4415 2585 4416
rect 2613 4415 2614 4416
rect 2668 4415 2669 4416
rect 2646 4417 2647 4418
rect 2755 4417 2756 4418
rect 2647 4419 2648 4420
rect 2734 4419 2735 4420
rect 2655 4421 2656 4422
rect 2665 4421 2666 4422
rect 2673 4421 2674 4422
rect 2727 4421 2728 4422
rect 2676 4423 2677 4424
rect 2724 4423 2725 4424
rect 2526 4425 2527 4426
rect 2723 4425 2724 4426
rect 2694 4427 2695 4428
rect 2741 4427 2742 4428
rect 2499 4429 2500 4430
rect 2742 4429 2743 4430
rect 2500 4431 2501 4432
rect 2505 4431 2506 4432
rect 2682 4431 2683 4432
rect 2693 4431 2694 4432
rect 2703 4431 2704 4432
rect 2726 4431 2727 4432
rect 2702 4433 2703 4434
rect 2785 4433 2786 4434
rect 2706 4435 2707 4436
rect 2729 4435 2730 4436
rect 2643 4437 2644 4438
rect 2705 4437 2706 4438
rect 2712 4437 2713 4438
rect 2756 4437 2757 4438
rect 2700 4439 2701 4440
rect 2711 4439 2712 4440
rect 2699 4441 2700 4442
rect 2715 4441 2716 4442
rect 2278 4443 2279 4444
rect 2714 4443 2715 4444
rect 2762 4443 2763 4444
rect 2766 4443 2767 4444
rect 2731 4445 2732 4446
rect 2763 4445 2764 4446
rect 2721 4447 2722 4448
rect 2732 4447 2733 4448
rect 2709 4449 2710 4450
rect 2720 4449 2721 4450
rect 2697 4451 2698 4452
rect 2708 4451 2709 4452
rect 2691 4453 2692 4454
rect 2696 4453 2697 4454
rect 2679 4455 2680 4456
rect 2690 4455 2691 4456
rect 2379 4457 2380 4458
rect 2680 4457 2681 4458
rect 2769 4457 2770 4458
rect 2787 4457 2788 4458
rect 2769 4459 2770 4460
rect 2776 4459 2777 4460
rect 2772 4461 2773 4462
rect 2782 4461 2783 4462
rect 2053 4470 2054 4471
rect 2060 4470 2061 4471
rect 2056 4472 2057 4473
rect 2188 4472 2189 4473
rect 2063 4474 2064 4475
rect 2199 4474 2200 4475
rect 2070 4476 2071 4477
rect 2206 4476 2207 4477
rect 2074 4478 2075 4479
rect 2227 4478 2228 4479
rect 2074 4480 2075 4481
rect 2299 4480 2300 4481
rect 2077 4482 2078 4483
rect 2221 4482 2222 4483
rect 2081 4484 2082 4485
rect 2193 4484 2194 4485
rect 2084 4486 2085 4487
rect 2272 4486 2273 4487
rect 2088 4488 2089 4489
rect 2311 4488 2312 4489
rect 2088 4490 2089 4491
rect 2205 4490 2206 4491
rect 2091 4492 2092 4493
rect 2335 4492 2336 4493
rect 2095 4494 2096 4495
rect 2302 4494 2303 4495
rect 2098 4496 2099 4497
rect 2254 4496 2255 4497
rect 2100 4498 2101 4499
rect 2107 4498 2108 4499
rect 2113 4498 2114 4499
rect 2135 4498 2136 4499
rect 2113 4500 2114 4501
rect 2317 4500 2318 4501
rect 2116 4502 2117 4503
rect 2296 4502 2297 4503
rect 2120 4504 2121 4505
rect 2308 4504 2309 4505
rect 2123 4506 2124 4507
rect 2256 4506 2257 4507
rect 2123 4508 2124 4509
rect 2290 4508 2291 4509
rect 2133 4510 2134 4511
rect 2157 4510 2158 4511
rect 2142 4512 2143 4513
rect 2176 4512 2177 4513
rect 2151 4514 2152 4515
rect 2356 4514 2357 4515
rect 2157 4516 2158 4517
rect 2203 4516 2204 4517
rect 2160 4518 2161 4519
rect 2245 4518 2246 4519
rect 2163 4520 2164 4521
rect 2353 4520 2354 4521
rect 2166 4522 2167 4523
rect 2251 4522 2252 4523
rect 2166 4524 2167 4525
rect 2233 4524 2234 4525
rect 2169 4526 2170 4527
rect 2305 4526 2306 4527
rect 2173 4528 2174 4529
rect 2284 4528 2285 4529
rect 2184 4530 2185 4531
rect 2275 4530 2276 4531
rect 2187 4532 2188 4533
rect 2371 4532 2372 4533
rect 2190 4534 2191 4535
rect 2271 4534 2272 4535
rect 2196 4536 2197 4537
rect 2293 4536 2294 4537
rect 2202 4538 2203 4539
rect 2338 4538 2339 4539
rect 2211 4540 2212 4541
rect 2283 4540 2284 4541
rect 2215 4542 2216 4543
rect 2220 4542 2221 4543
rect 2217 4544 2218 4545
rect 2314 4544 2315 4545
rect 2229 4546 2230 4547
rect 2278 4546 2279 4547
rect 2235 4548 2236 4549
rect 2326 4548 2327 4549
rect 2238 4550 2239 4551
rect 2320 4550 2321 4551
rect 2242 4552 2243 4553
rect 2629 4552 2630 4553
rect 2241 4554 2242 4555
rect 2323 4554 2324 4555
rect 2250 4556 2251 4557
rect 2684 4556 2685 4557
rect 2253 4558 2254 4559
rect 2347 4558 2348 4559
rect 2259 4560 2260 4561
rect 2341 4560 2342 4561
rect 2265 4562 2266 4563
rect 2365 4562 2366 4563
rect 2274 4564 2275 4565
rect 2368 4564 2369 4565
rect 2277 4566 2278 4567
rect 2359 4566 2360 4567
rect 2289 4568 2290 4569
rect 2386 4568 2387 4569
rect 2295 4570 2296 4571
rect 2389 4570 2390 4571
rect 2307 4572 2308 4573
rect 2749 4572 2750 4573
rect 2313 4574 2314 4575
rect 2687 4574 2688 4575
rect 2325 4576 2326 4577
rect 2413 4576 2414 4577
rect 2331 4578 2332 4579
rect 2680 4578 2681 4579
rect 2343 4580 2344 4581
rect 2699 4580 2700 4581
rect 2349 4582 2350 4583
rect 2461 4582 2462 4583
rect 2355 4584 2356 4585
rect 2437 4584 2438 4585
rect 2361 4586 2362 4587
rect 2449 4586 2450 4587
rect 2367 4588 2368 4589
rect 2455 4588 2456 4589
rect 2377 4590 2378 4591
rect 2383 4590 2384 4591
rect 2379 4592 2380 4593
rect 2711 4592 2712 4593
rect 2385 4594 2386 4595
rect 2745 4594 2746 4595
rect 2397 4596 2398 4597
rect 2723 4596 2724 4597
rect 2401 4598 2402 4599
rect 2641 4598 2642 4599
rect 2409 4600 2410 4601
rect 2491 4600 2492 4601
rect 2415 4602 2416 4603
rect 2503 4602 2504 4603
rect 2419 4604 2420 4605
rect 2608 4604 2609 4605
rect 2433 4606 2434 4607
rect 2497 4606 2498 4607
rect 2436 4608 2437 4609
rect 2500 4608 2501 4609
rect 2445 4610 2446 4611
rect 2581 4610 2582 4611
rect 2301 4612 2302 4613
rect 2580 4612 2581 4613
rect 2448 4614 2449 4615
rect 2584 4614 2585 4615
rect 2451 4616 2452 4617
rect 2533 4616 2534 4617
rect 2457 4618 2458 4619
rect 2530 4618 2531 4619
rect 2460 4620 2461 4621
rect 2679 4620 2680 4621
rect 2463 4622 2464 4623
rect 2539 4622 2540 4623
rect 2466 4624 2467 4625
rect 2542 4624 2543 4625
rect 2469 4626 2470 4627
rect 2551 4626 2552 4627
rect 2475 4628 2476 4629
rect 2545 4628 2546 4629
rect 2395 4630 2396 4631
rect 2544 4630 2545 4631
rect 2478 4632 2479 4633
rect 2512 4632 2513 4633
rect 2487 4634 2488 4635
rect 2617 4634 2618 4635
rect 2490 4636 2491 4637
rect 2620 4636 2621 4637
rect 2493 4638 2494 4639
rect 2563 4638 2564 4639
rect 2499 4640 2500 4641
rect 2569 4640 2570 4641
rect 2505 4642 2506 4643
rect 2593 4642 2594 4643
rect 2509 4644 2510 4645
rect 2538 4644 2539 4645
rect 2511 4646 2512 4647
rect 2715 4646 2716 4647
rect 2518 4648 2519 4649
rect 2805 4648 2806 4649
rect 2523 4650 2524 4651
rect 2599 4650 2600 4651
rect 2529 4652 2530 4653
rect 2759 4652 2760 4653
rect 2535 4654 2536 4655
rect 2789 4654 2790 4655
rect 2541 4656 2542 4657
rect 2547 4656 2548 4657
rect 2550 4656 2551 4657
rect 2623 4656 2624 4657
rect 2568 4658 2569 4659
rect 2650 4658 2651 4659
rect 2583 4660 2584 4661
rect 2665 4660 2666 4661
rect 2425 4662 2426 4663
rect 2665 4662 2666 4663
rect 2589 4664 2590 4665
rect 2729 4664 2730 4665
rect 2575 4666 2576 4667
rect 2729 4666 2730 4667
rect 2601 4668 2602 4669
rect 2647 4668 2648 4669
rect 2605 4670 2606 4671
rect 2735 4670 2736 4671
rect 2565 4672 2566 4673
rect 2604 4672 2605 4673
rect 2614 4672 2615 4673
rect 2690 4672 2691 4673
rect 2617 4674 2618 4675
rect 2693 4674 2694 4675
rect 2620 4676 2621 4677
rect 2696 4676 2697 4677
rect 2626 4678 2627 4679
rect 2644 4678 2645 4679
rect 2626 4680 2627 4681
rect 2720 4680 2721 4681
rect 2638 4682 2639 4683
rect 2799 4682 2800 4683
rect 2641 4684 2642 4685
rect 2708 4684 2709 4685
rect 2650 4686 2651 4687
rect 2732 4686 2733 4687
rect 2659 4688 2660 4689
rect 2785 4688 2786 4689
rect 2662 4690 2663 4691
rect 2726 4690 2727 4691
rect 2672 4692 2673 4693
rect 2705 4692 2706 4693
rect 2699 4694 2700 4695
rect 2769 4694 2770 4695
rect 2702 4696 2703 4697
rect 2766 4696 2767 4697
rect 2587 4698 2588 4699
rect 2702 4698 2703 4699
rect 2586 4700 2587 4701
rect 2668 4700 2669 4701
rect 2623 4702 2624 4703
rect 2668 4702 2669 4703
rect 2705 4702 2706 4703
rect 2772 4702 2773 4703
rect 2060 4711 2061 4712
rect 2225 4711 2226 4712
rect 2074 4713 2075 4714
rect 2191 4713 2192 4714
rect 2077 4715 2078 4716
rect 2188 4715 2189 4716
rect 2081 4717 2082 4718
rect 2166 4717 2167 4718
rect 2093 4719 2094 4720
rect 2100 4719 2101 4720
rect 2106 4719 2107 4720
rect 2235 4719 2236 4720
rect 2084 4721 2085 4722
rect 2105 4721 2106 4722
rect 2084 4723 2085 4724
rect 2133 4723 2134 4724
rect 2109 4725 2110 4726
rect 2234 4725 2235 4726
rect 2108 4727 2109 4728
rect 2125 4727 2126 4728
rect 2113 4729 2114 4730
rect 2141 4729 2142 4730
rect 2116 4731 2117 4732
rect 2157 4731 2158 4732
rect 2130 4733 2131 4734
rect 2289 4733 2290 4734
rect 2138 4735 2139 4736
rect 2207 4735 2208 4736
rect 2151 4737 2152 4738
rect 2295 4737 2296 4738
rect 2152 4739 2153 4740
rect 2184 4739 2185 4740
rect 2154 4741 2155 4742
rect 2466 4741 2467 4742
rect 2158 4743 2159 4744
rect 2169 4743 2170 4744
rect 2164 4745 2165 4746
rect 2241 4745 2242 4746
rect 2067 4747 2068 4748
rect 2240 4747 2241 4748
rect 2067 4749 2068 4750
rect 2182 4749 2183 4750
rect 2193 4749 2194 4750
rect 2243 4749 2244 4750
rect 2167 4751 2168 4752
rect 2194 4751 2195 4752
rect 2196 4751 2197 4752
rect 2246 4751 2247 4752
rect 2211 4753 2212 4754
rect 2620 4753 2621 4754
rect 2214 4755 2215 4756
rect 2650 4755 2651 4756
rect 2217 4757 2218 4758
rect 2261 4757 2262 4758
rect 2229 4759 2230 4760
rect 2288 4759 2289 4760
rect 2202 4761 2203 4762
rect 2228 4761 2229 4762
rect 2238 4761 2239 4762
rect 2285 4761 2286 4762
rect 2199 4763 2200 4764
rect 2237 4763 2238 4764
rect 2253 4763 2254 4764
rect 2303 4763 2304 4764
rect 2112 4765 2113 4766
rect 2252 4765 2253 4766
rect 2256 4765 2257 4766
rect 2297 4765 2298 4766
rect 2205 4767 2206 4768
rect 2255 4767 2256 4768
rect 2259 4767 2260 4768
rect 2580 4767 2581 4768
rect 2265 4769 2266 4770
rect 2318 4769 2319 4770
rect 2220 4771 2221 4772
rect 2264 4771 2265 4772
rect 2063 4773 2064 4774
rect 2219 4773 2220 4774
rect 2274 4773 2275 4774
rect 2321 4773 2322 4774
rect 2279 4775 2280 4776
rect 2643 4775 2644 4776
rect 2283 4777 2284 4778
rect 2550 4777 2551 4778
rect 2309 4779 2310 4780
rect 2490 4779 2491 4780
rect 2325 4781 2326 4782
rect 2647 4781 2648 4782
rect 2277 4783 2278 4784
rect 2324 4783 2325 4784
rect 2331 4783 2332 4784
rect 2372 4783 2373 4784
rect 2330 4785 2331 4786
rect 2349 4785 2350 4786
rect 2313 4787 2314 4788
rect 2348 4787 2349 4788
rect 2271 4789 2272 4790
rect 2312 4789 2313 4790
rect 2343 4789 2344 4790
rect 2715 4789 2716 4790
rect 2307 4791 2308 4792
rect 2342 4791 2343 4792
rect 2361 4791 2362 4792
rect 2390 4791 2391 4792
rect 2367 4793 2368 4794
rect 2402 4793 2403 4794
rect 2397 4795 2398 4796
rect 2712 4795 2713 4796
rect 2415 4797 2416 4798
rect 2429 4797 2430 4798
rect 2379 4799 2380 4800
rect 2414 4799 2415 4800
rect 2355 4801 2356 4802
rect 2378 4801 2379 4802
rect 2301 4803 2302 4804
rect 2354 4803 2355 4804
rect 2250 4805 2251 4806
rect 2300 4805 2301 4806
rect 2120 4807 2121 4808
rect 2249 4807 2250 4808
rect 2417 4807 2418 4808
rect 2445 4807 2446 4808
rect 2420 4809 2421 4810
rect 2448 4809 2449 4810
rect 2436 4811 2437 4812
rect 2438 4811 2439 4812
rect 2433 4813 2434 4814
rect 2435 4813 2436 4814
rect 2441 4813 2442 4814
rect 2457 4813 2458 4814
rect 2444 4815 2445 4816
rect 2460 4815 2461 4816
rect 2451 4817 2452 4818
rect 2465 4817 2466 4818
rect 2453 4819 2454 4820
rect 2478 4819 2479 4820
rect 2459 4821 2460 4822
rect 2463 4821 2464 4822
rect 2462 4823 2463 4824
rect 2577 4823 2578 4824
rect 2469 4825 2470 4826
rect 2477 4825 2478 4826
rect 2471 4827 2472 4828
rect 2568 4827 2569 4828
rect 2475 4829 2476 4830
rect 2483 4829 2484 4830
rect 2487 4829 2488 4830
rect 2507 4829 2508 4830
rect 2493 4831 2494 4832
rect 2576 4831 2577 4832
rect 2495 4833 2496 4834
rect 2668 4833 2669 4834
rect 2499 4835 2500 4836
rect 2519 4835 2520 4836
rect 2505 4837 2506 4838
rect 2513 4837 2514 4838
rect 2511 4839 2512 4840
rect 2531 4839 2532 4840
rect 2306 4841 2307 4842
rect 2510 4841 2511 4842
rect 2523 4841 2524 4842
rect 2708 4841 2709 4842
rect 2529 4843 2530 4844
rect 2693 4843 2694 4844
rect 2535 4845 2536 4846
rect 2555 4845 2556 4846
rect 2538 4847 2539 4848
rect 2558 4847 2559 4848
rect 2544 4849 2545 4850
rect 2612 4849 2613 4850
rect 2543 4851 2544 4852
rect 2547 4851 2548 4852
rect 2541 4853 2542 4854
rect 2546 4853 2547 4854
rect 2567 4853 2568 4854
rect 2629 4853 2630 4854
rect 2573 4855 2574 4856
rect 2617 4855 2618 4856
rect 2579 4857 2580 4858
rect 2604 4857 2605 4858
rect 2589 4859 2590 4860
rect 2594 4859 2595 4860
rect 2586 4861 2587 4862
rect 2588 4861 2589 4862
rect 2583 4863 2584 4864
rect 2585 4863 2586 4864
rect 2565 4865 2566 4866
rect 2582 4865 2583 4866
rect 2591 4865 2592 4866
rect 2708 4865 2709 4866
rect 2606 4867 2607 4868
rect 2623 4867 2624 4868
rect 2360 4869 2361 4870
rect 2624 4869 2625 4870
rect 2614 4871 2615 4872
rect 2729 4871 2730 4872
rect 2618 4873 2619 4874
rect 2696 4873 2697 4874
rect 2626 4875 2627 4876
rect 2652 4875 2653 4876
rect 2636 4877 2637 4878
rect 2672 4877 2673 4878
rect 2498 4879 2499 4880
rect 2673 4879 2674 4880
rect 2638 4881 2639 4882
rect 2736 4881 2737 4882
rect 2641 4883 2642 4884
rect 2733 4883 2734 4884
rect 2409 4885 2410 4886
rect 2734 4885 2735 4886
rect 2385 4887 2386 4888
rect 2408 4887 2409 4888
rect 2649 4887 2650 4888
rect 2694 4887 2695 4888
rect 2659 4889 2660 4890
rect 2667 4889 2668 4890
rect 2609 4891 2610 4892
rect 2658 4891 2659 4892
rect 2662 4891 2663 4892
rect 2687 4891 2688 4892
rect 2670 4893 2671 4894
rect 2690 4893 2691 4894
rect 2699 4893 2700 4894
rect 2714 4893 2715 4894
rect 2702 4895 2703 4896
rect 2717 4895 2718 4896
rect 2726 4895 2727 4896
rect 2737 4895 2738 4896
rect 2053 4904 2054 4905
rect 2225 4904 2226 4905
rect 2060 4906 2061 4907
rect 2240 4906 2241 4907
rect 2063 4908 2064 4909
rect 2164 4908 2165 4909
rect 2066 4910 2067 4911
rect 2188 4910 2189 4911
rect 2070 4912 2071 4913
rect 2237 4912 2238 4913
rect 2069 4914 2070 4915
rect 2081 4914 2082 4915
rect 2074 4916 2075 4917
rect 2182 4916 2183 4917
rect 2077 4918 2078 4919
rect 2191 4918 2192 4919
rect 2076 4920 2077 4921
rect 2080 4920 2081 4921
rect 2083 4920 2084 4921
rect 2200 4920 2201 4921
rect 2095 4922 2096 4923
rect 2246 4922 2247 4923
rect 2105 4924 2106 4925
rect 2234 4924 2235 4925
rect 2108 4926 2109 4927
rect 2264 4926 2265 4927
rect 2115 4928 2116 4929
rect 2255 4928 2256 4929
rect 2119 4930 2120 4931
rect 2234 4930 2235 4931
rect 2122 4932 2123 4933
rect 2243 4932 2244 4933
rect 2125 4934 2126 4935
rect 2138 4934 2139 4935
rect 2134 4936 2135 4937
rect 2207 4936 2208 4937
rect 2135 4938 2136 4939
rect 2158 4938 2159 4939
rect 2141 4940 2142 4941
rect 2151 4940 2152 4941
rect 2141 4942 2142 4943
rect 2396 4942 2397 4943
rect 2155 4944 2156 4945
rect 2324 4944 2325 4945
rect 2155 4946 2156 4947
rect 2285 4946 2286 4947
rect 2158 4948 2159 4949
rect 2279 4948 2280 4949
rect 2161 4950 2162 4951
rect 2219 4950 2220 4951
rect 2170 4952 2171 4953
rect 2216 4952 2217 4953
rect 2179 4954 2180 4955
rect 2228 4954 2229 4955
rect 2185 4956 2186 4957
rect 2249 4956 2250 4957
rect 2188 4958 2189 4959
rect 2252 4958 2253 4959
rect 2197 4960 2198 4961
rect 2387 4960 2388 4961
rect 2197 4962 2198 4963
rect 2261 4962 2262 4963
rect 2204 4964 2205 4965
rect 2579 4964 2580 4965
rect 2222 4966 2223 4967
rect 2288 4966 2289 4967
rect 2231 4968 2232 4969
rect 2297 4968 2298 4969
rect 2243 4970 2244 4971
rect 2300 4970 2301 4971
rect 2246 4972 2247 4973
rect 2303 4972 2304 4973
rect 2255 4974 2256 4975
rect 2318 4974 2319 4975
rect 2261 4976 2262 4977
rect 2330 4976 2331 4977
rect 2273 4978 2274 4979
rect 2360 4978 2361 4979
rect 2279 4980 2280 4981
rect 2615 4980 2616 4981
rect 2285 4982 2286 4983
rect 2348 4982 2349 4983
rect 2303 4984 2304 4985
rect 2372 4984 2373 4985
rect 2309 4986 2310 4987
rect 2378 4986 2379 4987
rect 2315 4988 2316 4989
rect 2599 4988 2600 4989
rect 2321 4990 2322 4991
rect 2399 4990 2400 4991
rect 2321 4992 2322 4993
rect 2390 4992 2391 4993
rect 2327 4994 2328 4995
rect 2444 4994 2445 4995
rect 2342 4996 2343 4997
rect 2549 4996 2550 4997
rect 2345 4998 2346 4999
rect 2408 4998 2409 4999
rect 2351 5000 2352 5001
rect 2414 5000 2415 5001
rect 2354 5002 2355 5003
rect 2580 5002 2581 5003
rect 2366 5004 2367 5005
rect 2429 5004 2430 5005
rect 2372 5006 2373 5007
rect 2435 5006 2436 5007
rect 2375 5008 2376 5009
rect 2438 5008 2439 5009
rect 2378 5010 2379 5011
rect 2616 5010 2617 5011
rect 2384 5012 2385 5013
rect 2558 5012 2559 5013
rect 2390 5014 2391 5015
rect 2459 5014 2460 5015
rect 2393 5016 2394 5017
rect 2680 5016 2681 5017
rect 2402 5018 2403 5019
rect 2737 5018 2738 5019
rect 2408 5020 2409 5021
rect 2477 5020 2478 5021
rect 2432 5022 2433 5023
rect 2495 5022 2496 5023
rect 2435 5024 2436 5025
rect 2498 5024 2499 5025
rect 2438 5026 2439 5027
rect 2576 5026 2577 5027
rect 2441 5028 2442 5029
rect 2444 5028 2445 5029
rect 2441 5030 2442 5031
rect 2465 5030 2466 5031
rect 2420 5032 2421 5033
rect 2465 5032 2466 5033
rect 2420 5034 2421 5035
rect 2483 5034 2484 5035
rect 2447 5036 2448 5037
rect 2552 5036 2553 5037
rect 2453 5038 2454 5039
rect 2701 5038 2702 5039
rect 2456 5040 2457 5041
rect 2519 5040 2520 5041
rect 2462 5042 2463 5043
rect 2646 5042 2647 5043
rect 2417 5044 2418 5045
rect 2462 5044 2463 5045
rect 2468 5044 2469 5045
rect 2727 5044 2728 5045
rect 2471 5046 2472 5047
rect 2519 5046 2520 5047
rect 2474 5048 2475 5049
rect 2531 5048 2532 5049
rect 2486 5050 2487 5051
rect 2507 5050 2508 5051
rect 2297 5052 2298 5053
rect 2507 5052 2508 5053
rect 2489 5054 2490 5055
rect 2510 5054 2511 5055
rect 2492 5056 2493 5057
rect 2546 5056 2547 5057
rect 2495 5058 2496 5059
rect 2571 5058 2572 5059
rect 2510 5060 2511 5061
rect 2567 5060 2568 5061
rect 2513 5062 2514 5063
rect 2624 5062 2625 5063
rect 2516 5064 2517 5065
rect 2582 5064 2583 5065
rect 2522 5066 2523 5067
rect 2585 5066 2586 5067
rect 2525 5068 2526 5069
rect 2588 5068 2589 5069
rect 2528 5070 2529 5071
rect 2591 5070 2592 5071
rect 2531 5072 2532 5073
rect 2620 5072 2621 5073
rect 2546 5074 2547 5075
rect 2609 5074 2610 5075
rect 2555 5076 2556 5077
rect 2642 5076 2643 5077
rect 2543 5078 2544 5079
rect 2556 5078 2557 5079
rect 2312 5080 2313 5081
rect 2543 5080 2544 5081
rect 2562 5080 2563 5081
rect 2618 5080 2619 5081
rect 2565 5082 2566 5083
rect 2594 5082 2595 5083
rect 2586 5084 2587 5085
rect 2649 5084 2650 5085
rect 2589 5086 2590 5087
rect 2652 5086 2653 5087
rect 2592 5088 2593 5089
rect 2670 5088 2671 5089
rect 2606 5090 2607 5091
rect 2655 5090 2656 5091
rect 2573 5092 2574 5093
rect 2606 5092 2607 5093
rect 2627 5092 2628 5093
rect 2639 5092 2640 5093
rect 2626 5094 2627 5095
rect 2720 5094 2721 5095
rect 2629 5096 2630 5097
rect 2717 5096 2718 5097
rect 2667 5098 2668 5099
rect 2690 5098 2691 5099
rect 2714 5098 2715 5099
rect 2723 5098 2724 5099
rect 2054 5107 2055 5108
rect 2161 5107 2162 5108
rect 2057 5109 2058 5110
rect 2119 5109 2120 5110
rect 2062 5111 2063 5112
rect 2164 5111 2165 5112
rect 2071 5113 2072 5114
rect 2135 5113 2136 5114
rect 2078 5115 2079 5116
rect 2092 5115 2093 5116
rect 2081 5117 2082 5118
rect 2095 5117 2096 5118
rect 2098 5117 2099 5118
rect 2200 5117 2201 5118
rect 2101 5119 2102 5120
rect 2197 5119 2198 5120
rect 2102 5121 2103 5122
rect 2114 5121 2115 5122
rect 2105 5123 2106 5124
rect 2131 5123 2132 5124
rect 2111 5125 2112 5126
rect 2185 5125 2186 5126
rect 2122 5127 2123 5128
rect 2138 5127 2139 5128
rect 2126 5129 2127 5130
rect 2144 5129 2145 5130
rect 2128 5131 2129 5132
rect 2275 5131 2276 5132
rect 2137 5133 2138 5134
rect 2151 5133 2152 5134
rect 2141 5135 2142 5136
rect 2234 5135 2235 5136
rect 2144 5137 2145 5138
rect 2516 5137 2517 5138
rect 2155 5139 2156 5140
rect 2586 5139 2587 5140
rect 2167 5141 2168 5142
rect 2399 5141 2400 5142
rect 2167 5143 2168 5144
rect 2179 5143 2180 5144
rect 2170 5145 2171 5146
rect 2396 5145 2397 5146
rect 2170 5147 2171 5148
rect 2188 5147 2189 5148
rect 2191 5147 2192 5148
rect 2222 5147 2223 5148
rect 2200 5149 2201 5150
rect 2231 5149 2232 5150
rect 2203 5151 2204 5152
rect 2243 5151 2244 5152
rect 2206 5153 2207 5154
rect 2246 5153 2247 5154
rect 2210 5155 2211 5156
rect 2281 5155 2282 5156
rect 2148 5157 2149 5158
rect 2209 5157 2210 5158
rect 2216 5157 2217 5158
rect 2218 5157 2219 5158
rect 2215 5159 2216 5160
rect 2255 5159 2256 5160
rect 2221 5161 2222 5162
rect 2261 5161 2262 5162
rect 2233 5163 2234 5164
rect 2279 5163 2280 5164
rect 2236 5165 2237 5166
rect 2465 5165 2466 5166
rect 2254 5167 2255 5168
rect 2303 5167 2304 5168
rect 2260 5169 2261 5170
rect 2327 5169 2328 5170
rect 2266 5171 2267 5172
rect 2602 5171 2603 5172
rect 2273 5173 2274 5174
rect 2552 5173 2553 5174
rect 2272 5175 2273 5176
rect 2462 5175 2463 5176
rect 2278 5177 2279 5178
rect 2486 5177 2487 5178
rect 2290 5179 2291 5180
rect 2321 5179 2322 5180
rect 2297 5181 2298 5182
rect 2540 5181 2541 5182
rect 2296 5183 2297 5184
rect 2595 5183 2596 5184
rect 2302 5185 2303 5186
rect 2345 5185 2346 5186
rect 2309 5187 2310 5188
rect 2571 5187 2572 5188
rect 2308 5189 2309 5190
rect 2568 5189 2569 5190
rect 2329 5191 2330 5192
rect 2384 5191 2385 5192
rect 2338 5193 2339 5194
rect 2606 5193 2607 5194
rect 2344 5195 2345 5196
rect 2387 5195 2388 5196
rect 2347 5197 2348 5198
rect 2444 5197 2445 5198
rect 2359 5199 2360 5200
rect 2432 5199 2433 5200
rect 2362 5201 2363 5202
rect 2366 5201 2367 5202
rect 2372 5201 2373 5202
rect 2497 5201 2498 5202
rect 2371 5203 2372 5204
rect 2592 5203 2593 5204
rect 2375 5205 2376 5206
rect 2485 5205 2486 5206
rect 2285 5207 2286 5208
rect 2374 5207 2375 5208
rect 2284 5209 2285 5210
rect 2315 5209 2316 5210
rect 2314 5211 2315 5212
rect 2351 5211 2352 5212
rect 2350 5213 2351 5214
rect 2447 5213 2448 5214
rect 2378 5215 2379 5216
rect 2609 5215 2610 5216
rect 2377 5217 2378 5218
rect 2456 5217 2457 5218
rect 2383 5219 2384 5220
rect 2438 5219 2439 5220
rect 2386 5221 2387 5222
rect 2457 5221 2458 5222
rect 2390 5223 2391 5224
rect 2556 5223 2557 5224
rect 2393 5225 2394 5226
rect 2424 5225 2425 5226
rect 2392 5227 2393 5228
rect 2642 5227 2643 5228
rect 2408 5229 2409 5230
rect 2433 5229 2434 5230
rect 2410 5231 2411 5232
rect 2549 5231 2550 5232
rect 2420 5233 2421 5234
rect 2515 5233 2516 5234
rect 2257 5235 2258 5236
rect 2420 5235 2421 5236
rect 2430 5235 2431 5236
rect 2522 5235 2523 5236
rect 2441 5237 2442 5238
rect 2543 5237 2544 5238
rect 2442 5239 2443 5240
rect 2546 5239 2547 5240
rect 2445 5241 2446 5242
rect 2460 5241 2461 5242
rect 2454 5243 2455 5244
rect 2528 5243 2529 5244
rect 2464 5245 2465 5246
rect 2525 5245 2526 5246
rect 2468 5247 2469 5248
rect 2529 5247 2530 5248
rect 2470 5249 2471 5250
rect 2562 5249 2563 5250
rect 2476 5251 2477 5252
rect 2632 5251 2633 5252
rect 2479 5253 2480 5254
rect 2629 5253 2630 5254
rect 2489 5255 2490 5256
rect 2504 5255 2505 5256
rect 2488 5257 2489 5258
rect 2589 5257 2590 5258
rect 2495 5259 2496 5260
rect 2507 5259 2508 5260
rect 2492 5261 2493 5262
rect 2494 5261 2495 5262
rect 2491 5263 2492 5264
rect 2510 5263 2511 5264
rect 2482 5265 2483 5266
rect 2511 5265 2512 5266
rect 2519 5265 2520 5266
rect 2536 5265 2537 5266
rect 2435 5267 2436 5268
rect 2518 5267 2519 5268
rect 2531 5267 2532 5268
rect 2613 5267 2614 5268
rect 2474 5269 2475 5270
rect 2532 5269 2533 5270
rect 2473 5271 2474 5272
rect 2565 5271 2566 5272
rect 2620 5271 2621 5272
rect 2626 5271 2627 5272
rect 2047 5280 2048 5281
rect 2119 5280 2120 5281
rect 2074 5282 2075 5283
rect 2092 5282 2093 5283
rect 2075 5284 2076 5285
rect 2122 5284 2123 5285
rect 2079 5286 2080 5287
rect 2085 5286 2086 5287
rect 2082 5288 2083 5289
rect 2089 5288 2090 5289
rect 2092 5288 2093 5289
rect 2099 5288 2100 5289
rect 2102 5288 2103 5289
rect 2170 5288 2171 5289
rect 2106 5290 2107 5291
rect 2218 5290 2219 5291
rect 2113 5292 2114 5293
rect 2134 5292 2135 5293
rect 2116 5294 2117 5295
rect 2196 5294 2197 5295
rect 2119 5296 2120 5297
rect 2151 5296 2152 5297
rect 2122 5298 2123 5299
rect 2128 5298 2129 5299
rect 2128 5300 2129 5301
rect 2131 5300 2132 5301
rect 2131 5302 2132 5303
rect 2141 5302 2142 5303
rect 2138 5304 2139 5305
rect 2226 5304 2227 5305
rect 2148 5306 2149 5307
rect 2163 5306 2164 5307
rect 2155 5308 2156 5309
rect 2221 5308 2222 5309
rect 2157 5310 2158 5311
rect 2272 5310 2273 5311
rect 2167 5312 2168 5313
rect 2175 5312 2176 5313
rect 2169 5314 2170 5315
rect 2209 5314 2210 5315
rect 2203 5316 2204 5317
rect 2208 5316 2209 5317
rect 2206 5318 2207 5319
rect 2211 5318 2212 5319
rect 2215 5318 2216 5319
rect 2223 5318 2224 5319
rect 2200 5320 2201 5321
rect 2214 5320 2215 5321
rect 2191 5322 2192 5323
rect 2199 5322 2200 5323
rect 2217 5322 2218 5323
rect 2247 5322 2248 5323
rect 2229 5324 2230 5325
rect 2278 5324 2279 5325
rect 2233 5326 2234 5327
rect 2244 5326 2245 5327
rect 2238 5328 2239 5329
rect 2275 5328 2276 5329
rect 2241 5330 2242 5331
rect 2281 5330 2282 5331
rect 2254 5332 2255 5333
rect 2286 5332 2287 5333
rect 2257 5334 2258 5335
rect 2508 5334 2509 5335
rect 2260 5336 2261 5337
rect 2410 5336 2411 5337
rect 2259 5338 2260 5339
rect 2374 5338 2375 5339
rect 2266 5340 2267 5341
rect 2277 5340 2278 5341
rect 2265 5342 2266 5343
rect 2350 5342 2351 5343
rect 2271 5344 2272 5345
rect 2402 5344 2403 5345
rect 2296 5346 2297 5347
rect 2331 5346 2332 5347
rect 2302 5348 2303 5349
rect 2546 5348 2547 5349
rect 2308 5350 2309 5351
rect 2334 5350 2335 5351
rect 2290 5352 2291 5353
rect 2307 5352 2308 5353
rect 2289 5354 2290 5355
rect 2511 5354 2512 5355
rect 2314 5356 2315 5357
rect 2522 5356 2523 5357
rect 2319 5358 2320 5359
rect 2398 5358 2399 5359
rect 2322 5360 2323 5361
rect 2347 5360 2348 5361
rect 2325 5362 2326 5363
rect 2362 5362 2363 5363
rect 2338 5364 2339 5365
rect 2340 5364 2341 5365
rect 2344 5364 2345 5365
rect 2352 5364 2353 5365
rect 2359 5364 2360 5365
rect 2515 5364 2516 5365
rect 2368 5366 2369 5367
rect 2417 5366 2418 5367
rect 2367 5368 2368 5369
rect 2460 5368 2461 5369
rect 2371 5370 2372 5371
rect 2379 5370 2380 5371
rect 2370 5372 2371 5373
rect 2445 5372 2446 5373
rect 2386 5374 2387 5375
rect 2525 5374 2526 5375
rect 2383 5376 2384 5377
rect 2385 5376 2386 5377
rect 2382 5378 2383 5379
rect 2395 5378 2396 5379
rect 2388 5380 2389 5381
rect 2442 5380 2443 5381
rect 2392 5382 2393 5383
rect 2529 5382 2530 5383
rect 2414 5384 2415 5385
rect 2430 5384 2431 5385
rect 2417 5386 2418 5387
rect 2433 5386 2434 5387
rect 2420 5388 2421 5389
rect 2476 5388 2477 5389
rect 2313 5390 2314 5391
rect 2420 5390 2421 5391
rect 2427 5390 2428 5391
rect 2442 5390 2443 5391
rect 2430 5392 2431 5393
rect 2482 5392 2483 5393
rect 2329 5394 2330 5395
rect 2482 5394 2483 5395
rect 2328 5396 2329 5397
rect 2485 5396 2486 5397
rect 2433 5398 2434 5399
rect 2470 5398 2471 5399
rect 2436 5400 2437 5401
rect 2501 5400 2502 5401
rect 2445 5402 2446 5403
rect 2488 5402 2489 5403
rect 2448 5404 2449 5405
rect 2491 5404 2492 5405
rect 2454 5406 2455 5407
rect 2465 5406 2466 5407
rect 2473 5406 2474 5407
rect 2536 5406 2537 5407
rect 2284 5408 2285 5409
rect 2472 5408 2473 5409
rect 2283 5410 2284 5411
rect 2424 5410 2425 5411
rect 2377 5412 2378 5413
rect 2423 5412 2424 5413
rect 2479 5412 2480 5413
rect 2532 5412 2533 5413
rect 2491 5414 2492 5415
rect 2500 5414 2501 5415
rect 2494 5416 2495 5417
rect 2497 5416 2498 5417
rect 2065 5425 2066 5426
rect 2072 5425 2073 5426
rect 2079 5425 2080 5426
rect 2128 5425 2129 5426
rect 2099 5427 2100 5428
rect 2113 5427 2114 5428
rect 2106 5429 2107 5430
rect 2172 5429 2173 5430
rect 2111 5431 2112 5432
rect 2178 5431 2179 5432
rect 2115 5433 2116 5434
rect 2214 5433 2215 5434
rect 2119 5435 2120 5436
rect 2181 5435 2182 5436
rect 2125 5437 2126 5438
rect 2251 5437 2252 5438
rect 2127 5439 2128 5440
rect 2208 5439 2209 5440
rect 2131 5441 2132 5442
rect 2220 5441 2221 5442
rect 2130 5443 2131 5444
rect 2211 5443 2212 5444
rect 2141 5445 2142 5446
rect 2232 5445 2233 5446
rect 2145 5447 2146 5448
rect 2157 5447 2158 5448
rect 2138 5449 2139 5450
rect 2144 5449 2145 5450
rect 2148 5449 2149 5450
rect 2241 5449 2242 5450
rect 2151 5451 2152 5452
rect 2257 5451 2258 5452
rect 2163 5453 2164 5454
rect 2166 5453 2167 5454
rect 2175 5453 2176 5454
rect 2205 5453 2206 5454
rect 2196 5455 2197 5456
rect 2221 5455 2222 5456
rect 2118 5457 2119 5458
rect 2196 5457 2197 5458
rect 2223 5457 2224 5458
rect 2254 5457 2255 5458
rect 2199 5459 2200 5460
rect 2224 5459 2225 5460
rect 2184 5461 2185 5462
rect 2199 5461 2200 5462
rect 2169 5463 2170 5464
rect 2184 5463 2185 5464
rect 2229 5463 2230 5464
rect 2305 5463 2306 5464
rect 2238 5465 2239 5466
rect 2275 5465 2276 5466
rect 2247 5467 2248 5468
rect 2265 5467 2266 5468
rect 2248 5469 2249 5470
rect 2322 5469 2323 5470
rect 2134 5471 2135 5472
rect 2323 5471 2324 5472
rect 2259 5473 2260 5474
rect 2468 5473 2469 5474
rect 2260 5475 2261 5476
rect 2382 5475 2383 5476
rect 2218 5477 2219 5478
rect 2383 5477 2384 5478
rect 2277 5479 2278 5480
rect 2338 5479 2339 5480
rect 2215 5481 2216 5482
rect 2278 5481 2279 5482
rect 2283 5481 2284 5482
rect 2391 5481 2392 5482
rect 2284 5483 2285 5484
rect 2359 5483 2360 5484
rect 2286 5485 2287 5486
rect 2296 5485 2297 5486
rect 2287 5487 2288 5488
rect 2313 5487 2314 5488
rect 2289 5489 2290 5490
rect 2419 5489 2420 5490
rect 2307 5491 2308 5492
rect 2454 5491 2455 5492
rect 2244 5493 2245 5494
rect 2308 5493 2309 5494
rect 2245 5495 2246 5496
rect 2319 5495 2320 5496
rect 2317 5497 2318 5498
rect 2389 5497 2390 5498
rect 2328 5499 2329 5500
rect 2410 5499 2411 5500
rect 2271 5501 2272 5502
rect 2329 5501 2330 5502
rect 2235 5503 2236 5504
rect 2272 5503 2273 5504
rect 2347 5503 2348 5504
rect 2423 5503 2424 5504
rect 2352 5505 2353 5506
rect 2404 5505 2405 5506
rect 2370 5507 2371 5508
rect 2402 5507 2403 5508
rect 2374 5509 2375 5510
rect 2417 5509 2418 5510
rect 2379 5511 2380 5512
rect 2395 5511 2396 5512
rect 2380 5513 2381 5514
rect 2438 5513 2439 5514
rect 2385 5515 2386 5516
rect 2483 5515 2484 5516
rect 2365 5517 2366 5518
rect 2386 5517 2387 5518
rect 2407 5517 2408 5518
rect 2430 5517 2431 5518
rect 2340 5519 2341 5520
rect 2431 5519 2432 5520
rect 2341 5521 2342 5522
rect 2422 5521 2423 5522
rect 2414 5523 2415 5524
rect 2455 5523 2456 5524
rect 2413 5525 2414 5526
rect 2433 5525 2434 5526
rect 2353 5527 2354 5528
rect 2434 5527 2435 5528
rect 2416 5529 2417 5530
rect 2436 5529 2437 5530
rect 2425 5531 2426 5532
rect 2452 5531 2453 5532
rect 2428 5533 2429 5534
rect 2445 5533 2446 5534
rect 2367 5535 2368 5536
rect 2445 5535 2446 5536
rect 2441 5537 2442 5538
rect 2448 5537 2449 5538
rect 2325 5539 2326 5540
rect 2448 5539 2449 5540
rect 2326 5541 2327 5542
rect 2398 5541 2399 5542
rect 2331 5543 2332 5544
rect 2398 5543 2399 5544
rect 2476 5543 2477 5544
rect 2494 5543 2495 5544
rect 2487 5545 2488 5546
rect 2494 5545 2495 5546
rect 2491 5547 2492 5548
rect 2514 5547 2515 5548
rect 2500 5549 2501 5550
rect 2504 5549 2505 5550
rect 2089 5558 2090 5559
rect 2192 5558 2193 5559
rect 2092 5560 2093 5561
rect 2189 5560 2190 5561
rect 2101 5562 2102 5563
rect 2205 5562 2206 5563
rect 2111 5564 2112 5565
rect 2172 5564 2173 5565
rect 2104 5566 2105 5567
rect 2111 5566 2112 5567
rect 2118 5566 2119 5567
rect 2196 5566 2197 5567
rect 2132 5568 2133 5569
rect 2153 5568 2154 5569
rect 2134 5570 2135 5571
rect 2248 5570 2249 5571
rect 2137 5572 2138 5573
rect 2221 5572 2222 5573
rect 2141 5574 2142 5575
rect 2278 5574 2279 5575
rect 2148 5576 2149 5577
rect 2272 5576 2273 5577
rect 2159 5578 2160 5579
rect 2199 5578 2200 5579
rect 2162 5580 2163 5581
rect 2184 5580 2185 5581
rect 2166 5582 2167 5583
rect 2222 5582 2223 5583
rect 2171 5584 2172 5585
rect 2178 5584 2179 5585
rect 2174 5586 2175 5587
rect 2181 5586 2182 5587
rect 2183 5586 2184 5587
rect 2257 5586 2258 5587
rect 2195 5588 2196 5589
rect 2211 5588 2212 5589
rect 2198 5590 2199 5591
rect 2438 5590 2439 5591
rect 2204 5592 2205 5593
rect 2224 5592 2225 5593
rect 2208 5594 2209 5595
rect 2326 5594 2327 5595
rect 2144 5596 2145 5597
rect 2207 5596 2208 5597
rect 2216 5596 2217 5597
rect 2227 5596 2228 5597
rect 2225 5598 2226 5599
rect 2275 5598 2276 5599
rect 2228 5600 2229 5601
rect 2254 5600 2255 5601
rect 2231 5602 2232 5603
rect 2241 5602 2242 5603
rect 2233 5604 2234 5605
rect 2289 5604 2290 5605
rect 2234 5606 2235 5607
rect 2251 5606 2252 5607
rect 2236 5608 2237 5609
rect 2292 5608 2293 5609
rect 2237 5610 2238 5611
rect 2262 5610 2263 5611
rect 2247 5612 2248 5613
rect 2305 5612 2306 5613
rect 2245 5614 2246 5615
rect 2304 5614 2305 5615
rect 2284 5616 2285 5617
rect 2323 5616 2324 5617
rect 2283 5618 2284 5619
rect 2338 5618 2339 5619
rect 2287 5620 2288 5621
rect 2317 5620 2318 5621
rect 2286 5622 2287 5623
rect 2329 5622 2330 5623
rect 2296 5624 2297 5625
rect 2298 5624 2299 5625
rect 2260 5626 2261 5627
rect 2295 5626 2296 5627
rect 2259 5628 2260 5629
rect 2308 5628 2309 5629
rect 2307 5630 2308 5631
rect 2365 5630 2366 5631
rect 2310 5632 2311 5633
rect 2419 5632 2420 5633
rect 2322 5634 2323 5635
rect 2448 5634 2449 5635
rect 2325 5636 2326 5637
rect 2341 5636 2342 5637
rect 2335 5638 2336 5639
rect 2365 5638 2366 5639
rect 2340 5640 2341 5641
rect 2344 5640 2345 5641
rect 2347 5640 2348 5641
rect 2393 5640 2394 5641
rect 2350 5642 2351 5643
rect 2416 5642 2417 5643
rect 2353 5644 2354 5645
rect 2400 5644 2401 5645
rect 2356 5646 2357 5647
rect 2383 5646 2384 5647
rect 2359 5648 2360 5649
rect 2378 5648 2379 5649
rect 2359 5650 2360 5651
rect 2374 5650 2375 5651
rect 2369 5652 2370 5653
rect 2380 5652 2381 5653
rect 2372 5654 2373 5655
rect 2387 5654 2388 5655
rect 2375 5656 2376 5657
rect 2407 5656 2408 5657
rect 2390 5658 2391 5659
rect 2413 5658 2414 5659
rect 2404 5660 2405 5661
rect 2487 5660 2488 5661
rect 2406 5662 2407 5663
rect 2425 5662 2426 5663
rect 2410 5664 2411 5665
rect 2445 5664 2446 5665
rect 2428 5666 2429 5667
rect 2441 5666 2442 5667
rect 2473 5666 2474 5667
rect 2483 5666 2484 5667
rect 2089 5675 2090 5676
rect 2192 5675 2193 5676
rect 2092 5677 2093 5678
rect 2099 5677 2100 5678
rect 2104 5677 2105 5678
rect 2171 5677 2172 5678
rect 2096 5679 2097 5680
rect 2103 5679 2104 5680
rect 2106 5679 2107 5680
rect 2216 5679 2217 5680
rect 2108 5681 2109 5682
rect 2174 5681 2175 5682
rect 2109 5683 2110 5684
rect 2189 5683 2190 5684
rect 2115 5685 2116 5686
rect 2122 5685 2123 5686
rect 2118 5687 2119 5688
rect 2195 5687 2196 5688
rect 2125 5689 2126 5690
rect 2153 5689 2154 5690
rect 2126 5691 2127 5692
rect 2204 5691 2205 5692
rect 2129 5693 2130 5694
rect 2207 5693 2208 5694
rect 2138 5695 2139 5696
rect 2198 5695 2199 5696
rect 2141 5697 2142 5698
rect 2183 5697 2184 5698
rect 2132 5699 2133 5700
rect 2141 5699 2142 5700
rect 2144 5699 2145 5700
rect 2231 5699 2232 5700
rect 2144 5701 2145 5702
rect 2228 5701 2229 5702
rect 2151 5703 2152 5704
rect 2190 5703 2191 5704
rect 2154 5705 2155 5706
rect 2225 5705 2226 5706
rect 2157 5707 2158 5708
rect 2259 5707 2260 5708
rect 2163 5709 2164 5710
rect 2262 5709 2263 5710
rect 2172 5711 2173 5712
rect 2289 5711 2290 5712
rect 2181 5713 2182 5714
rect 2295 5713 2296 5714
rect 2184 5715 2185 5716
rect 2298 5715 2299 5716
rect 2193 5717 2194 5718
rect 2362 5717 2363 5718
rect 2196 5719 2197 5720
rect 2283 5719 2284 5720
rect 2205 5721 2206 5722
rect 2292 5721 2293 5722
rect 2208 5723 2209 5724
rect 2247 5723 2248 5724
rect 2211 5725 2212 5726
rect 2359 5725 2360 5726
rect 2222 5727 2223 5728
rect 2400 5727 2401 5728
rect 2221 5729 2222 5730
rect 2322 5729 2323 5730
rect 2228 5731 2229 5732
rect 2325 5731 2326 5732
rect 2234 5733 2235 5734
rect 2375 5733 2376 5734
rect 2237 5735 2238 5736
rect 2378 5735 2379 5736
rect 2244 5737 2245 5738
rect 2304 5737 2305 5738
rect 2246 5739 2247 5740
rect 2396 5739 2397 5740
rect 2249 5741 2250 5742
rect 2387 5741 2388 5742
rect 2255 5743 2256 5744
rect 2310 5743 2311 5744
rect 2262 5745 2263 5746
rect 2390 5745 2391 5746
rect 2286 5747 2287 5748
rect 2340 5747 2341 5748
rect 2307 5749 2308 5750
rect 2413 5749 2414 5750
rect 2350 5751 2351 5752
rect 2393 5751 2394 5752
rect 2356 5753 2357 5754
rect 2369 5753 2370 5754
rect 2065 5762 2066 5763
rect 2072 5762 2073 5763
rect 2089 5762 2090 5763
rect 2109 5762 2110 5763
rect 2119 5762 2120 5763
rect 2141 5762 2142 5763
rect 2122 5764 2123 5765
rect 2157 5764 2158 5765
rect 2126 5766 2127 5767
rect 2138 5766 2139 5767
rect 2147 5766 2148 5767
rect 2151 5766 2152 5767
rect 2153 5766 2154 5767
rect 2156 5766 2157 5767
rect 2159 5766 2160 5767
rect 2234 5766 2235 5767
rect 2166 5768 2167 5769
rect 2181 5768 2182 5769
rect 2169 5770 2170 5771
rect 2214 5770 2215 5771
rect 2172 5772 2173 5773
rect 2190 5772 2191 5773
rect 2184 5774 2185 5775
rect 2221 5774 2222 5775
rect 2193 5776 2194 5777
rect 2208 5776 2209 5777
rect 2196 5778 2197 5779
rect 2224 5778 2225 5779
rect 2211 5780 2212 5781
rect 2231 5780 2232 5781
rect 2237 5780 2238 5781
rect 2255 5780 2256 5781
rect 2246 5782 2247 5783
rect 2262 5782 2263 5783
rect 2249 5784 2250 5785
rect 2259 5784 2260 5785
rect 2146 5793 2147 5794
rect 2150 5793 2151 5794
rect 2156 5793 2157 5794
rect 2159 5793 2160 5794
rect 2143 5802 2144 5803
rect 2153 5802 2154 5803
<< end >>
