magic
tech scmos
timestamp 1395743079
<< m1p >>
use CELL  1
transform -1 0 1058 0 1 2363
box 0 0 6 6
use CELL  2
transform -1 0 1088 0 1 713
box 0 0 6 6
use CELL  3
transform 1 0 1475 0 1 1388
box 0 0 6 6
use CELL  4
transform -1 0 1086 0 1 1388
box 0 0 6 6
use CELL  5
transform -1 0 1356 0 1 1668
box 0 0 6 6
use CELL  6
transform -1 0 1042 0 1 713
box 0 0 6 6
use CELL  7
transform 1 0 1071 0 1 2449
box 0 0 6 6
use CELL  8
transform 1 0 1128 0 -1 512
box 0 0 6 6
use CELL  9
transform -1 0 1281 0 1 1936
box 0 0 6 6
use CELL  10
transform 1 0 1336 0 -1 719
box 0 0 6 6
use CELL  11
transform 1 0 1101 0 1 506
box 0 0 6 6
use CELL  12
transform -1 0 1172 0 1 2363
box 0 0 6 6
use CELL  13
transform 1 0 1346 0 1 1821
box 0 0 6 6
use CELL  14
transform 1 0 1137 0 1 2047
box 0 0 6 6
use CELL  15
transform -1 0 1393 0 1 1821
box 0 0 6 6
use CELL  16
transform -1 0 1300 0 1 1821
box 0 0 6 6
use CELL  17
transform 1 0 1272 0 1 620
box 0 0 6 6
use CELL  18
transform 1 0 1392 0 -1 818
box 0 0 6 6
use CELL  19
transform -1 0 1349 0 1 713
box 0 0 6 6
use CELL  20
transform -1 0 1026 0 1 2235
box 0 0 6 6
use CELL  21
transform 1 0 1431 0 1 1535
box 0 0 6 6
use CELL  22
transform -1 0 1398 0 1 1092
box 0 0 6 6
use CELL  23
transform -1 0 1218 0 1 557
box 0 0 6 6
use CELL  24
transform -1 0 1156 0 -1 2134
box 0 0 6 6
use CELL  25
transform 1 0 1442 0 1 959
box 0 0 6 6
use CELL  26
transform -1 0 1015 0 1 1668
box 0 0 6 6
use CELL  27
transform -1 0 1153 0 1 557
box 0 0 6 6
use CELL  28
transform 1 0 990 0 1 1388
box 0 0 6 6
use CELL  29
transform -1 0 1088 0 1 1668
box 0 0 6 6
use CELL  30
transform -1 0 1010 0 1 1388
box 0 0 6 6
use CELL  31
transform -1 0 1008 0 1 1253
box 0 0 6 6
use CELL  32
transform 1 0 1008 0 1 620
box 0 0 6 6
use CELL  33
transform -1 0 1462 0 1 959
box 0 0 6 6
use CELL  34
transform -1 0 1420 0 1 1092
box 0 0 6 6
use CELL  35
transform -1 0 960 0 1 959
box 0 0 6 6
use CELL  36
transform -1 0 1039 0 1 2300
box 0 0 6 6
use CELL  37
transform -1 0 1108 0 1 1821
box 0 0 6 6
use CELL  38
transform -1 0 1087 0 1 2128
box 0 0 6 6
use CELL  39
transform -1 0 1398 0 1 959
box 0 0 6 6
use CELL  40
transform -1 0 1224 0 1 2047
box 0 0 6 6
use CELL  41
transform -1 0 1071 0 1 2128
box 0 0 6 6
use CELL  42
transform 1 0 1235 0 1 620
box 0 0 6 6
use CELL  43
transform -1 0 1002 0 1 1535
box 0 0 6 6
use CELL  44
transform -1 0 1042 0 1 959
box 0 0 6 6
use CELL  45
transform 1 0 1071 0 1 1821
box 0 0 6 6
use CELL  46
transform -1 0 1059 0 1 1936
box 0 0 6 6
use CELL  47
transform -1 0 1382 0 1 1388
box 0 0 6 6
use CELL  48
transform 1 0 1276 0 1 2235
box 0 0 6 6
use CELL  49
transform -1 0 1021 0 1 1821
box 0 0 6 6
use CELL  50
transform 1 0 1345 0 -1 2053
box 0 0 6 6
use CELL  51
transform -1 0 1061 0 -1 719
box 0 0 6 6
use CELL  52
transform 1 0 1037 0 -1 2053
box 0 0 6 6
use CELL  53
transform -1 0 1073 0 -1 626
box 0 0 6 6
use CELL  54
transform -1 0 1339 0 1 1535
box 0 0 6 6
use CELL  55
transform -1 0 1412 0 1 812
box 0 0 6 6
use CELL  56
transform -1 0 1074 0 1 2235
box 0 0 6 6
use CELL  57
transform -1 0 1409 0 1 1535
box 0 0 6 6
use CELL  58
transform 1 0 1381 0 -1 1541
box 0 0 6 6
use CELL  59
transform -1 0 1399 0 -1 1827
box 0 0 6 6
use CELL  60
transform -1 0 1030 0 1 620
box 0 0 6 6
use CELL  61
transform 1 0 1058 0 1 2128
box 0 0 6 6
use CELL  62
transform -1 0 1333 0 1 1936
box 0 0 6 6
use CELL  63
transform 1 0 1420 0 1 812
box 0 0 6 6
use CELL  64
transform 1 0 1449 0 1 959
box 0 0 6 6
use CELL  65
transform -1 0 1022 0 1 1668
box 0 0 6 6
use CELL  66
transform -1 0 1026 0 1 506
box 0 0 6 6
use CELL  67
transform -1 0 1026 0 1 713
box 0 0 6 6
use CELL  68
transform -1 0 1188 0 1 1936
box 0 0 6 6
use CELL  69
transform 1 0 1089 0 1 1668
box 0 0 6 6
use CELL  70
transform -1 0 1083 0 1 1092
box 0 0 6 6
use CELL  71
transform -1 0 1427 0 1 1668
box 0 0 6 6
use CELL  72
transform -1 0 1036 0 1 1668
box 0 0 6 6
use CELL  73
transform -1 0 1014 0 1 1092
box 0 0 6 6
use CELL  74
transform 1 0 1021 0 1 812
box 0 0 6 6
use CELL  75
transform -1 0 1015 0 1 1253
box 0 0 6 6
use CELL  76
transform -1 0 1440 0 1 1668
box 0 0 6 6
use CELL  77
transform -1 0 1061 0 1 1821
box 0 0 6 6
use CELL  78
transform -1 0 1042 0 1 1092
box 0 0 6 6
use CELL  79
transform -1 0 1246 0 1 2047
box 0 0 6 6
use CELL  80
transform -1 0 1180 0 1 1535
box 0 0 6 6
use CELL  81
transform 1 0 1309 0 1 2047
box 0 0 6 6
use CELL  82
transform 1 0 1244 0 1 620
box 0 0 6 6
use CELL  83
transform -1 0 1046 0 1 2363
box 0 0 6 6
use CELL  84
transform -1 0 1433 0 1 1253
box 0 0 6 6
use CELL  85
transform -1 0 1052 0 1 2128
box 0 0 6 6
use CELL  86
transform -1 0 1066 0 1 620
box 0 0 6 6
use CELL  87
transform -1 0 1053 0 1 2300
box 0 0 6 6
use CELL  88
transform -1 0 1345 0 1 2047
box 0 0 6 6
use CELL  89
transform 1 0 1156 0 -1 563
box 0 0 6 6
use CELL  90
transform -1 0 1421 0 1 1253
box 0 0 6 6
use CELL  91
transform -1 0 1097 0 -1 818
box 0 0 6 6
use CELL  92
transform -1 0 1358 0 1 2047
box 0 0 6 6
use CELL  93
transform -1 0 1003 0 1 1388
box 0 0 6 6
use CELL  94
transform -1 0 1509 0 1 1388
box 0 0 6 6
use CELL  95
transform 1 0 1011 0 1 1388
box 0 0 6 6
use CELL  96
transform -1 0 1064 0 -1 1098
box 0 0 6 6
use CELL  97
transform -1 0 1061 0 1 1388
box 0 0 6 6
use CELL  98
transform -1 0 1345 0 1 1936
box 0 0 6 6
use CELL  99
transform -1 0 1379 0 1 1936
box 0 0 6 6
use CELL  100
transform 1 0 1410 0 1 1535
box 0 0 6 6
use CELL  101
transform -1 0 1130 0 1 1388
box 0 0 6 6
use CELL  102
transform 1 0 1489 0 -1 1394
box 0 0 6 6
use CELL  103
transform -1 0 1033 0 1 713
box 0 0 6 6
use CELL  104
transform -1 0 1092 0 1 557
box 0 0 6 6
use CELL  105
transform 1 0 1104 0 -1 563
box 0 0 6 6
use CELL  106
transform 1 0 1041 0 -1 1942
box 0 0 6 6
use CELL  107
transform -1 0 1055 0 1 506
box 0 0 6 6
use CELL  108
transform -1 0 1047 0 1 2449
box 0 0 6 6
use CELL  109
transform 1 0 1065 0 -1 2053
box 0 0 6 6
use CELL  110
transform -1 0 1078 0 1 2128
box 0 0 6 6
use CELL  111
transform -1 0 1334 0 1 2128
box 0 0 6 6
use CELL  112
transform -1 0 1386 0 1 959
box 0 0 6 6
use CELL  113
transform -1 0 1368 0 1 1668
box 0 0 6 6
use CELL  114
transform 1 0 1332 0 1 2047
box 0 0 6 6
use CELL  115
transform -1 0 1230 0 1 1936
box 0 0 6 6
use CELL  116
transform -1 0 1312 0 1 713
box 0 0 6 6
use CELL  117
transform -1 0 1020 0 -1 2134
box 0 0 6 6
use CELL  118
transform 1 0 1215 0 1 2300
box 0 0 6 6
use CELL  119
transform -1 0 1029 0 1 1668
box 0 0 6 6
use CELL  120
transform -1 0 1027 0 1 2128
box 0 0 6 6
use CELL  121
transform -1 0 1033 0 1 506
box 0 0 6 6
use CELL  122
transform -1 0 1368 0 1 812
box 0 0 6 6
use CELL  123
transform -1 0 1463 0 1 1388
box 0 0 6 6
use CELL  124
transform -1 0 1309 0 1 1535
box 0 0 6 6
use CELL  125
transform -1 0 1107 0 1 2047
box 0 0 6 6
use CELL  126
transform 1 0 1163 0 -1 563
box 0 0 6 6
use CELL  127
transform -1 0 1053 0 1 1253
box 0 0 6 6
use CELL  128
transform 1 0 1228 0 1 2300
box 0 0 6 6
use CELL  129
transform -1 0 1044 0 1 620
box 0 0 6 6
use CELL  130
transform -1 0 1184 0 1 2363
box 0 0 6 6
use CELL  131
transform -1 0 1033 0 1 557
box 0 0 6 6
use CELL  132
transform -1 0 1228 0 1 2300
box 0 0 6 6
use CELL  133
transform -1 0 1231 0 1 2047
box 0 0 6 6
use CELL  134
transform -1 0 1471 0 1 959
box 0 0 6 6
use CELL  135
transform -1 0 1081 0 1 1253
box 0 0 6 6
use CELL  136
transform -1 0 1246 0 -1 2241
box 0 0 6 6
use CELL  137
transform -1 0 1234 0 1 2128
box 0 0 6 6
use CELL  138
transform -1 0 1088 0 1 2235
box 0 0 6 6
use CELL  139
transform -1 0 1091 0 1 2363
box 0 0 6 6
use CELL  140
transform 1 0 1061 0 1 959
box 0 0 6 6
use CELL  141
transform -1 0 1039 0 1 2363
box 0 0 6 6
use CELL  142
transform -1 0 1049 0 1 1821
box 0 0 6 6
use CELL  143
transform -1 0 1270 0 1 2235
box 0 0 6 6
use CELL  144
transform -1 0 1042 0 1 1821
box 0 0 6 6
use CELL  145
transform -1 0 1091 0 1 620
box 0 0 6 6
use CELL  146
transform -1 0 1202 0 1 2300
box 0 0 6 6
use CELL  147
transform -1 0 1062 0 1 1535
box 0 0 6 6
use CELL  148
transform -1 0 1002 0 1 2047
box 0 0 6 6
use CELL  149
transform -1 0 1209 0 1 2300
box 0 0 6 6
use CELL  150
transform -1 0 1451 0 1 1388
box 0 0 6 6
use CELL  151
transform -1 0 1075 0 1 812
box 0 0 6 6
use CELL  152
transform 1 0 1265 0 1 620
box 0 0 6 6
use CELL  153
transform -1 0 1296 0 1 812
box 0 0 6 6
use CELL  154
transform 1 0 1366 0 -1 1942
box 0 0 6 6
use CELL  155
transform -1 0 1248 0 1 713
box 0 0 6 6
use CELL  156
transform 1 0 1135 0 -1 512
box 0 0 6 6
use CELL  157
transform 1 0 1399 0 -1 818
box 0 0 6 6
use CELL  158
transform -1 0 1190 0 1 557
box 0 0 6 6
use CELL  159
transform -1 0 1063 0 1 2449
box 0 0 6 6
use CELL  160
transform -1 0 1038 0 1 2408
box 0 0 6 6
use CELL  161
transform -1 0 1021 0 1 2047
box 0 0 6 6
use CELL  162
transform -1 0 1035 0 1 959
box 0 0 6 6
use CELL  163
transform -1 0 1042 0 1 2235
box 0 0 6 6
use CELL  164
transform -1 0 1193 0 1 2363
box 0 0 6 6
use CELL  165
transform -1 0 1033 0 1 2235
box 0 0 6 6
use CELL  166
transform -1 0 1061 0 1 1668
box 0 0 6 6
use CELL  167
transform 1 0 1108 0 -1 1259
box 0 0 6 6
use CELL  168
transform 1 0 1464 0 1 1092
box 0 0 6 6
use CELL  169
transform -1 0 1327 0 1 1821
box 0 0 6 6
use CELL  170
transform -1 0 1241 0 -1 2306
box 0 0 6 6
use CELL  171
transform -1 0 1206 0 1 1092
box 0 0 6 6
use CELL  172
transform -1 0 1119 0 1 713
box 0 0 6 6
use CELL  173
transform -1 0 1034 0 1 812
box 0 0 6 6
use CELL  174
transform 1 0 1441 0 -1 1674
box 0 0 6 6
use CELL  175
transform -1 0 1123 0 1 1388
box 0 0 6 6
use CELL  176
transform -1 0 1381 0 1 1253
box 0 0 6 6
use CELL  177
transform -1 0 1028 0 1 1092
box 0 0 6 6
use CELL  178
transform -1 0 1263 0 1 1936
box 0 0 6 6
use CELL  179
transform -1 0 1020 0 1 812
box 0 0 6 6
use CELL  180
transform -1 0 1043 0 1 812
box 0 0 6 6
use CELL  181
transform -1 0 1105 0 1 1535
box 0 0 6 6
use CELL  182
transform 1 0 1284 0 -1 626
box 0 0 6 6
use CELL  183
transform 1 0 978 0 -1 965
box 0 0 6 6
use CELL  184
transform -1 0 1516 0 1 1388
box 0 0 6 6
use CELL  185
transform -1 0 1060 0 -1 965
box 0 0 6 6
use CELL  186
transform -1 0 1124 0 1 2408
box 0 0 6 6
use CELL  187
transform -1 0 1423 0 1 1535
box 0 0 6 6
use CELL  188
transform -1 0 1074 0 1 1253
box 0 0 6 6
use CELL  189
transform 1 0 1299 0 -1 719
box 0 0 6 6
use CELL  190
transform 1 0 1313 0 1 713
box 0 0 6 6
use CELL  191
transform 1 0 1022 0 1 1821
box 0 0 6 6
use CELL  192
transform -1 0 1117 0 1 557
box 0 0 6 6
use CELL  193
transform -1 0 1421 0 1 1388
box 0 0 6 6
use CELL  194
transform 1 0 992 0 1 959
box 0 0 6 6
use CELL  195
transform -1 0 1264 0 1 620
box 0 0 6 6
use CELL  196
transform -1 0 1093 0 1 1388
box 0 0 6 6
use CELL  197
transform -1 0 1228 0 1 1253
box 0 0 6 6
use CELL  198
transform -1 0 967 0 -1 965
box 0 0 6 6
use CELL  199
transform -1 0 1405 0 1 1821
box 0 0 6 6
use CELL  200
transform -1 0 1083 0 1 959
box 0 0 6 6
use CELL  201
transform -1 0 1359 0 1 1821
box 0 0 6 6
use CELL  202
transform -1 0 1305 0 -1 965
box 0 0 6 6
use CELL  203
transform -1 0 1095 0 1 713
box 0 0 6 6
use CELL  204
transform -1 0 1204 0 1 1535
box 0 0 6 6
use CELL  205
transform -1 0 1413 0 1 1668
box 0 0 6 6
use CELL  206
transform -1 0 1211 0 1 557
box 0 0 6 6
use CELL  207
transform -1 0 1079 0 1 1668
box 0 0 6 6
use CELL  208
transform -1 0 1419 0 1 812
box 0 0 6 6
use CELL  209
transform 1 0 1339 0 -1 1827
box 0 0 6 6
use CELL  210
transform -1 0 1014 0 1 1821
box 0 0 6 6
use CELL  211
transform -1 0 1245 0 1 1092
box 0 0 6 6
use CELL  212
transform -1 0 1444 0 1 1535
box 0 0 6 6
use CELL  213
transform -1 0 1021 0 1 1936
box 0 0 6 6
use CELL  214
transform 1 0 1320 0 1 1936
box 0 0 6 6
use CELL  215
transform -1 0 1028 0 -1 1541
box 0 0 6 6
use CELL  216
transform -1 0 1049 0 1 2235
box 0 0 6 6
use CELL  217
transform -1 0 1225 0 1 557
box 0 0 6 6
use CELL  218
transform -1 0 1056 0 1 2449
box 0 0 6 6
use CELL  219
transform -1 0 1214 0 1 620
box 0 0 6 6
use CELL  220
transform -1 0 1416 0 1 959
box 0 0 6 6
use CELL  221
transform 1 0 1327 0 1 713
box 0 0 6 6
use CELL  222
transform -1 0 1075 0 1 1936
box 0 0 6 6
use CELL  223
transform -1 0 1107 0 1 1668
box 0 0 6 6
use CELL  224
transform -1 0 1289 0 1 2235
box 0 0 6 6
use CELL  225
transform -1 0 1026 0 1 557
box 0 0 6 6
use CELL  226
transform -1 0 1082 0 -1 1942
box 0 0 6 6
use CELL  227
transform 1 0 1042 0 1 557
box 0 0 6 6
use CELL  228
transform -1 0 1081 0 1 2235
box 0 0 6 6
use CELL  229
transform -1 0 1213 0 1 1253
box 0 0 6 6
use CELL  230
transform -1 0 1287 0 1 713
box 0 0 6 6
use CELL  231
transform -1 0 1082 0 1 506
box 0 0 6 6
use CELL  232
transform -1 0 1184 0 1 2300
box 0 0 6 6
use CELL  233
transform -1 0 1024 0 1 1388
box 0 0 6 6
use CELL  234
transform 1 0 1224 0 -1 2241
box 0 0 6 6
use CELL  235
transform -1 0 1064 0 1 2047
box 0 0 6 6
use CELL  236
transform -1 0 1084 0 1 1821
box 0 0 6 6
use CELL  237
transform -1 0 1071 0 1 1092
box 0 0 6 6
use CELL  238
transform -1 0 1200 0 1 2363
box 0 0 6 6
use CELL  239
transform -1 0 1046 0 1 506
box 0 0 6 6
use CELL  240
transform 1 0 1177 0 -1 2134
box 0 0 6 6
use CELL  241
transform -1 0 1076 0 1 713
box 0 0 6 6
use CELL  242
transform -1 0 1057 0 1 812
box 0 0 6 6
use CELL  243
transform -1 0 1070 0 1 1821
box 0 0 6 6
use CELL  244
transform 1 0 1231 0 -1 563
box 0 0 6 6
use CELL  245
transform -1 0 1068 0 1 1388
box 0 0 6 6
use CELL  246
transform -1 0 1386 0 1 1821
box 0 0 6 6
use CELL  247
transform -1 0 1359 0 1 1936
box 0 0 6 6
use CELL  248
transform -1 0 1502 0 1 1388
box 0 0 6 6
use CELL  249
transform -1 0 1078 0 1 2300
box 0 0 6 6
use CELL  250
transform -1 0 1388 0 1 1253
box 0 0 6 6
use CELL  251
transform 1 0 1299 0 -1 1942
box 0 0 6 6
use CELL  252
transform 1 0 1008 0 1 1535
box 0 0 6 6
use CELL  253
transform -1 0 1226 0 1 620
box 0 0 6 6
use CELL  254
transform -1 0 1104 0 1 812
box 0 0 6 6
use CELL  255
transform -1 0 1014 0 1 2047
box 0 0 6 6
use CELL  256
transform 1 0 1217 0 -1 2241
box 0 0 6 6
use CELL  257
transform 1 0 1059 0 1 1253
box 0 0 6 6
use CELL  258
transform -1 0 1463 0 1 1092
box 0 0 6 6
use CELL  259
transform -1 0 1031 0 1 1388
box 0 0 6 6
use CELL  260
transform -1 0 1055 0 1 1535
box 0 0 6 6
use CELL  261
transform 1 0 985 0 -1 965
box 0 0 6 6
use CELL  262
transform -1 0 1054 0 1 1668
box 0 0 6 6
use CELL  263
transform -1 0 1402 0 1 1535
box 0 0 6 6
use CELL  264
transform -1 0 1319 0 1 1936
box 0 0 6 6
use CELL  265
transform -1 0 1341 0 1 2128
box 0 0 6 6
use CELL  266
transform -1 0 1076 0 1 959
box 0 0 6 6
use CELL  267
transform -1 0 1057 0 1 2047
box 0 0 6 6
use CELL  268
transform -1 0 1435 0 1 812
box 0 0 6 6
use CELL  269
transform -1 0 1052 0 1 2408
box 0 0 6 6
use CELL  270
transform -1 0 1089 0 1 1936
box 0 0 6 6
use CELL  271
transform -1 0 1240 0 1 1821
box 0 0 6 6
use CELL  272
transform -1 0 1154 0 1 2408
box 0 0 6 6
use CELL  273
transform 1 0 1427 0 -1 1674
box 0 0 6 6
use CELL  274
transform -1 0 1449 0 1 812
box 0 0 6 6
use CELL  275
transform -1 0 1032 0 1 2363
box 0 0 6 6
use CELL  276
transform 1 0 1441 0 1 1253
box 0 0 6 6
use CELL  277
transform 1 0 1448 0 1 1253
box 0 0 6 6
use CELL  278
transform -1 0 1046 0 1 1253
box 0 0 6 6
use CELL  279
transform -1 0 1247 0 -1 2306
box 0 0 6 6
use CELL  280
transform -1 0 1045 0 1 2128
box 0 0 6 6
use CELL  281
transform -1 0 1049 0 1 1092
box 0 0 6 6
use CELL  282
transform -1 0 1021 0 1 959
box 0 0 6 6
use CELL  283
transform -1 0 1050 0 1 2047
box 0 0 6 6
use CELL  284
transform -1 0 1488 0 1 1388
box 0 0 6 6
use CELL  285
transform -1 0 1098 0 1 506
box 0 0 6 6
use CELL  286
transform 1 0 1065 0 -1 2306
box 0 0 6 6
use CELL  287
transform 1 0 1273 0 1 2128
box 0 0 6 6
use CELL  288
transform -1 0 1148 0 1 2408
box 0 0 6 6
use CELL  289
transform -1 0 1352 0 -1 1942
box 0 0 6 6
use CELL  290
transform -1 0 1055 0 -1 563
box 0 0 6 6
use CELL  291
transform 1 0 1248 0 1 2300
box 0 0 6 6
use CELL  292
transform 1 0 1130 0 1 2408
box 0 0 6 6
use CELL  293
transform -1 0 1035 0 1 1092
box 0 0 6 6
use CELL  294
transform -1 0 1050 0 1 812
box 0 0 6 6
use CELL  295
transform 1 0 1424 0 -1 1541
box 0 0 6 6
use CELL  296
transform 1 0 1261 0 1 2047
box 0 0 6 6
use CELL  297
transform -1 0 1312 0 1 1936
box 0 0 6 6
use CELL  298
transform -1 0 1386 0 1 812
box 0 0 6 6
use CELL  299
transform -1 0 1395 0 1 1668
box 0 0 6 6
use CELL  300
transform 1 0 1079 0 1 2300
box 0 0 6 6
use CELL  301
transform -1 0 1100 0 -1 2414
box 0 0 6 6
use CELL  302
transform -1 0 1348 0 1 2128
box 0 0 6 6
use CELL  303
transform -1 0 1014 0 -1 1942
box 0 0 6 6
use CELL  304
transform 1 0 1092 0 -1 1541
box 0 0 6 6
use CELL  305
transform -1 0 1326 0 1 713
box 0 0 6 6
use CELL  306
transform -1 0 1269 0 1 1668
box 0 0 6 6
use CELL  307
transform -1 0 1322 0 1 2047
box 0 0 6 6
use CELL  308
transform 1 0 1079 0 1 557
box 0 0 6 6
use CELL  309
transform -1 0 1070 0 1 2363
box 0 0 6 6
use CELL  310
transform 1 0 1064 0 1 2449
box 0 0 6 6
use CELL  311
transform 1 0 1233 0 -1 2241
box 0 0 6 6
use CELL  312
transform -1 0 1248 0 1 1668
box 0 0 6 6
use CELL  313
transform -1 0 1028 0 1 2047
box 0 0 6 6
use CELL  314
transform -1 0 1046 0 1 2300
box 0 0 6 6
use CELL  315
transform -1 0 1405 0 1 1092
box 0 0 6 6
use CELL  316
transform -1 0 1477 0 1 1092
box 0 0 6 6
use CELL  317
transform -1 0 1427 0 1 1092
box 0 0 6 6
use CELL  318
transform -1 0 1128 0 1 1936
box 0 0 6 6
use CELL  319
transform -1 0 1059 0 1 620
box 0 0 6 6
use CELL  320
transform -1 0 1028 0 1 1936
box 0 0 6 6
use CELL  321
transform 1 0 1349 0 1 713
box 0 0 6 6
use CELL  322
transform -1 0 1022 0 1 1253
box 0 0 6 6
use CELL  323
transform -1 0 1008 0 1 1668
box 0 0 6 6
use CELL  324
transform -1 0 1032 0 1 2300
box 0 0 6 6
use CELL  325
transform -1 0 1442 0 -1 818
box 0 0 6 6
use CELL  326
transform -1 0 1350 0 1 959
box 0 0 6 6
use CELL  327
transform -1 0 1045 0 1 2408
box 0 0 6 6
use CELL  328
transform -1 0 1021 0 1 1092
box 0 0 6 6
use CELL  329
transform -1 0 1327 0 1 2128
box 0 0 6 6
use CELL  330
transform -1 0 1255 0 1 2128
box 0 0 6 6
use CELL  331
transform -1 0 1035 0 1 1821
box 0 0 6 6
use CELL  332
transform -1 0 1021 0 1 1535
box 0 0 6 6
use CELL  333
transform -1 0 1054 0 1 713
box 0 0 6 6
use CELL  334
transform -1 0 1040 0 1 1535
box 0 0 6 6
use CELL  335
transform 1 0 1251 0 1 620
box 0 0 6 6
use CELL  336
transform -1 0 1478 0 1 959
box 0 0 6 6
use CELL  337
transform -1 0 1028 0 1 959
box 0 0 6 6
use CELL  338
transform -1 0 1023 0 1 620
box 0 0 6 6
use CELL  339
transform -1 0 1441 0 1 959
box 0 0 6 6
use CELL  340
transform 1 0 1445 0 -1 1098
box 0 0 6 6
use CELL  341
transform -1 0 1067 0 1 2235
box 0 0 6 6
use CELL  342
transform -1 0 1366 0 1 1936
box 0 0 6 6
use CELL  343
transform -1 0 1262 0 1 1388
box 0 0 6 6
use CELL  344
transform 1 0 1349 0 1 2128
box 0 0 6 6
use CELL  345
transform -1 0 1312 0 1 2128
box 0 0 6 6
use CELL  346
transform -1 0 1014 0 1 959
box 0 0 6 6
use CELL  347
transform -1 0 1212 0 1 713
box 0 0 6 6
use CELL  348
transform -1 0 1082 0 1 812
box 0 0 6 6
use CELL  349
transform -1 0 1035 0 1 1936
box 0 0 6 6
use CELL  350
transform -1 0 1037 0 1 620
box 0 0 6 6
use CELL  351
transform -1 0 1434 0 1 959
box 0 0 6 6
use CELL  352
transform -1 0 1440 0 1 1253
box 0 0 6 6
use CELL  353
transform -1 0 1068 0 1 1936
box 0 0 6 6
use CELL  354
transform -1 0 1420 0 1 1668
box 0 0 6 6
use CELL  355
transform 1 0 1325 0 1 2047
box 0 0 6 6
use CELL  356
transform -1 0 1130 0 1 620
box 0 0 6 6
use CELL  357
transform -1 0 1040 0 1 506
box 0 0 6 6
use CELL  358
transform 1 0 1213 0 1 1821
box 0 0 6 6
use CELL  359
transform -1 0 1406 0 1 1253
box 0 0 6 6
use CELL  360
transform -1 0 1089 0 1 506
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 1103 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 1094 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 1097 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 1167 0 1 812
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 1278 0 1 959
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 1197 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 1192 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 1253 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 1469 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 1406 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 1189 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 1185 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 1174 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 1175 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 1086 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 1067 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 1332 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 1375 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 1439 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 1378 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 1442 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 1339 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 1079 0 1 713
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 1136 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 1172 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 1175 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 1291 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 1297 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 1294 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 1300 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 1246 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 1209 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 1263 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 1279 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 1306 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 1278 0 1 620
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 1225 0 1 557
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 1098 0 1 506
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 1181 0 1 557
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 1160 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 1121 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 1211 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 1163 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 1118 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 1121 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 1124 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 1398 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 1390 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 1463 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 1421 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 1451 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 1215 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 1210 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 1239 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 1374 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 1377 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 1362 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 1333 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 1264 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 1344 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 1354 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 1427 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 1388 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 1405 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 1398 0 1 959
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 1374 0 1 812
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 1272 0 1 713
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 1226 0 1 620
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 1248 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 1267 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 1251 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 1255 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 1255 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 1333 0 1 713
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 1426 0 1 812
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 1462 0 1 959
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 1033 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 1105 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 1033 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 1092 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 1143 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 1300 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 1403 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 1317 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 1362 0 1 959
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 1202 0 1 557
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 1241 0 1 620
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 1293 0 1 713
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 1386 0 1 812
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 1404 0 1 959
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 1408 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 1394 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 1433 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 1369 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 1214 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 1149 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 1042 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 1126 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 1077 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 1056 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 1202 0 1 620
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 1188 0 1 713
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 1245 0 1 812
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 1141 0 1 557
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 1205 0 1 620
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 1173 0 1 713
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 1206 0 1 812
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 1305 0 1 959
box 0 0 3 6
use FEEDTHRU  F-109
transform 1 0 1119 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-110
transform 1 0 1120 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-111
transform 1 0 1117 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-112
transform 1 0 1229 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-113
transform 1 0 1120 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-114
transform 1 0 1052 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-115
transform 1 0 1037 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-116
transform 1 0 1043 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-117
transform 1 0 1040 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-118
transform 1 0 1034 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-119
transform 1 0 1049 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-120
transform 1 0 1014 0 1 620
box 0 0 3 6
use FEEDTHRU  F-121
transform 1 0 1033 0 1 713
box 0 0 3 6
use FEEDTHRU  F-122
transform 1 0 1034 0 1 812
box 0 0 3 6
use FEEDTHRU  F-123
transform 1 0 1439 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-124
transform 1 0 1422 0 1 959
box 0 0 3 6
use FEEDTHRU  F-125
transform 1 0 1442 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-126
transform 1 0 1425 0 1 959
box 0 0 3 6
use FEEDTHRU  F-127
transform 1 0 1427 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-128
transform 1 0 1412 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-129
transform 1 0 1451 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-130
transform 1 0 1387 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-131
transform 1 0 1404 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-132
transform 1 0 1327 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-133
transform 1 0 1287 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-134
transform 1 0 1303 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-135
transform 1 0 1315 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-136
transform 1 0 1270 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-137
transform 1 0 1401 0 1 959
box 0 0 3 6
use FEEDTHRU  F-138
transform 1 0 1377 0 1 812
box 0 0 3 6
use FEEDTHRU  F-139
transform 1 0 1088 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-140
transform 1 0 1091 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-141
transform 1 0 1141 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-142
transform 1 0 1073 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-143
transform 1 0 1055 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-144
transform 1 0 1227 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-145
transform 1 0 1255 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-146
transform 1 0 1168 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-147
transform 1 0 1161 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-148
transform 1 0 1108 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-149
transform 1 0 1139 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-150
transform 1 0 1157 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-151
transform 1 0 1109 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-152
transform 1 0 1144 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-153
transform 1 0 1136 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-154
transform 1 0 1347 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-155
transform 1 0 1351 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-156
transform 1 0 1409 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-157
transform 1 0 1315 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-158
transform 1 0 1344 0 1 812
box 0 0 3 6
use FEEDTHRU  F-159
transform 1 0 1197 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-160
transform 1 0 1221 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-161
transform 1 0 1204 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-162
transform 1 0 1164 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-163
transform 1 0 1201 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-164
transform 1 0 1224 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-165
transform 1 0 1252 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-166
transform 1 0 1352 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-167
transform 1 0 1097 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-168
transform 1 0 1094 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-169
transform 1 0 1079 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-170
transform 1 0 1162 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-171
transform 1 0 1065 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-172
transform 1 0 1074 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-173
transform 1 0 1355 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-174
transform 1 0 1258 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-175
transform 1 0 1261 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-176
transform 1 0 1303 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-177
transform 1 0 1119 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-178
transform 1 0 1322 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-179
transform 1 0 1078 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-180
transform 1 0 1109 0 1 620
box 0 0 3 6
use FEEDTHRU  F-181
transform 1 0 1152 0 1 713
box 0 0 3 6
use FEEDTHRU  F-182
transform 1 0 1104 0 1 812
box 0 0 3 6
use FEEDTHRU  F-183
transform 1 0 1275 0 1 959
box 0 0 3 6
use FEEDTHRU  F-184
transform 1 0 1089 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-185
transform 1 0 1183 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-186
transform 1 0 1250 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-187
transform 1 0 1222 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-188
transform 1 0 1200 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-189
transform 1 0 1198 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-190
transform 1 0 1406 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-191
transform 1 0 1303 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-192
transform 1 0 1320 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-193
transform 1 0 1365 0 1 959
box 0 0 3 6
use FEEDTHRU  F-194
transform 1 0 1251 0 1 812
box 0 0 3 6
use FEEDTHRU  F-195
transform 1 0 1200 0 1 713
box 0 0 3 6
use FEEDTHRU  F-196
transform 1 0 1172 0 1 620
box 0 0 3 6
use FEEDTHRU  F-197
transform 1 0 1386 0 1 959
box 0 0 3 6
use FEEDTHRU  F-198
transform 1 0 1287 0 1 713
box 0 0 3 6
use FEEDTHRU  F-199
transform 1 0 1229 0 1 620
box 0 0 3 6
use FEEDTHRU  F-200
transform 1 0 1196 0 1 557
box 0 0 3 6
use FEEDTHRU  F-201
transform 1 0 1127 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-202
transform 1 0 1174 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-203
transform 1 0 1173 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-204
transform 1 0 1113 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-205
transform 1 0 1114 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-206
transform 1 0 1116 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-207
transform 1 0 1472 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-208
transform 1 0 1382 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-209
transform 1 0 1409 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-210
transform 1 0 1386 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-211
transform 1 0 1368 0 1 959
box 0 0 3 6
use FEEDTHRU  F-212
transform 1 0 1356 0 1 812
box 0 0 3 6
use FEEDTHRU  F-213
transform 1 0 1266 0 1 713
box 0 0 3 6
use FEEDTHRU  F-214
transform 1 0 1309 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-215
transform 1 0 1346 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-216
transform 1 0 1354 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-217
transform 1 0 1350 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-218
transform 1 0 1320 0 1 959
box 0 0 3 6
use FEEDTHRU  F-219
transform 1 0 1347 0 1 812
box 0 0 3 6
use FEEDTHRU  F-220
transform 1 0 1110 0 1 713
box 0 0 3 6
use FEEDTHRU  F-221
transform 1 0 1076 0 1 557
box 0 0 3 6
use FEEDTHRU  F-222
transform 1 0 1082 0 1 620
box 0 0 3 6
use FEEDTHRU  F-223
transform 1 0 1094 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-224
transform 1 0 1296 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-225
transform 1 0 1300 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-226
transform 1 0 1312 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-227
transform 1 0 1033 0 1 557
box 0 0 3 6
use FEEDTHRU  F-228
transform 1 0 1044 0 1 620
box 0 0 3 6
use FEEDTHRU  F-229
transform 1 0 1061 0 1 713
box 0 0 3 6
use FEEDTHRU  F-230
transform 1 0 1066 0 1 812
box 0 0 3 6
use FEEDTHRU  F-231
transform 1 0 1051 0 1 959
box 0 0 3 6
use FEEDTHRU  F-232
transform 1 0 1049 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-233
transform 1 0 1065 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-234
transform 1 0 1063 0 1 812
box 0 0 3 6
use FEEDTHRU  F-235
transform 1 0 1185 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-236
transform 1 0 1201 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-237
transform 1 0 1175 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-238
transform 1 0 1169 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-239
transform 1 0 1151 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-240
transform 1 0 1209 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-241
transform 1 0 1219 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-242
transform 1 0 1248 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-243
transform 1 0 1258 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-244
transform 1 0 1289 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-245
transform 1 0 1206 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-246
transform 1 0 1182 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-247
transform 1 0 1146 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-248
transform 1 0 1263 0 1 959
box 0 0 3 6
use FEEDTHRU  F-249
transform 1 0 1158 0 1 812
box 0 0 3 6
use FEEDTHRU  F-250
transform 1 0 1383 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-251
transform 1 0 1345 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-252
transform 1 0 1388 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-253
transform 1 0 1312 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-254
transform 1 0 1272 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-255
transform 1 0 1273 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-256
transform 1 0 1386 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-257
transform 1 0 1048 0 1 959
box 0 0 3 6
use FEEDTHRU  F-258
transform 1 0 1068 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-259
transform 1 0 1053 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-260
transform 1 0 1074 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-261
transform 1 0 1074 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-262
transform 1 0 1395 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-263
transform 1 0 1366 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-264
transform 1 0 1186 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-265
transform 1 0 1221 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-266
transform 1 0 1176 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-267
transform 1 0 1071 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-268
transform 1 0 1067 0 1 959
box 0 0 3 6
use FEEDTHRU  F-269
transform 1 0 1088 0 1 812
box 0 0 3 6
use FEEDTHRU  F-270
transform 1 0 1076 0 1 713
box 0 0 3 6
use FEEDTHRU  F-271
transform 1 0 1117 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-272
transform 1 0 1203 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-273
transform 1 0 1225 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-274
transform 1 0 1187 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-275
transform 1 0 1061 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-276
transform 1 0 1076 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-277
transform 1 0 1058 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-278
transform 1 0 1038 0 1 2449
box 0 0 3 6
use FEEDTHRU  F-279
transform 1 0 1091 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-280
transform 1 0 1397 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-281
transform 1 0 1411 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-282
transform 1 0 1357 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-283
transform 1 0 1374 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-284
transform 1 0 1356 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-285
transform 1 0 1407 0 1 959
box 0 0 3 6
use FEEDTHRU  F-286
transform 1 0 1389 0 1 812
box 0 0 3 6
use FEEDTHRU  F-287
transform 1 0 1088 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-288
transform 1 0 1085 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-289
transform 1 0 1070 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-290
transform 1 0 1128 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-291
transform 1 0 1155 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-292
transform 1 0 1150 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-293
transform 1 0 1167 0 1 713
box 0 0 3 6
use FEEDTHRU  F-294
transform 1 0 1197 0 1 812
box 0 0 3 6
use FEEDTHRU  F-295
transform 1 0 1203 0 1 959
box 0 0 3 6
use FEEDTHRU  F-296
transform 1 0 1155 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-297
transform 1 0 1140 0 1 713
box 0 0 3 6
use FEEDTHRU  F-298
transform 1 0 1128 0 1 812
box 0 0 3 6
use FEEDTHRU  F-299
transform 1 0 1200 0 1 959
box 0 0 3 6
use FEEDTHRU  F-300
transform 1 0 1140 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-301
transform 1 0 1121 0 1 620
box 0 0 3 6
use FEEDTHRU  F-302
transform 1 0 1097 0 1 620
box 0 0 3 6
use FEEDTHRU  F-303
transform 1 0 1146 0 1 713
box 0 0 3 6
use FEEDTHRU  F-304
transform 1 0 1134 0 1 812
box 0 0 3 6
use FEEDTHRU  F-305
transform 1 0 1318 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-306
transform 1 0 1306 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-307
transform 1 0 1285 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-308
transform 1 0 1330 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-309
transform 1 0 1389 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-310
transform 1 0 1371 0 1 959
box 0 0 3 6
use FEEDTHRU  F-311
transform 1 0 1359 0 1 812
box 0 0 3 6
use FEEDTHRU  F-312
transform 1 0 1269 0 1 713
box 0 0 3 6
use FEEDTHRU  F-313
transform 1 0 1214 0 1 620
box 0 0 3 6
use FEEDTHRU  F-314
transform 1 0 1324 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-315
transform 1 0 1297 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-316
transform 1 0 1062 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-317
transform 1 0 1079 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-318
transform 1 0 1061 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-319
transform 1 0 1059 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-320
transform 1 0 1034 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-321
transform 1 0 1454 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-322
transform 1 0 1080 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-323
transform 1 0 1191 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-324
transform 1 0 1164 0 1 959
box 0 0 3 6
use FEEDTHRU  F-325
transform 1 0 1157 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-326
transform 1 0 1102 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-327
transform 1 0 1333 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-328
transform 1 0 1359 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-329
transform 1 0 1189 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-330
transform 1 0 1158 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-331
transform 1 0 1212 0 1 959
box 0 0 3 6
use FEEDTHRU  F-332
transform 1 0 1164 0 1 812
box 0 0 3 6
use FEEDTHRU  F-333
transform 1 0 1238 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-334
transform 1 0 1225 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-335
transform 1 0 1466 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-336
transform 1 0 1393 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-337
transform 1 0 1401 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-338
transform 1 0 1300 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-339
transform 1 0 1095 0 1 713
box 0 0 3 6
use FEEDTHRU  F-340
transform 1 0 1101 0 1 557
box 0 0 3 6
use FEEDTHRU  F-341
transform 1 0 1103 0 1 620
box 0 0 3 6
use FEEDTHRU  F-342
transform 1 0 1098 0 1 557
box 0 0 3 6
use FEEDTHRU  F-343
transform 1 0 1083 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-344
transform 1 0 1073 0 1 506
box 0 0 3 6
use FEEDTHRU  F-345
transform 1 0 1061 0 1 506
box 0 0 3 6
use FEEDTHRU  F-346
transform 1 0 1070 0 1 506
box 0 0 3 6
use FEEDTHRU  F-347
transform 1 0 1047 0 1 2449
box 0 0 3 6
use FEEDTHRU  F-348
transform 1 0 1076 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-349
transform 1 0 1088 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-350
transform 1 0 1120 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-351
transform 1 0 1131 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-352
transform 1 0 1126 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-353
transform 1 0 1106 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-354
transform 1 0 1151 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-355
transform 1 0 1267 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-356
transform 1 0 1252 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-357
transform 1 0 1270 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-358
transform 1 0 1230 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-359
transform 1 0 1212 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-360
transform 1 0 1184 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-361
transform 1 0 1347 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-362
transform 1 0 1357 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-363
transform 1 0 1430 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-364
transform 1 0 1391 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-365
transform 1 0 1239 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-366
transform 1 0 1200 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-367
transform 1 0 1222 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-368
transform 1 0 1190 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-369
transform 1 0 1190 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-370
transform 1 0 1157 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-371
transform 1 0 1139 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-372
transform 1 0 1332 0 1 812
box 0 0 3 6
use FEEDTHRU  F-373
transform 1 0 1332 0 1 959
box 0 0 3 6
use FEEDTHRU  F-374
transform 1 0 1341 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-375
transform 1 0 1312 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-376
transform 1 0 1296 0 1 713
box 0 0 3 6
use FEEDTHRU  F-377
transform 1 0 1326 0 1 812
box 0 0 3 6
use FEEDTHRU  F-378
transform 1 0 1326 0 1 959
box 0 0 3 6
use FEEDTHRU  F-379
transform 1 0 1335 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-380
transform 1 0 1306 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-381
transform 1 0 1436 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-382
transform 1 0 1093 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-383
transform 1 0 1098 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-384
transform 1 0 1099 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-385
transform 1 0 1095 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-386
transform 1 0 1107 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-387
transform 1 0 1096 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-388
transform 1 0 1101 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-389
transform 1 0 1089 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-390
transform 1 0 1102 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-391
transform 1 0 1055 0 1 557
box 0 0 3 6
use FEEDTHRU  F-392
transform 1 0 1073 0 1 620
box 0 0 3 6
use FEEDTHRU  F-393
transform 1 0 1101 0 1 713
box 0 0 3 6
use FEEDTHRU  F-394
transform 1 0 1119 0 1 812
box 0 0 3 6
use FEEDTHRU  F-395
transform 1 0 1134 0 1 959
box 0 0 3 6
use FEEDTHRU  F-396
transform 1 0 1104 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-397
transform 1 0 1093 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-398
transform 1 0 1061 0 1 557
box 0 0 3 6
use FEEDTHRU  F-399
transform 1 0 1079 0 1 620
box 0 0 3 6
use FEEDTHRU  F-400
transform 1 0 1107 0 1 713
box 0 0 3 6
use FEEDTHRU  F-401
transform 1 0 1116 0 1 812
box 0 0 3 6
use FEEDTHRU  F-402
transform 1 0 1089 0 1 959
box 0 0 3 6
use FEEDTHRU  F-403
transform 1 0 1101 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-404
transform 1 0 1099 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-405
transform 1 0 1105 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-406
transform 1 0 1046 0 1 506
box 0 0 3 6
use FEEDTHRU  F-407
transform 1 0 1067 0 1 557
box 0 0 3 6
use FEEDTHRU  F-408
transform 1 0 1254 0 1 812
box 0 0 3 6
use FEEDTHRU  F-409
transform 1 0 1301 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-410
transform 1 0 1240 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-411
transform 1 0 1158 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-412
transform 1 0 1165 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-413
transform 1 0 1118 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-414
transform 1 0 1124 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-415
transform 1 0 1197 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-416
transform 1 0 1195 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-417
transform 1 0 1114 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-418
transform 1 0 1137 0 1 713
box 0 0 3 6
use FEEDTHRU  F-419
transform 1 0 1155 0 1 812
box 0 0 3 6
use FEEDTHRU  F-420
transform 1 0 1146 0 1 959
box 0 0 3 6
use FEEDTHRU  F-421
transform 1 0 1185 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-422
transform 1 0 1134 0 1 713
box 0 0 3 6
use FEEDTHRU  F-423
transform 1 0 1146 0 1 812
box 0 0 3 6
use FEEDTHRU  F-424
transform 1 0 1137 0 1 959
box 0 0 3 6
use FEEDTHRU  F-425
transform 1 0 1128 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-426
transform 1 0 1175 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-427
transform 1 0 1073 0 1 557
box 0 0 3 6
use FEEDTHRU  F-428
transform 1 0 1249 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-429
transform 1 0 1368 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-430
transform 1 0 1345 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-431
transform 1 0 1364 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-432
transform 1 0 1327 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-433
transform 1 0 1368 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-434
transform 1 0 1315 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-435
transform 1 0 1350 0 1 959
box 0 0 3 6
use FEEDTHRU  F-436
transform 1 0 1371 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-437
transform 1 0 1348 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-438
transform 1 0 1367 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-439
transform 1 0 1189 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-440
transform 1 0 1178 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-441
transform 1 0 1142 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-442
transform 1 0 1154 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-443
transform 1 0 1112 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-444
transform 1 0 1115 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-445
transform 1 0 1161 0 1 959
box 0 0 3 6
use FEEDTHRU  F-446
transform 1 0 1085 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-447
transform 1 0 1126 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-448
transform 1 0 1134 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-449
transform 1 0 1132 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-450
transform 1 0 1152 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-451
transform 1 0 1135 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-452
transform 1 0 1130 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-453
transform 1 0 1174 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-454
transform 1 0 1134 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-455
transform 1 0 1143 0 1 959
box 0 0 3 6
use FEEDTHRU  F-456
transform 1 0 1152 0 1 812
box 0 0 3 6
use FEEDTHRU  F-457
transform 1 0 1234 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-458
transform 1 0 1231 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-459
transform 1 0 1254 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-460
transform 1 0 1288 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-461
transform 1 0 1338 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-462
transform 1 0 1372 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-463
transform 1 0 1319 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-464
transform 1 0 1128 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-465
transform 1 0 1167 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-466
transform 1 0 1144 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-467
transform 1 0 1148 0 1 620
box 0 0 3 6
use FEEDTHRU  F-468
transform 1 0 1161 0 1 713
box 0 0 3 6
use FEEDTHRU  F-469
transform 1 0 1126 0 1 557
box 0 0 3 6
use FEEDTHRU  F-470
transform 1 0 1160 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-471
transform 1 0 1163 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-472
transform 1 0 1198 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-473
transform 1 0 1166 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-474
transform 1 0 1133 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-475
transform 1 0 1127 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-476
transform 1 0 1077 0 1 2449
box 0 0 3 6
use FEEDTHRU  F-477
transform 1 0 1170 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-478
transform 1 0 1153 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-479
transform 1 0 1173 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-480
transform 1 0 1147 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-481
transform 1 0 1136 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-482
transform 1 0 1193 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-483
transform 1 0 1169 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-484
transform 1 0 1204 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-485
transform 1 0 1283 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-486
transform 1 0 1261 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-487
transform 1 0 1299 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-488
transform 1 0 1323 0 1 959
box 0 0 3 6
use FEEDTHRU  F-489
transform 1 0 1246 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-490
transform 1 0 1284 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-491
transform 1 0 1281 0 1 959
box 0 0 3 6
use FEEDTHRU  F-492
transform 1 0 1176 0 1 812
box 0 0 3 6
use FEEDTHRU  F-493
transform 1 0 1188 0 1 812
box 0 0 3 6
use FEEDTHRU  F-494
transform 1 0 1194 0 1 812
box 0 0 3 6
use FEEDTHRU  F-495
transform 1 0 1167 0 1 959
box 0 0 3 6
use FEEDTHRU  F-496
transform 1 0 1152 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-497
transform 1 0 1227 0 1 812
box 0 0 3 6
use FEEDTHRU  F-498
transform 1 0 1197 0 1 713
box 0 0 3 6
use FEEDTHRU  F-499
transform 1 0 1233 0 1 812
box 0 0 3 6
use FEEDTHRU  F-500
transform 1 0 1257 0 1 959
box 0 0 3 6
use FEEDTHRU  F-501
transform 1 0 1263 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-502
transform 1 0 1266 0 1 812
box 0 0 3 6
use FEEDTHRU  F-503
transform 1 0 1193 0 1 620
box 0 0 3 6
use FEEDTHRU  F-504
transform 1 0 1153 0 1 557
box 0 0 3 6
use FEEDTHRU  F-505
transform 1 0 1320 0 1 812
box 0 0 3 6
use FEEDTHRU  F-506
transform 1 0 1112 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-507
transform 1 0 1103 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-508
transform 1 0 1154 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-509
transform 1 0 1130 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-510
transform 1 0 1082 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-511
transform 1 0 1095 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-512
transform 1 0 1116 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-513
transform 1 0 1117 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-514
transform 1 0 1197 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-515
transform 1 0 1168 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-516
transform 1 0 1145 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-517
transform 1 0 1105 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-518
transform 1 0 1119 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-519
transform 1 0 1122 0 1 959
box 0 0 3 6
use FEEDTHRU  F-520
transform 1 0 1185 0 1 812
box 0 0 3 6
use FEEDTHRU  F-521
transform 1 0 1125 0 1 713
box 0 0 3 6
use FEEDTHRU  F-522
transform 1 0 1132 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-523
transform 1 0 1119 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-524
transform 1 0 1146 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-525
transform 1 0 1141 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-526
transform 1 0 1158 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-527
transform 1 0 1138 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-528
transform 1 0 1125 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-529
transform 1 0 1152 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-530
transform 1 0 1147 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-531
transform 1 0 1164 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-532
transform 1 0 1141 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-533
transform 1 0 1159 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-534
transform 1 0 1153 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-535
transform 1 0 1148 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-536
transform 1 0 1129 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-537
transform 1 0 1194 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-538
transform 1 0 1309 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-539
transform 1 0 1311 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-540
transform 1 0 1261 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-541
transform 1 0 1314 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-542
transform 1 0 1212 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-543
transform 1 0 1154 0 1 620
box 0 0 3 6
use FEEDTHRU  F-544
transform 1 0 1144 0 1 557
box 0 0 3 6
use FEEDTHRU  F-545
transform 1 0 1185 0 1 713
box 0 0 3 6
use FEEDTHRU  F-546
transform 1 0 1242 0 1 812
box 0 0 3 6
use FEEDTHRU  F-547
transform 1 0 1308 0 1 959
box 0 0 3 6
use FEEDTHRU  F-548
transform 1 0 1131 0 1 959
box 0 0 3 6
use FEEDTHRU  F-549
transform 1 0 1226 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-550
transform 1 0 1257 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-551
transform 1 0 1224 0 1 959
box 0 0 3 6
use FEEDTHRU  F-552
transform 1 0 1248 0 1 812
box 0 0 3 6
use FEEDTHRU  F-553
transform 1 0 1191 0 1 713
box 0 0 3 6
use FEEDTHRU  F-554
transform 1 0 1258 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-555
transform 1 0 1258 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-556
transform 1 0 1212 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-557
transform 1 0 1182 0 1 812
box 0 0 3 6
use FEEDTHRU  F-558
transform 1 0 1107 0 1 959
box 0 0 3 6
use FEEDTHRU  F-559
transform 1 0 1275 0 1 713
box 0 0 3 6
use FEEDTHRU  F-560
transform 1 0 1338 0 1 812
box 0 0 3 6
use FEEDTHRU  F-561
transform 1 0 1353 0 1 959
box 0 0 3 6
use FEEDTHRU  F-562
transform 1 0 1331 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-563
transform 1 0 1318 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-564
transform 1 0 1329 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-565
transform 1 0 1326 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-566
transform 1 0 1307 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-567
transform 1 0 1424 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-568
transform 1 0 1190 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-569
transform 1 0 1180 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-570
transform 1 0 1164 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-571
transform 1 0 1155 0 1 959
box 0 0 3 6
use FEEDTHRU  F-572
transform 1 0 1218 0 1 713
box 0 0 3 6
use FEEDTHRU  F-573
transform 1 0 1278 0 1 812
box 0 0 3 6
use FEEDTHRU  F-574
transform 1 0 1251 0 1 959
box 0 0 3 6
use FEEDTHRU  F-575
transform 1 0 1140 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-576
transform 1 0 1151 0 1 620
box 0 0 3 6
use FEEDTHRU  F-577
transform 1 0 1123 0 1 557
box 0 0 3 6
use FEEDTHRU  F-578
transform 1 0 1130 0 1 620
box 0 0 3 6
use FEEDTHRU  F-579
transform 1 0 1244 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-580
transform 1 0 1228 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-581
transform 1 0 1245 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-582
transform 1 0 1206 0 1 959
box 0 0 3 6
use FEEDTHRU  F-583
transform 1 0 1193 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-584
transform 1 0 1147 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-585
transform 1 0 1170 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-586
transform 1 0 1159 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-587
transform 1 0 1219 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-588
transform 1 0 1218 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-589
transform 1 0 1336 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-590
transform 1 0 1380 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-591
transform 1 0 1351 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-592
transform 1 0 1343 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-593
transform 1 0 1336 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-594
transform 1 0 1353 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-595
transform 1 0 1317 0 1 959
box 0 0 3 6
use FEEDTHRU  F-596
transform 1 0 1220 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-597
transform 1 0 1201 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-598
transform 1 0 1341 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-599
transform 1 0 1217 0 1 620
box 0 0 3 6
use FEEDTHRU  F-600
transform 1 0 1212 0 1 713
box 0 0 3 6
use FEEDTHRU  F-601
transform 1 0 1177 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-602
transform 1 0 1194 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-603
transform 1 0 1152 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-604
transform 1 0 1159 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-605
transform 1 0 1188 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-606
transform 1 0 1291 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-607
transform 1 0 1287 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-608
transform 1 0 1138 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-609
transform 1 0 1146 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-610
transform 1 0 1123 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-611
transform 1 0 1182 0 1 959
box 0 0 3 6
use FEEDTHRU  F-612
transform 1 0 1295 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-613
transform 1 0 1288 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-614
transform 1 0 1311 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-615
transform 1 0 1269 0 1 959
box 0 0 3 6
use FEEDTHRU  F-616
transform 1 0 1156 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-617
transform 1 0 1149 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-618
transform 1 0 1170 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-619
transform 1 0 1171 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-620
transform 1 0 1182 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-621
transform 1 0 1159 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-622
transform 1 0 1160 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-623
transform 1 0 1153 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-624
transform 1 0 1232 0 1 620
box 0 0 3 6
use FEEDTHRU  F-625
transform 1 0 1290 0 1 713
box 0 0 3 6
use FEEDTHRU  F-626
transform 1 0 1302 0 1 812
box 0 0 3 6
use FEEDTHRU  F-627
transform 1 0 1389 0 1 959
box 0 0 3 6
use FEEDTHRU  F-628
transform 1 0 1454 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-629
transform 1 0 1255 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-630
transform 1 0 1262 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-631
transform 1 0 1285 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-632
transform 1 0 1293 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-633
transform 1 0 1303 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-634
transform 1 0 1199 0 1 557
box 0 0 3 6
use FEEDTHRU  F-635
transform 1 0 1181 0 1 620
box 0 0 3 6
use FEEDTHRU  F-636
transform 1 0 1230 0 1 713
box 0 0 3 6
use FEEDTHRU  F-637
transform 1 0 1305 0 1 812
box 0 0 3 6
use FEEDTHRU  F-638
transform 1 0 1272 0 1 812
box 0 0 3 6
use FEEDTHRU  F-639
transform 1 0 1164 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-640
transform 1 0 1171 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-641
transform 1 0 1124 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-642
transform 1 0 1148 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-643
transform 1 0 1170 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-644
transform 1 0 1230 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-645
transform 1 0 1216 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-646
transform 1 0 1223 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-647
transform 1 0 1273 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-648
transform 1 0 1243 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-649
transform 1 0 1246 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-650
transform 1 0 1290 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-651
transform 1 0 1330 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-652
transform 1 0 1199 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-653
transform 1 0 1237 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-654
transform 1 0 1172 0 1 2300
box 0 0 3 6
use FEEDTHRU  F-655
transform 1 0 1148 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-656
transform 1 0 1195 0 1 2128
box 0 0 3 6
use FEEDTHRU  F-657
transform 1 0 1194 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-658
transform 1 0 1218 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-659
transform 1 0 1115 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-660
transform 1 0 1151 0 1 2235
box 0 0 3 6
use FEEDTHRU  F-661
transform 1 0 1191 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-662
transform 1 0 1183 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-663
transform 1 0 1206 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-664
transform 1 0 1195 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-665
transform 1 0 1178 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-666
transform 1 0 1165 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-667
transform 1 0 1176 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-668
transform 1 0 1236 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-669
transform 1 0 1219 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-670
transform 1 0 1202 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-671
transform 1 0 1204 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-672
transform 1 0 1215 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-673
transform 1 0 1173 0 1 959
box 0 0 3 6
use FEEDTHRU  F-674
transform 1 0 1239 0 1 812
box 0 0 3 6
use FEEDTHRU  F-675
transform 1 0 1067 0 1 506
box 0 0 3 6
use FEEDTHRU  F-676
transform 1 0 1164 0 1 713
box 0 0 3 6
use FEEDTHRU  F-677
transform 1 0 1112 0 1 620
box 0 0 3 6
use FEEDTHRU  F-678
transform 1 0 1118 0 1 620
box 0 0 3 6
use FEEDTHRU  F-679
transform 1 0 1224 0 1 812
box 0 0 3 6
use FEEDTHRU  F-680
transform 1 0 1149 0 1 959
box 0 0 3 6
use FEEDTHRU  F-681
transform 1 0 1188 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-682
transform 1 0 1177 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-683
transform 1 0 1184 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-684
transform 1 0 1192 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-685
transform 1 0 1218 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-686
transform 1 0 1228 0 1 557
box 0 0 3 6
use FEEDTHRU  F-687
transform 1 0 1281 0 1 620
box 0 0 3 6
use FEEDTHRU  F-688
transform 1 0 1278 0 1 713
box 0 0 3 6
use FEEDTHRU  F-689
transform 1 0 1341 0 1 812
box 0 0 3 6
use FEEDTHRU  F-690
transform 1 0 1242 0 1 959
box 0 0 3 6
use FEEDTHRU  F-691
transform 1 0 1293 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-692
transform 1 0 1267 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-693
transform 1 0 1268 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-694
transform 1 0 1330 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-695
transform 1 0 1371 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-696
transform 1 0 1318 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-697
transform 1 0 1293 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-698
transform 1 0 1348 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-699
transform 1 0 1264 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-700
transform 1 0 1299 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-701
transform 1 0 1252 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-702
transform 1 0 1275 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-703
transform 1 0 1203 0 1 713
box 0 0 3 6
use FEEDTHRU  F-704
transform 1 0 1260 0 1 812
box 0 0 3 6
use FEEDTHRU  F-705
transform 1 0 1188 0 1 959
box 0 0 3 6
use FEEDTHRU  F-706
transform 1 0 1227 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-707
transform 1 0 1218 0 1 959
box 0 0 3 6
use FEEDTHRU  F-708
transform 1 0 1284 0 1 812
box 0 0 3 6
use FEEDTHRU  F-709
transform 1 0 1224 0 1 713
box 0 0 3 6
use FEEDTHRU  F-710
transform 1 0 1175 0 1 620
box 0 0 3 6
use FEEDTHRU  F-711
transform 1 0 1169 0 1 557
box 0 0 3 6
use FEEDTHRU  F-712
transform 1 0 1276 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-713
transform 1 0 1100 0 1 2408
box 0 0 3 6
use FEEDTHRU  F-714
transform 1 0 1091 0 1 2363
box 0 0 3 6
use FEEDTHRU  F-715
transform 1 0 1212 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-716
transform 1 0 1207 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-717
transform 1 0 1236 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-718
transform 1 0 1228 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-719
transform 1 0 1335 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-720
transform 1 0 1234 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-721
transform 1 0 1248 0 1 959
box 0 0 3 6
use FEEDTHRU  F-722
transform 1 0 1290 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-723
transform 1 0 1273 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-724
transform 1 0 1280 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-725
transform 1 0 1282 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-726
transform 1 0 1317 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-727
transform 1 0 1282 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-728
transform 1 0 1336 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-729
transform 1 0 1154 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-730
transform 1 0 1171 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-731
transform 1 0 1203 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-732
transform 1 0 1155 0 1 2047
box 0 0 3 6
use FEEDTHRU  F-733
transform 1 0 1188 0 1 1936
box 0 0 3 6
use FEEDTHRU  F-734
transform 1 0 1182 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-735
transform 1 0 1171 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-736
transform 1 0 1172 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-737
transform 1 0 1186 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-738
transform 1 0 1119 0 1 959
box 0 0 3 6
use FEEDTHRU  F-739
transform 1 0 1234 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-740
transform 1 0 1251 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-741
transform 1 0 1269 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-742
transform 1 0 1221 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-743
transform 1 0 1213 0 1 1253
box 0 0 3 6
use FEEDTHRU  F-744
transform 1 0 1214 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-745
transform 1 0 1228 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-746
transform 1 0 1251 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-747
transform 1 0 1231 0 1 1821
box 0 0 3 6
use FEEDTHRU  F-748
transform 1 0 1233 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-749
transform 1 0 1194 0 1 959
box 0 0 3 6
use FEEDTHRU  F-750
transform 1 0 1170 0 1 713
box 0 0 3 6
use FEEDTHRU  F-751
transform 1 0 1142 0 1 1388
box 0 0 3 6
use FEEDTHRU  F-752
transform 1 0 1165 0 1 1535
box 0 0 3 6
use FEEDTHRU  F-753
transform 1 0 1194 0 1 1668
box 0 0 3 6
use FEEDTHRU  F-754
transform 1 0 1136 0 1 620
box 0 0 3 6
use FEEDTHRU  F-755
transform 1 0 1129 0 1 557
box 0 0 3 6
use FEEDTHRU  F-756
transform 1 0 1089 0 1 506
box 0 0 3 6
<< metal1 >>
rect 1028 497 1048 498
rect 1038 499 1069 500
rect 1041 501 1063 502
rect 1050 503 1072 504
rect 1074 503 1078 504
rect 1084 503 1091 504
rect 1099 503 1103 504
rect 1132 503 1140 504
rect 1021 513 1035 514
rect 1031 515 1057 516
rect 1044 517 1069 518
rect 1047 519 1069 520
rect 1046 521 1072 522
rect 1050 523 1063 524
rect 1028 525 1063 526
rect 1053 527 1075 528
rect 1028 529 1075 530
rect 1031 531 1054 532
rect 1077 531 1158 532
rect 1021 533 1078 534
rect 1080 533 1128 534
rect 1087 535 1171 536
rect 1090 537 1131 538
rect 1090 539 1103 540
rect 1093 541 1155 542
rect 1099 543 1183 544
rect 1087 545 1100 546
rect 1105 545 1227 546
rect 1112 547 1125 548
rect 1115 549 1146 550
rect 1142 551 1152 552
rect 1164 551 1198 552
rect 1167 553 1189 554
rect 1200 553 1221 554
rect 1203 555 1217 556
rect 1229 555 1236 556
rect 1009 564 1016 565
rect 1024 564 1029 565
rect 1028 566 1078 567
rect 1032 568 1100 569
rect 1034 570 1046 571
rect 1039 572 1069 573
rect 1043 574 1075 575
rect 1042 576 1216 577
rect 1056 578 1075 579
rect 1057 580 1114 581
rect 1062 582 1081 583
rect 1061 584 1099 585
rect 1064 586 1123 587
rect 1071 588 1111 589
rect 1083 590 1120 591
rect 1025 592 1084 593
rect 1086 592 1128 593
rect 1102 594 1105 595
rect 1115 594 1153 595
rect 1130 596 1138 597
rect 1124 598 1132 599
rect 1154 598 1195 599
rect 1145 600 1156 601
rect 1170 600 1177 601
rect 1173 602 1210 603
rect 1182 604 1186 605
rect 1182 606 1201 607
rect 1203 606 1243 607
rect 1148 608 1204 609
rect 1089 610 1150 611
rect 1206 610 1219 611
rect 1142 612 1207 613
rect 1223 612 1234 613
rect 1226 614 1280 615
rect 1220 616 1228 617
rect 1229 616 1283 617
rect 1197 618 1231 619
rect 1021 627 1097 628
rect 1035 629 1084 630
rect 1015 631 1035 632
rect 1039 631 1136 632
rect 1049 633 1123 634
rect 1052 635 1078 636
rect 1054 637 1172 638
rect 1057 639 1084 640
rect 1061 641 1142 642
rect 1045 643 1063 644
rect 1064 643 1169 644
rect 1071 645 1120 646
rect 1074 647 1103 648
rect 1080 649 1109 650
rect 1040 651 1081 652
rect 1089 651 1268 652
rect 1090 653 1105 654
rect 1098 655 1148 656
rect 1113 657 1166 658
rect 1114 659 1187 660
rect 1117 661 1156 662
rect 1125 663 1153 664
rect 1110 665 1154 666
rect 1025 667 1112 668
rect 1024 669 1038 670
rect 1126 669 1225 670
rect 1128 671 1138 672
rect 1042 673 1139 674
rect 1149 673 1163 674
rect 1173 673 1202 674
rect 1174 675 1207 676
rect 1176 677 1226 678
rect 1189 679 1204 680
rect 1192 681 1213 682
rect 1194 683 1247 684
rect 1204 685 1222 686
rect 1207 687 1210 688
rect 1131 689 1211 690
rect 1213 689 1219 690
rect 1215 691 1271 692
rect 1219 693 1301 694
rect 1227 695 1274 696
rect 1233 697 1292 698
rect 1242 699 1295 700
rect 1259 701 1286 702
rect 1276 703 1289 704
rect 1230 705 1289 706
rect 1182 707 1232 708
rect 1279 707 1338 708
rect 1279 709 1283 710
rect 1198 711 1283 712
rect 1297 711 1308 712
rect 1334 711 1345 712
rect 1015 720 1184 721
rect 1018 722 1112 723
rect 1021 724 1065 725
rect 1031 726 1097 727
rect 1028 728 1033 729
rect 1049 728 1172 729
rect 1048 730 1178 731
rect 1059 732 1081 733
rect 1062 734 1068 735
rect 1071 734 1166 735
rect 1070 736 1196 737
rect 1074 738 1160 739
rect 1090 740 1166 741
rect 1077 742 1090 743
rect 1102 742 1121 743
rect 1105 744 1154 745
rect 1041 746 1154 747
rect 1108 748 1118 749
rect 1114 750 1163 751
rect 1129 752 1142 753
rect 1138 754 1157 755
rect 1186 754 1244 755
rect 1126 756 1187 757
rect 1192 756 1250 757
rect 1198 758 1229 759
rect 1168 760 1199 761
rect 1083 762 1169 763
rect 1201 762 1253 763
rect 1204 764 1262 765
rect 1213 766 1286 767
rect 1225 768 1286 769
rect 1052 770 1226 771
rect 1240 770 1434 771
rect 1255 772 1367 773
rect 1267 774 1358 775
rect 1246 776 1268 777
rect 1189 778 1247 779
rect 1073 780 1190 781
rect 1270 780 1361 781
rect 1273 782 1376 783
rect 1207 784 1274 785
rect 1174 786 1208 787
rect 1276 786 1340 787
rect 1279 788 1343 789
rect 1219 790 1280 791
rect 1288 790 1411 791
rect 1294 792 1388 793
rect 1297 794 1328 795
rect 1303 796 1322 797
rect 1291 798 1304 799
rect 1234 800 1292 801
rect 1307 800 1391 801
rect 1231 802 1307 803
rect 1324 802 1349 803
rect 1334 804 1428 805
rect 1310 806 1334 807
rect 1344 806 1351 807
rect 1345 808 1408 809
rect 1378 810 1385 811
rect 955 819 963 820
rect 993 819 1036 820
rect 1012 821 1027 822
rect 1016 823 1065 824
rect 1029 825 1133 826
rect 1019 827 1031 828
rect 1038 827 1053 828
rect 1033 829 1038 830
rect 1052 829 1068 830
rect 1055 831 1307 832
rect 1058 833 1136 834
rect 1065 835 1163 836
rect 1068 837 1090 838
rect 1070 839 1178 840
rect 1071 841 1394 842
rect 1077 843 1190 844
rect 1078 845 1325 846
rect 1080 847 1096 848
rect 1090 849 1118 850
rect 1105 851 1277 852
rect 1108 853 1184 854
rect 1120 855 1136 856
rect 1009 857 1121 858
rect 1123 857 1187 858
rect 1129 859 1202 860
rect 1138 861 1148 862
rect 1144 863 1154 864
rect 1147 865 1157 866
rect 1074 867 1157 868
rect 1150 869 1226 870
rect 1159 871 1265 872
rect 1165 873 1214 874
rect 1048 875 1166 876
rect 1022 877 1050 878
rect 1174 877 1241 878
rect 1183 879 1382 880
rect 1189 881 1262 882
rect 1198 883 1205 884
rect 1207 883 1307 884
rect 1219 885 1286 886
rect 1225 887 1250 888
rect 1228 889 1295 890
rect 1234 891 1259 892
rect 1243 893 1310 894
rect 1243 895 1343 896
rect 1246 897 1364 898
rect 1249 899 1448 900
rect 1252 901 1367 902
rect 1252 903 1280 904
rect 1168 905 1280 906
rect 1168 907 1196 908
rect 1195 909 1440 910
rect 1255 911 1385 912
rect 1267 913 1415 914
rect 1270 915 1474 916
rect 1282 917 1301 918
rect 1318 917 1418 918
rect 1321 919 1401 920
rect 1321 921 1349 922
rect 1207 923 1349 924
rect 1339 925 1355 926
rect 1351 927 1470 928
rect 1357 929 1370 930
rect 1360 931 1373 932
rect 1363 933 1385 934
rect 1375 935 1400 936
rect 1378 937 1403 938
rect 1387 939 1406 940
rect 1387 941 1411 942
rect 1273 943 1412 944
rect 1390 945 1409 946
rect 1303 947 1391 948
rect 1396 947 1433 948
rect 1345 949 1397 950
rect 1102 951 1346 952
rect 1423 951 1461 952
rect 1427 953 1464 954
rect 1426 955 1458 956
rect 1437 957 1445 958
rect 979 966 987 967
rect 989 966 994 967
rect 1012 966 1109 967
rect 1019 968 1121 969
rect 1023 970 1050 971
rect 1026 972 1133 973
rect 1030 974 1056 975
rect 1030 976 1163 977
rect 1033 978 1172 979
rect 1050 980 1053 981
rect 1068 980 1073 981
rect 1074 980 1310 981
rect 1037 982 1076 983
rect 1037 984 1079 985
rect 1090 984 1103 985
rect 1090 986 1277 987
rect 1105 988 1136 989
rect 1120 990 1124 991
rect 1129 990 1139 991
rect 1135 992 1145 993
rect 1141 994 1202 995
rect 1147 996 1187 997
rect 1147 998 1265 999
rect 1153 1000 1169 1001
rect 1159 1002 1214 1003
rect 1066 1004 1214 1005
rect 1165 1006 1193 1007
rect 1156 1008 1166 1009
rect 1156 1010 1205 1011
rect 1174 1012 1217 1013
rect 1177 1014 1437 1015
rect 1183 1016 1241 1017
rect 1047 1018 1184 1019
rect 1189 1018 1229 1019
rect 1150 1020 1190 1021
rect 1195 1020 1235 1021
rect 1195 1022 1202 1023
rect 1198 1024 1280 1025
rect 1207 1026 1247 1027
rect 1243 1028 1295 1029
rect 1249 1030 1292 1031
rect 1258 1032 1265 1033
rect 1225 1034 1259 1035
rect 1270 1034 1313 1035
rect 1276 1036 1459 1037
rect 1282 1038 1286 1039
rect 1300 1038 1325 1039
rect 1306 1040 1385 1041
rect 1327 1042 1337 1043
rect 1333 1044 1343 1045
rect 1348 1044 1397 1045
rect 1354 1046 1477 1047
rect 1318 1048 1355 1049
rect 1318 1050 1364 1051
rect 1357 1052 1409 1053
rect 1375 1054 1415 1055
rect 1387 1056 1450 1057
rect 1369 1058 1388 1059
rect 1369 1060 1470 1061
rect 1390 1062 1456 1063
rect 1372 1064 1391 1065
rect 1351 1066 1373 1067
rect 1321 1068 1352 1069
rect 1321 1070 1367 1071
rect 1402 1070 1419 1071
rect 1222 1072 1404 1073
rect 1405 1072 1410 1073
rect 1399 1074 1407 1075
rect 1330 1076 1401 1077
rect 1412 1076 1433 1077
rect 1423 1078 1444 1079
rect 1252 1080 1423 1081
rect 1252 1082 1476 1083
rect 1426 1084 1429 1085
rect 1440 1084 1461 1085
rect 1219 1086 1462 1087
rect 1081 1088 1220 1089
rect 1452 1088 1467 1089
rect 1463 1090 1466 1091
rect 1006 1099 1036 1100
rect 1012 1101 1058 1102
rect 1013 1103 1055 1104
rect 1033 1105 1157 1106
rect 1037 1107 1119 1108
rect 1040 1109 1073 1110
rect 1041 1111 1061 1112
rect 1047 1113 1076 1114
rect 1048 1115 1116 1116
rect 1050 1117 1067 1118
rect 1062 1119 1193 1120
rect 1069 1121 1142 1122
rect 1038 1123 1070 1124
rect 1076 1123 1244 1124
rect 1078 1125 1384 1126
rect 1081 1127 1148 1128
rect 1094 1129 1106 1130
rect 1100 1131 1103 1132
rect 1019 1133 1104 1134
rect 1020 1135 1265 1136
rect 1106 1137 1121 1138
rect 1026 1139 1122 1140
rect 1109 1141 1196 1142
rect 1129 1143 1205 1144
rect 1135 1145 1176 1146
rect 1148 1147 1172 1148
rect 1153 1149 1227 1150
rect 1154 1151 1423 1152
rect 1165 1153 1182 1154
rect 1166 1155 1178 1156
rect 1172 1157 1184 1158
rect 1090 1159 1185 1160
rect 1178 1161 1190 1162
rect 1159 1163 1191 1164
rect 1063 1165 1161 1166
rect 1186 1165 1212 1166
rect 1193 1167 1199 1168
rect 1201 1167 1214 1168
rect 1044 1169 1203 1170
rect 1044 1171 1131 1172
rect 1205 1171 1217 1172
rect 1214 1173 1223 1174
rect 1228 1175 1401 1176
rect 1229 1177 1247 1178
rect 1234 1179 1426 1180
rect 1235 1181 1253 1182
rect 1247 1183 1286 1184
rect 1253 1185 1277 1186
rect 1256 1187 1456 1188
rect 1262 1189 1301 1190
rect 1268 1191 1295 1192
rect 1274 1193 1292 1194
rect 1289 1195 1313 1196
rect 1301 1197 1397 1198
rect 1304 1199 1322 1200
rect 1307 1201 1337 1202
rect 1313 1203 1343 1204
rect 1318 1205 1394 1206
rect 1319 1207 1331 1208
rect 1325 1209 1417 1210
rect 1331 1211 1391 1212
rect 1337 1213 1355 1214
rect 1346 1215 1370 1216
rect 1351 1217 1356 1218
rect 1348 1219 1353 1220
rect 1349 1221 1373 1222
rect 1357 1223 1432 1224
rect 1358 1225 1376 1226
rect 1258 1227 1377 1228
rect 1389 1227 1407 1228
rect 1392 1229 1447 1230
rect 1395 1231 1410 1232
rect 1387 1233 1411 1234
rect 1386 1235 1444 1236
rect 1398 1237 1413 1238
rect 1401 1239 1419 1240
rect 1404 1241 1426 1242
rect 1407 1243 1476 1244
rect 1413 1245 1429 1246
rect 1422 1247 1453 1248
rect 1438 1249 1466 1250
rect 1440 1251 1473 1252
rect 994 1260 999 1261
rect 1006 1260 1052 1261
rect 1013 1262 1030 1263
rect 1020 1264 1144 1265
rect 1008 1266 1020 1267
rect 1022 1266 1159 1267
rect 1026 1268 1119 1269
rect 1035 1270 1051 1271
rect 1066 1270 1212 1271
rect 1069 1272 1182 1273
rect 1010 1274 1070 1275
rect 1076 1274 1209 1275
rect 1054 1276 1076 1277
rect 1038 1278 1054 1279
rect 1091 1278 1161 1279
rect 1094 1280 1261 1281
rect 1106 1282 1147 1283
rect 1100 1284 1107 1285
rect 1115 1284 1387 1285
rect 1125 1286 1240 1287
rect 1128 1288 1191 1289
rect 1072 1290 1192 1291
rect 1154 1292 1162 1293
rect 1044 1294 1156 1295
rect 1005 1296 1045 1297
rect 1184 1296 1252 1297
rect 1178 1298 1186 1299
rect 1166 1300 1180 1301
rect 1220 1300 1224 1301
rect 1202 1302 1222 1303
rect 1203 1304 1206 1305
rect 1224 1304 1384 1305
rect 1226 1306 1474 1307
rect 1088 1308 1228 1309
rect 1229 1308 1246 1309
rect 1121 1310 1231 1311
rect 1121 1312 1138 1313
rect 1235 1312 1487 1313
rect 1247 1314 1447 1315
rect 1253 1316 1498 1317
rect 1193 1318 1255 1319
rect 1148 1320 1195 1321
rect 1130 1322 1150 1323
rect 1131 1324 1176 1325
rect 1081 1326 1177 1327
rect 1262 1326 1285 1327
rect 1256 1328 1264 1329
rect 1274 1328 1282 1329
rect 1289 1328 1297 1329
rect 1079 1330 1291 1331
rect 1057 1332 1079 1333
rect 1056 1334 1104 1335
rect 1307 1334 1438 1335
rect 1308 1336 1426 1337
rect 1313 1338 1436 1339
rect 1325 1340 1405 1341
rect 1301 1342 1405 1343
rect 1302 1344 1462 1345
rect 1331 1346 1417 1347
rect 1319 1348 1333 1349
rect 1320 1350 1515 1351
rect 1337 1352 1345 1353
rect 1346 1352 1366 1353
rect 1347 1354 1356 1355
rect 1349 1356 1369 1357
rect 1356 1358 1381 1359
rect 1358 1360 1429 1361
rect 1383 1362 1411 1363
rect 1352 1364 1411 1365
rect 1353 1366 1377 1367
rect 1389 1366 1429 1367
rect 1389 1368 1505 1369
rect 1395 1370 1435 1371
rect 1398 1372 1432 1373
rect 1392 1374 1432 1375
rect 1401 1376 1444 1377
rect 1407 1378 1471 1379
rect 1304 1380 1408 1381
rect 1416 1380 1441 1381
rect 1422 1382 1465 1383
rect 1452 1384 1456 1385
rect 1413 1386 1453 1387
rect 1467 1386 1494 1387
rect 1008 1395 1054 1396
rect 1015 1397 1082 1398
rect 1019 1399 1125 1400
rect 1019 1401 1070 1402
rect 1038 1403 1067 1404
rect 998 1405 1067 1406
rect 1041 1407 1045 1408
rect 1053 1407 1094 1408
rect 1059 1409 1159 1410
rect 1063 1411 1192 1412
rect 1001 1413 1064 1414
rect 1000 1415 1051 1416
rect 1084 1415 1191 1416
rect 1088 1417 1195 1418
rect 1087 1419 1177 1420
rect 1106 1421 1122 1422
rect 1100 1423 1122 1424
rect 1118 1425 1228 1426
rect 1118 1427 1231 1428
rect 1143 1429 1167 1430
rect 1016 1431 1143 1432
rect 1146 1431 1170 1432
rect 1057 1433 1146 1434
rect 1173 1433 1188 1434
rect 1155 1435 1173 1436
rect 1149 1437 1155 1438
rect 1137 1439 1149 1440
rect 1131 1441 1137 1442
rect 1179 1441 1197 1442
rect 1178 1443 1341 1444
rect 1185 1445 1194 1446
rect 1199 1445 1357 1446
rect 1215 1447 1230 1448
rect 1217 1449 1225 1450
rect 1223 1451 1252 1452
rect 1226 1453 1240 1454
rect 1235 1455 1258 1456
rect 1128 1457 1257 1458
rect 1078 1459 1128 1460
rect 1241 1459 1305 1460
rect 1245 1461 1420 1462
rect 1254 1463 1335 1464
rect 1253 1465 1354 1466
rect 1260 1467 1378 1468
rect 1259 1469 1291 1470
rect 1263 1471 1287 1472
rect 1265 1473 1498 1474
rect 1284 1475 1450 1476
rect 1281 1477 1284 1478
rect 1308 1477 1419 1478
rect 1302 1479 1308 1480
rect 1310 1479 1348 1480
rect 1316 1481 1411 1482
rect 1320 1483 1374 1484
rect 1328 1485 1366 1486
rect 1332 1487 1515 1488
rect 1269 1489 1332 1490
rect 1337 1489 1408 1490
rect 1344 1491 1353 1492
rect 1346 1493 1390 1494
rect 1349 1495 1501 1496
rect 1355 1497 1429 1498
rect 1262 1499 1429 1500
rect 1358 1501 1432 1502
rect 1368 1503 1398 1504
rect 1370 1505 1435 1506
rect 1376 1507 1441 1508
rect 1296 1509 1440 1510
rect 1380 1511 1484 1512
rect 1379 1513 1444 1514
rect 1367 1515 1443 1516
rect 1388 1517 1453 1518
rect 1391 1519 1465 1520
rect 1394 1521 1468 1522
rect 1400 1523 1447 1524
rect 1404 1525 1487 1526
rect 1383 1527 1405 1528
rect 1407 1527 1474 1528
rect 1437 1529 1459 1530
rect 1455 1531 1508 1532
rect 1470 1533 1480 1534
rect 997 1542 1067 1543
rect 1016 1544 1082 1545
rect 1024 1546 1109 1547
rect 1031 1548 1039 1549
rect 1035 1550 1054 1551
rect 1026 1552 1035 1553
rect 1027 1554 1076 1555
rect 1041 1556 1176 1557
rect 1043 1558 1128 1559
rect 1052 1560 1242 1561
rect 1057 1562 1149 1563
rect 1056 1564 1155 1565
rect 1063 1566 1081 1567
rect 1068 1568 1088 1569
rect 1086 1570 1119 1571
rect 1019 1572 1118 1573
rect 1020 1574 1151 1575
rect 1100 1576 1227 1577
rect 1102 1578 1241 1579
rect 1124 1580 1148 1581
rect 1136 1582 1154 1583
rect 1160 1582 1184 1583
rect 1012 1584 1160 1585
rect 1169 1584 1199 1585
rect 1145 1586 1169 1587
rect 1172 1586 1205 1587
rect 1060 1588 1172 1589
rect 1059 1590 1136 1591
rect 1177 1590 1305 1591
rect 1187 1592 1247 1593
rect 1186 1594 1191 1595
rect 1074 1596 1190 1597
rect 1196 1596 1208 1597
rect 1166 1598 1196 1599
rect 1142 1600 1166 1601
rect 1201 1600 1224 1601
rect 1050 1602 1223 1603
rect 1217 1604 1232 1605
rect 1220 1606 1238 1607
rect 1193 1608 1220 1609
rect 1225 1608 1254 1609
rect 1229 1610 1253 1611
rect 1228 1612 1257 1613
rect 1235 1614 1337 1615
rect 1249 1616 1260 1617
rect 1262 1616 1313 1617
rect 1265 1618 1301 1619
rect 1243 1620 1265 1621
rect 1283 1620 1319 1621
rect 1286 1622 1295 1623
rect 1310 1622 1386 1623
rect 1316 1624 1335 1625
rect 1315 1626 1419 1627
rect 1333 1628 1377 1629
rect 1346 1630 1385 1631
rect 1345 1632 1356 1633
rect 1349 1634 1416 1635
rect 1348 1636 1359 1637
rect 1352 1638 1382 1639
rect 1340 1640 1352 1641
rect 1339 1642 1374 1643
rect 1331 1644 1373 1645
rect 1354 1646 1380 1647
rect 1367 1648 1397 1649
rect 1370 1650 1401 1651
rect 1328 1652 1370 1653
rect 1327 1654 1422 1655
rect 1388 1656 1406 1657
rect 1387 1658 1426 1659
rect 1391 1660 1400 1661
rect 1270 1662 1391 1663
rect 1394 1662 1403 1663
rect 1288 1664 1394 1665
rect 1407 1664 1423 1665
rect 1342 1666 1409 1667
rect 1006 1675 1196 1676
rect 1010 1677 1044 1678
rect 1013 1679 1151 1680
rect 1003 1681 1152 1682
rect 1017 1683 1050 1684
rect 1020 1685 1035 1686
rect 1009 1687 1020 1688
rect 1024 1687 1101 1688
rect 1030 1689 1205 1690
rect 1037 1691 1169 1692
rect 1059 1693 1069 1694
rect 1059 1695 1178 1696
rect 1062 1697 1081 1698
rect 1068 1699 1197 1700
rect 1077 1701 1179 1702
rect 1079 1703 1190 1704
rect 1083 1705 1121 1706
rect 1082 1707 1238 1708
rect 1097 1709 1109 1710
rect 1102 1711 1232 1712
rect 1105 1713 1308 1714
rect 1106 1715 1229 1716
rect 1115 1717 1118 1718
rect 1118 1719 1199 1720
rect 1127 1721 1136 1722
rect 1133 1723 1154 1724
rect 1139 1725 1148 1726
rect 1142 1727 1160 1728
rect 1056 1729 1161 1730
rect 1148 1731 1166 1732
rect 1154 1733 1172 1734
rect 1172 1735 1184 1736
rect 1175 1737 1187 1738
rect 1184 1739 1208 1740
rect 1187 1741 1223 1742
rect 1199 1743 1202 1744
rect 1202 1745 1226 1746
rect 1205 1747 1364 1748
rect 1208 1749 1247 1750
rect 1211 1751 1241 1752
rect 1219 1753 1236 1754
rect 1220 1755 1250 1756
rect 1229 1757 1337 1758
rect 1232 1759 1253 1760
rect 1265 1759 1346 1760
rect 1267 1761 1271 1762
rect 1268 1763 1299 1764
rect 1283 1765 1319 1766
rect 1288 1767 1293 1768
rect 1289 1769 1340 1770
rect 1294 1771 1305 1772
rect 1295 1773 1323 1774
rect 1300 1775 1391 1776
rect 1301 1777 1403 1778
rect 1310 1779 1313 1780
rect 1313 1781 1423 1782
rect 1315 1783 1326 1784
rect 1316 1785 1370 1786
rect 1319 1787 1373 1788
rect 1327 1789 1419 1790
rect 1328 1791 1406 1792
rect 1331 1793 1429 1794
rect 1333 1795 1355 1796
rect 1337 1797 1382 1798
rect 1334 1799 1382 1800
rect 1342 1801 1394 1802
rect 1348 1803 1367 1804
rect 1347 1805 1400 1806
rect 1354 1807 1388 1808
rect 1360 1809 1404 1810
rect 1363 1811 1389 1812
rect 1375 1813 1436 1814
rect 1378 1815 1443 1816
rect 1384 1817 1426 1818
rect 1396 1819 1439 1820
rect 1012 1828 1140 1829
rect 1012 1830 1020 1831
rect 1016 1832 1121 1833
rect 1023 1834 1031 1835
rect 1033 1834 1190 1835
rect 1040 1836 1130 1837
rect 1044 1838 1134 1839
rect 1047 1840 1128 1841
rect 1056 1842 1145 1843
rect 1059 1844 1188 1845
rect 1060 1846 1063 1847
rect 1063 1848 1161 1849
rect 1065 1850 1176 1851
rect 1066 1852 1214 1853
rect 1070 1854 1305 1855
rect 1080 1856 1302 1857
rect 1084 1858 1209 1859
rect 1103 1860 1127 1861
rect 1097 1862 1103 1863
rect 1096 1864 1101 1865
rect 1151 1864 1157 1865
rect 1154 1866 1175 1867
rect 1148 1868 1154 1869
rect 1142 1870 1148 1871
rect 1026 1872 1142 1873
rect 1165 1872 1203 1873
rect 1184 1874 1193 1875
rect 1183 1876 1208 1877
rect 1205 1878 1223 1879
rect 1217 1880 1233 1881
rect 1211 1882 1217 1883
rect 1210 1884 1221 1885
rect 1123 1886 1220 1887
rect 1229 1886 1236 1887
rect 1228 1888 1241 1889
rect 1249 1890 1296 1891
rect 1252 1892 1269 1893
rect 1255 1894 1290 1895
rect 1265 1896 1299 1897
rect 1264 1898 1280 1899
rect 1273 1900 1314 1901
rect 1276 1902 1308 1903
rect 1288 1904 1329 1905
rect 1292 1906 1341 1907
rect 1291 1908 1332 1909
rect 1294 1910 1358 1911
rect 1297 1912 1332 1913
rect 1303 1914 1320 1915
rect 1310 1916 1326 1917
rect 1199 1918 1325 1919
rect 1196 1920 1199 1921
rect 1178 1922 1196 1923
rect 1314 1922 1317 1923
rect 1334 1922 1341 1923
rect 1334 1924 1364 1925
rect 1337 1926 1404 1927
rect 1283 1928 1338 1929
rect 1347 1928 1382 1929
rect 1364 1930 1398 1931
rect 1375 1932 1392 1933
rect 1360 1934 1375 1935
rect 1378 1934 1389 1935
rect 997 1943 1010 1944
rect 1019 1943 1175 1944
rect 1012 1945 1020 1946
rect 1023 1945 1100 1946
rect 1023 1947 1121 1948
rect 1030 1949 1142 1950
rect 1033 1951 1130 1952
rect 1035 1953 1061 1954
rect 1052 1955 1097 1956
rect 1057 1957 1163 1958
rect 1059 1959 1193 1960
rect 1066 1961 1133 1962
rect 1087 1963 1214 1964
rect 1090 1965 1103 1966
rect 1093 1967 1145 1968
rect 1096 1969 1118 1970
rect 1102 1971 1199 1972
rect 1105 1973 1160 1974
rect 1114 1975 1175 1976
rect 1120 1977 1148 1978
rect 1126 1979 1154 1980
rect 1129 1981 1157 1982
rect 1141 1983 1217 1984
rect 1150 1985 1172 1986
rect 1070 1987 1172 1988
rect 1063 1989 1070 1990
rect 1153 1989 1196 1990
rect 1156 1991 1190 1992
rect 1183 1993 1211 1994
rect 1183 1995 1208 1996
rect 1195 1997 1220 1998
rect 1084 1999 1220 2000
rect 1045 2001 1085 2002
rect 1198 2001 1223 2002
rect 1165 2003 1223 2004
rect 1073 2005 1166 2006
rect 1201 2005 1241 2006
rect 1204 2007 1242 2008
rect 1213 2009 1259 2010
rect 1228 2011 1250 2012
rect 1232 2013 1256 2014
rect 1237 2015 1318 2016
rect 1247 2017 1292 2018
rect 1252 2019 1257 2020
rect 1229 2021 1254 2022
rect 1259 2021 1262 2022
rect 1226 2023 1263 2024
rect 1279 2023 1293 2024
rect 1264 2025 1281 2026
rect 1288 2025 1305 2026
rect 1294 2027 1362 2028
rect 1276 2029 1296 2030
rect 1277 2031 1315 2032
rect 1297 2033 1302 2034
rect 1298 2035 1358 2036
rect 1307 2037 1338 2038
rect 1323 2039 1354 2040
rect 1328 2041 1341 2042
rect 1334 2043 1344 2044
rect 1307 2045 1344 2046
rect 1367 2045 1378 2046
rect 1000 2054 1036 2055
rect 1016 2056 1097 2057
rect 1026 2058 1067 2059
rect 1034 2060 1094 2061
rect 1041 2062 1080 2063
rect 1043 2064 1157 2065
rect 1045 2066 1143 2067
rect 1048 2068 1085 2069
rect 1050 2070 1130 2071
rect 1052 2072 1172 2073
rect 1059 2074 1107 2075
rect 1082 2076 1146 2077
rect 1085 2078 1110 2079
rect 1094 2080 1100 2081
rect 1102 2080 1230 2081
rect 1090 2082 1104 2083
rect 1126 2082 1140 2083
rect 1073 2084 1128 2085
rect 1150 2084 1158 2085
rect 1162 2084 1170 2085
rect 1055 2086 1164 2087
rect 1165 2086 1173 2087
rect 1159 2088 1167 2089
rect 1153 2090 1161 2091
rect 1178 2090 1281 2091
rect 1183 2092 1227 2093
rect 1198 2094 1223 2095
rect 1201 2096 1224 2097
rect 1186 2098 1203 2099
rect 1204 2098 1227 2099
rect 1205 2100 1251 2101
rect 1232 2102 1236 2103
rect 1190 2104 1233 2105
rect 1244 2104 1311 2105
rect 1244 2106 1248 2107
rect 1253 2106 1269 2107
rect 1271 2106 1333 2107
rect 1274 2108 1344 2109
rect 1277 2110 1326 2111
rect 1199 2112 1278 2113
rect 1286 2112 1308 2113
rect 1213 2114 1308 2115
rect 1298 2116 1357 2117
rect 1292 2118 1299 2119
rect 1301 2118 1314 2119
rect 1295 2120 1302 2121
rect 1304 2120 1317 2121
rect 1319 2120 1341 2121
rect 1304 2122 1340 2123
rect 1323 2124 1347 2125
rect 1238 2126 1347 2127
rect 1015 2135 1095 2136
rect 1022 2137 1080 2138
rect 1025 2139 1104 2140
rect 1024 2141 1035 2142
rect 1031 2143 1041 2144
rect 1034 2145 1107 2146
rect 1037 2147 1140 2148
rect 1040 2149 1134 2150
rect 1044 2151 1158 2152
rect 1047 2153 1090 2154
rect 1062 2155 1096 2156
rect 1066 2157 1164 2158
rect 1065 2159 1132 2160
rect 1069 2161 1099 2162
rect 1056 2163 1070 2164
rect 1073 2163 1122 2164
rect 1079 2165 1213 2166
rect 1085 2167 1170 2168
rect 1092 2169 1143 2170
rect 1107 2171 1128 2172
rect 1109 2173 1141 2174
rect 1119 2175 1167 2176
rect 1125 2177 1173 2178
rect 1128 2179 1176 2180
rect 1137 2181 1146 2182
rect 1149 2181 1197 2182
rect 1154 2183 1216 2184
rect 1160 2185 1254 2186
rect 1164 2187 1200 2188
rect 1170 2189 1206 2190
rect 1176 2191 1203 2192
rect 1179 2193 1191 2194
rect 1188 2195 1227 2196
rect 1191 2197 1224 2198
rect 1200 2199 1351 2200
rect 1221 2201 1299 2202
rect 1225 2203 1266 2204
rect 1231 2205 1272 2206
rect 1241 2207 1251 2208
rect 1244 2209 1275 2210
rect 1247 2211 1302 2212
rect 1256 2213 1311 2214
rect 1259 2215 1323 2216
rect 1259 2217 1281 2218
rect 1262 2219 1305 2220
rect 1268 2221 1330 2222
rect 1235 2223 1269 2224
rect 1152 2225 1235 2226
rect 1271 2225 1317 2226
rect 1286 2227 1340 2228
rect 1238 2229 1288 2230
rect 1313 2229 1344 2230
rect 1319 2231 1347 2232
rect 1332 2233 1337 2234
rect 1021 2242 1035 2243
rect 1037 2242 1057 2243
rect 1044 2244 1096 2245
rect 1044 2246 1048 2247
rect 1051 2246 1272 2247
rect 1062 2248 1067 2249
rect 1069 2248 1129 2249
rect 1073 2250 1084 2251
rect 1086 2250 1189 2251
rect 1086 2252 1090 2253
rect 1089 2254 1093 2255
rect 1028 2256 1093 2257
rect 1027 2258 1138 2259
rect 1095 2260 1099 2261
rect 1079 2262 1099 2263
rect 1122 2262 1213 2263
rect 1131 2264 1156 2265
rect 1140 2266 1159 2267
rect 1143 2268 1180 2269
rect 1149 2270 1174 2271
rect 1125 2272 1150 2273
rect 1119 2274 1126 2275
rect 1080 2276 1120 2277
rect 1152 2276 1226 2277
rect 1107 2278 1153 2279
rect 1161 2278 1165 2279
rect 1170 2278 1205 2279
rect 1170 2280 1177 2281
rect 1176 2282 1227 2283
rect 1182 2284 1216 2285
rect 1194 2286 1208 2287
rect 1200 2288 1285 2289
rect 1167 2290 1201 2291
rect 1210 2290 1248 2291
rect 1213 2292 1232 2293
rect 1223 2294 1251 2295
rect 1259 2294 1278 2295
rect 1262 2296 1281 2297
rect 1274 2298 1288 2299
rect 1027 2307 1150 2308
rect 1037 2309 1090 2310
rect 1041 2311 1093 2312
rect 1027 2313 1093 2314
rect 1044 2315 1126 2316
rect 1051 2317 1074 2318
rect 1034 2319 1075 2320
rect 1034 2321 1153 2322
rect 1056 2323 1077 2324
rect 1044 2325 1078 2326
rect 1071 2327 1087 2328
rect 1080 2329 1096 2330
rect 1089 2331 1114 2332
rect 1095 2333 1099 2334
rect 1104 2333 1156 2334
rect 1110 2335 1159 2336
rect 1116 2337 1180 2338
rect 1119 2339 1165 2340
rect 1134 2341 1168 2342
rect 1143 2343 1156 2344
rect 1152 2345 1171 2346
rect 1158 2347 1192 2348
rect 1161 2349 1198 2350
rect 1122 2351 1162 2352
rect 1122 2353 1171 2354
rect 1173 2353 1183 2354
rect 1173 2355 1177 2356
rect 1176 2357 1183 2358
rect 1185 2357 1214 2358
rect 1200 2359 1211 2360
rect 1204 2361 1217 2362
rect 1232 2361 1240 2362
rect 1245 2361 1253 2362
rect 1030 2370 1084 2371
rect 1033 2372 1075 2373
rect 1041 2374 1063 2375
rect 1050 2376 1072 2377
rect 1053 2378 1096 2379
rect 1040 2380 1096 2381
rect 1059 2382 1078 2383
rect 1065 2384 1156 2385
rect 1068 2386 1090 2387
rect 1080 2388 1087 2389
rect 1037 2390 1087 2391
rect 1036 2392 1078 2393
rect 1092 2392 1102 2393
rect 1110 2392 1189 2393
rect 1116 2394 1150 2395
rect 1113 2396 1117 2397
rect 1104 2398 1114 2399
rect 1056 2400 1105 2401
rect 1122 2400 1126 2401
rect 1128 2400 1135 2401
rect 1137 2400 1174 2401
rect 1140 2402 1159 2403
rect 1161 2402 1171 2403
rect 1164 2404 1168 2405
rect 1176 2404 1192 2405
rect 1182 2406 1186 2407
rect 1033 2415 1084 2416
rect 1040 2417 1063 2418
rect 1039 2419 1060 2420
rect 1042 2421 1090 2422
rect 1045 2423 1078 2424
rect 1047 2425 1105 2426
rect 1048 2427 1055 2428
rect 1050 2429 1102 2430
rect 1058 2431 1114 2432
rect 1065 2433 1117 2434
rect 1072 2435 1138 2436
rect 1078 2437 1129 2438
rect 1086 2439 1120 2440
rect 1098 2441 1132 2442
rect 1122 2443 1141 2444
rect 1125 2445 1147 2446
rect 1143 2447 1150 2448
rect 1039 2456 1062 2457
rect 1045 2458 1049 2459
rect 1054 2458 1073 2459
rect 1058 2460 1079 2461
<< metal2 >>
rect 1028 497 1029 507
rect 1047 497 1048 507
rect 1038 499 1039 507
rect 1068 499 1069 507
rect 1041 501 1042 507
rect 1062 501 1063 507
rect 1050 503 1051 507
rect 1071 503 1072 507
rect 1074 503 1075 507
rect 1077 503 1078 507
rect 1084 503 1085 507
rect 1090 503 1091 507
rect 1099 503 1100 507
rect 1102 503 1103 507
rect 1132 503 1133 507
rect 1139 503 1140 507
rect 1021 511 1022 514
rect 1034 513 1035 558
rect 1031 511 1032 516
rect 1056 515 1057 558
rect 1044 511 1045 518
rect 1068 511 1069 518
rect 1047 511 1048 520
rect 1068 519 1069 558
rect 1046 521 1047 558
rect 1071 511 1072 522
rect 1050 511 1051 524
rect 1062 511 1063 524
rect 1028 511 1029 526
rect 1062 525 1063 558
rect 1053 511 1054 528
rect 1074 511 1075 528
rect 1028 529 1029 558
rect 1074 529 1075 558
rect 1031 531 1032 558
rect 1053 531 1054 558
rect 1077 511 1078 532
rect 1157 531 1158 558
rect 1021 533 1022 558
rect 1077 533 1078 558
rect 1080 511 1081 534
rect 1127 533 1128 558
rect 1087 511 1088 536
rect 1170 535 1171 558
rect 1090 511 1091 538
rect 1130 537 1131 558
rect 1090 539 1091 558
rect 1102 539 1103 558
rect 1093 511 1094 542
rect 1154 541 1155 558
rect 1099 511 1100 544
rect 1182 543 1183 558
rect 1087 545 1088 558
rect 1099 545 1100 558
rect 1105 545 1106 558
rect 1226 545 1227 558
rect 1112 547 1113 558
rect 1124 547 1125 558
rect 1115 549 1116 558
rect 1145 549 1146 558
rect 1142 551 1143 558
rect 1151 551 1152 558
rect 1164 551 1165 558
rect 1197 551 1198 558
rect 1167 553 1168 558
rect 1188 553 1189 558
rect 1200 553 1201 558
rect 1220 553 1221 558
rect 1203 555 1204 558
rect 1216 555 1217 558
rect 1229 555 1230 558
rect 1235 555 1236 558
rect 1009 564 1010 621
rect 1015 564 1016 621
rect 1024 562 1025 565
rect 1028 562 1029 565
rect 1028 566 1029 621
rect 1077 562 1078 567
rect 1032 568 1033 621
rect 1099 562 1100 569
rect 1034 562 1035 571
rect 1045 570 1046 621
rect 1039 572 1040 621
rect 1068 562 1069 573
rect 1043 562 1044 575
rect 1074 562 1075 575
rect 1042 576 1043 621
rect 1215 576 1216 621
rect 1056 562 1057 579
rect 1074 578 1075 621
rect 1057 580 1058 621
rect 1113 580 1114 621
rect 1062 562 1063 583
rect 1080 582 1081 621
rect 1061 584 1062 621
rect 1098 584 1099 621
rect 1064 586 1065 621
rect 1122 586 1123 621
rect 1071 588 1072 621
rect 1110 588 1111 621
rect 1083 562 1084 591
rect 1119 590 1120 621
rect 1025 592 1026 621
rect 1083 592 1084 621
rect 1086 592 1087 621
rect 1127 562 1128 593
rect 1102 562 1103 595
rect 1104 594 1105 621
rect 1115 562 1116 595
rect 1152 594 1153 621
rect 1130 562 1131 597
rect 1137 596 1138 621
rect 1124 562 1125 599
rect 1131 598 1132 621
rect 1154 562 1155 599
rect 1194 598 1195 621
rect 1145 562 1146 601
rect 1155 600 1156 621
rect 1170 562 1171 601
rect 1176 600 1177 621
rect 1173 602 1174 621
rect 1209 602 1210 621
rect 1182 562 1183 605
rect 1185 562 1186 605
rect 1182 606 1183 621
rect 1200 562 1201 607
rect 1203 562 1204 607
rect 1242 606 1243 621
rect 1148 562 1149 609
rect 1203 608 1204 621
rect 1089 610 1090 621
rect 1149 610 1150 621
rect 1206 562 1207 611
rect 1218 610 1219 621
rect 1142 562 1143 613
rect 1206 612 1207 621
rect 1223 562 1224 613
rect 1233 612 1234 621
rect 1226 562 1227 615
rect 1279 614 1280 621
rect 1220 562 1221 617
rect 1227 616 1228 621
rect 1229 562 1230 617
rect 1282 616 1283 621
rect 1197 562 1198 619
rect 1230 618 1231 621
rect 1021 625 1022 628
rect 1096 627 1097 714
rect 1035 625 1036 630
rect 1083 625 1084 630
rect 1015 625 1016 632
rect 1034 631 1035 714
rect 1039 625 1040 632
rect 1135 631 1136 714
rect 1049 633 1050 714
rect 1122 625 1123 634
rect 1052 635 1053 714
rect 1077 635 1078 714
rect 1054 625 1055 638
rect 1171 637 1172 714
rect 1057 625 1058 640
rect 1083 639 1084 714
rect 1061 625 1062 642
rect 1141 641 1142 714
rect 1045 625 1046 644
rect 1062 643 1063 714
rect 1064 625 1065 644
rect 1168 643 1169 714
rect 1071 645 1072 714
rect 1119 625 1120 646
rect 1074 625 1075 648
rect 1102 647 1103 714
rect 1080 625 1081 650
rect 1108 649 1109 714
rect 1040 651 1041 714
rect 1080 651 1081 714
rect 1089 625 1090 652
rect 1267 651 1268 714
rect 1090 653 1091 714
rect 1104 625 1105 654
rect 1098 625 1099 656
rect 1147 655 1148 714
rect 1113 625 1114 658
rect 1165 657 1166 714
rect 1114 659 1115 714
rect 1186 659 1187 714
rect 1117 661 1118 714
rect 1155 625 1156 662
rect 1125 625 1126 664
rect 1152 625 1153 664
rect 1110 625 1111 666
rect 1153 665 1154 714
rect 1025 625 1026 668
rect 1111 667 1112 714
rect 1024 669 1025 714
rect 1037 669 1038 714
rect 1126 669 1127 714
rect 1224 625 1225 670
rect 1128 625 1129 672
rect 1137 625 1138 672
rect 1042 625 1043 674
rect 1138 673 1139 714
rect 1149 625 1150 674
rect 1162 673 1163 714
rect 1173 625 1174 674
rect 1201 673 1202 714
rect 1174 675 1175 714
rect 1206 625 1207 676
rect 1176 625 1177 678
rect 1225 677 1226 714
rect 1189 679 1190 714
rect 1203 625 1204 680
rect 1192 681 1193 714
rect 1212 625 1213 682
rect 1194 625 1195 684
rect 1246 683 1247 714
rect 1204 685 1205 714
rect 1221 625 1222 686
rect 1207 687 1208 714
rect 1209 625 1210 688
rect 1131 625 1132 690
rect 1210 689 1211 714
rect 1213 689 1214 714
rect 1218 625 1219 690
rect 1215 625 1216 692
rect 1270 691 1271 714
rect 1219 693 1220 714
rect 1300 693 1301 714
rect 1227 625 1228 696
rect 1273 695 1274 714
rect 1233 625 1234 698
rect 1291 697 1292 714
rect 1242 625 1243 700
rect 1294 699 1295 714
rect 1259 625 1260 702
rect 1285 701 1286 714
rect 1276 703 1277 714
rect 1288 625 1289 704
rect 1230 625 1231 706
rect 1288 705 1289 714
rect 1182 625 1183 708
rect 1231 707 1232 714
rect 1279 625 1280 708
rect 1337 707 1338 714
rect 1279 709 1280 714
rect 1282 625 1283 710
rect 1198 711 1199 714
rect 1282 711 1283 714
rect 1297 711 1298 714
rect 1307 711 1308 714
rect 1334 711 1335 714
rect 1344 711 1345 714
rect 1015 720 1016 813
rect 1183 720 1184 813
rect 1018 722 1019 813
rect 1111 718 1112 723
rect 1021 718 1022 725
rect 1064 724 1065 813
rect 1031 718 1032 727
rect 1096 718 1097 727
rect 1028 718 1029 729
rect 1032 728 1033 813
rect 1034 718 1035 729
rect 1035 728 1036 813
rect 1049 718 1050 729
rect 1171 718 1172 729
rect 1048 730 1049 813
rect 1177 730 1178 813
rect 1059 718 1060 733
rect 1080 718 1081 733
rect 1062 718 1063 735
rect 1067 734 1068 813
rect 1071 718 1072 735
rect 1165 718 1166 735
rect 1070 736 1071 813
rect 1195 736 1196 813
rect 1074 718 1075 739
rect 1159 738 1160 813
rect 1090 718 1091 741
rect 1165 740 1166 813
rect 1077 718 1078 743
rect 1089 742 1090 813
rect 1102 718 1103 743
rect 1120 742 1121 813
rect 1105 744 1106 813
rect 1153 718 1154 745
rect 1041 746 1042 813
rect 1153 746 1154 813
rect 1108 718 1109 749
rect 1117 748 1118 813
rect 1114 718 1115 751
rect 1162 718 1163 751
rect 1129 752 1130 813
rect 1141 718 1142 753
rect 1138 718 1139 755
rect 1156 754 1157 813
rect 1186 718 1187 755
rect 1243 754 1244 813
rect 1126 718 1127 757
rect 1186 756 1187 813
rect 1192 718 1193 757
rect 1249 756 1250 813
rect 1198 718 1199 759
rect 1228 758 1229 813
rect 1168 718 1169 761
rect 1198 760 1199 813
rect 1083 718 1084 763
rect 1168 762 1169 813
rect 1201 718 1202 763
rect 1252 762 1253 813
rect 1204 718 1205 765
rect 1261 764 1262 813
rect 1213 718 1214 767
rect 1285 718 1286 767
rect 1225 718 1226 769
rect 1285 768 1286 813
rect 1052 770 1053 813
rect 1225 770 1226 813
rect 1240 770 1241 813
rect 1433 770 1434 813
rect 1255 772 1256 813
rect 1366 772 1367 813
rect 1267 718 1268 775
rect 1357 774 1358 813
rect 1246 718 1247 777
rect 1267 776 1268 813
rect 1189 718 1190 779
rect 1246 778 1247 813
rect 1073 780 1074 813
rect 1189 780 1190 813
rect 1270 718 1271 781
rect 1360 780 1361 813
rect 1273 718 1274 783
rect 1375 782 1376 813
rect 1207 718 1208 785
rect 1273 784 1274 813
rect 1174 718 1175 787
rect 1207 786 1208 813
rect 1276 718 1277 787
rect 1339 786 1340 813
rect 1279 718 1280 789
rect 1342 788 1343 813
rect 1219 718 1220 791
rect 1279 790 1280 813
rect 1288 718 1289 791
rect 1410 790 1411 813
rect 1294 718 1295 793
rect 1387 792 1388 813
rect 1297 718 1298 795
rect 1327 794 1328 813
rect 1303 718 1304 797
rect 1321 796 1322 813
rect 1291 718 1292 799
rect 1303 798 1304 813
rect 1234 800 1235 813
rect 1291 800 1292 813
rect 1307 718 1308 801
rect 1390 800 1391 813
rect 1231 718 1232 803
rect 1306 802 1307 813
rect 1324 718 1325 803
rect 1348 802 1349 813
rect 1334 718 1335 805
rect 1427 804 1428 813
rect 1310 718 1311 807
rect 1333 806 1334 813
rect 1344 718 1345 807
rect 1350 718 1351 807
rect 1345 808 1346 813
rect 1407 808 1408 813
rect 1378 810 1379 813
rect 1384 810 1385 813
rect 955 819 956 960
rect 962 819 963 960
rect 993 819 994 960
rect 1035 817 1036 820
rect 1012 821 1013 960
rect 1026 821 1027 960
rect 1016 823 1017 960
rect 1064 817 1065 824
rect 1029 817 1030 826
rect 1132 825 1133 960
rect 1019 827 1020 960
rect 1030 827 1031 960
rect 1038 817 1039 828
rect 1052 817 1053 828
rect 1033 829 1034 960
rect 1037 829 1038 960
rect 1052 829 1053 960
rect 1067 817 1068 830
rect 1055 817 1056 832
rect 1306 817 1307 832
rect 1058 833 1059 960
rect 1135 817 1136 834
rect 1065 835 1066 960
rect 1162 835 1163 960
rect 1068 837 1069 960
rect 1089 817 1090 838
rect 1070 817 1071 840
rect 1177 817 1178 840
rect 1071 841 1072 960
rect 1393 841 1394 960
rect 1077 817 1078 844
rect 1189 817 1190 844
rect 1078 845 1079 960
rect 1324 845 1325 960
rect 1080 817 1081 848
rect 1095 817 1096 848
rect 1090 849 1091 960
rect 1117 817 1118 850
rect 1105 817 1106 852
rect 1276 851 1277 960
rect 1108 853 1109 960
rect 1183 817 1184 854
rect 1120 817 1121 856
rect 1135 855 1136 960
rect 1009 857 1010 960
rect 1120 857 1121 960
rect 1123 857 1124 960
rect 1186 817 1187 858
rect 1129 817 1130 860
rect 1201 859 1202 960
rect 1138 861 1139 960
rect 1147 817 1148 862
rect 1144 863 1145 960
rect 1153 817 1154 864
rect 1147 865 1148 960
rect 1156 817 1157 866
rect 1074 867 1075 960
rect 1156 867 1157 960
rect 1150 869 1151 960
rect 1225 817 1226 870
rect 1159 817 1160 872
rect 1264 871 1265 960
rect 1165 817 1166 874
rect 1213 873 1214 960
rect 1048 817 1049 876
rect 1165 875 1166 960
rect 1022 817 1023 878
rect 1049 877 1050 960
rect 1174 877 1175 960
rect 1240 817 1241 878
rect 1183 879 1184 960
rect 1381 817 1382 880
rect 1189 881 1190 960
rect 1261 817 1262 882
rect 1198 817 1199 884
rect 1204 883 1205 960
rect 1207 817 1208 884
rect 1306 883 1307 960
rect 1219 885 1220 960
rect 1285 817 1286 886
rect 1225 887 1226 960
rect 1249 817 1250 888
rect 1228 817 1229 890
rect 1294 817 1295 890
rect 1234 817 1235 892
rect 1258 891 1259 960
rect 1243 817 1244 894
rect 1309 893 1310 960
rect 1243 895 1244 960
rect 1342 817 1343 896
rect 1246 817 1247 898
rect 1363 817 1364 898
rect 1249 899 1250 960
rect 1447 817 1448 900
rect 1252 817 1253 902
rect 1366 901 1367 960
rect 1252 903 1253 960
rect 1279 817 1280 904
rect 1168 817 1169 906
rect 1279 905 1280 960
rect 1168 907 1169 960
rect 1195 817 1196 908
rect 1195 909 1196 960
rect 1439 909 1440 960
rect 1255 817 1256 912
rect 1384 817 1385 912
rect 1267 817 1268 914
rect 1414 913 1415 960
rect 1270 915 1271 960
rect 1473 915 1474 960
rect 1282 917 1283 960
rect 1300 917 1301 960
rect 1318 917 1319 960
rect 1417 817 1418 918
rect 1321 817 1322 920
rect 1400 817 1401 920
rect 1321 921 1322 960
rect 1348 817 1349 922
rect 1207 923 1208 960
rect 1348 923 1349 960
rect 1327 923 1328 960
rect 1327 817 1328 924
rect 1333 923 1334 960
rect 1333 817 1334 924
rect 1339 817 1340 926
rect 1354 925 1355 960
rect 1351 927 1352 960
rect 1469 927 1470 960
rect 1357 817 1358 930
rect 1369 929 1370 960
rect 1360 817 1361 932
rect 1372 931 1373 960
rect 1363 933 1364 960
rect 1384 933 1385 960
rect 1375 817 1376 936
rect 1399 935 1400 960
rect 1378 817 1379 938
rect 1402 937 1403 960
rect 1387 817 1388 940
rect 1405 939 1406 960
rect 1387 941 1388 960
rect 1410 817 1411 942
rect 1273 817 1274 944
rect 1411 943 1412 960
rect 1390 817 1391 946
rect 1408 945 1409 960
rect 1303 817 1304 948
rect 1390 947 1391 960
rect 1396 817 1397 948
rect 1432 947 1433 960
rect 1345 817 1346 950
rect 1396 949 1397 960
rect 1102 817 1103 952
rect 1345 951 1346 960
rect 1423 951 1424 960
rect 1460 951 1461 960
rect 1427 817 1428 954
rect 1463 953 1464 960
rect 1426 955 1427 960
rect 1457 955 1458 960
rect 1437 817 1438 958
rect 1444 817 1445 958
rect 979 964 980 967
rect 986 964 987 967
rect 989 964 990 967
rect 993 964 994 967
rect 1009 966 1010 1093
rect 1009 964 1010 967
rect 1012 964 1013 967
rect 1108 964 1109 967
rect 1019 964 1020 969
rect 1120 964 1121 969
rect 1023 964 1024 971
rect 1049 964 1050 971
rect 1026 964 1027 973
rect 1132 964 1133 973
rect 1030 964 1031 975
rect 1055 964 1056 975
rect 1030 976 1031 1093
rect 1162 964 1163 977
rect 1033 978 1034 1093
rect 1171 978 1172 1093
rect 1050 980 1051 1093
rect 1052 964 1053 981
rect 1068 964 1069 981
rect 1072 980 1073 1093
rect 1074 964 1075 981
rect 1309 964 1310 981
rect 1037 964 1038 983
rect 1075 982 1076 1093
rect 1037 984 1038 1093
rect 1078 964 1079 985
rect 1090 964 1091 985
rect 1102 984 1103 1093
rect 1090 986 1091 1093
rect 1276 964 1277 987
rect 1105 988 1106 1093
rect 1135 964 1136 989
rect 1120 990 1121 1093
rect 1123 964 1124 991
rect 1129 990 1130 1093
rect 1138 964 1139 991
rect 1135 992 1136 1093
rect 1144 964 1145 993
rect 1141 994 1142 1093
rect 1201 964 1202 995
rect 1147 964 1148 997
rect 1186 996 1187 1093
rect 1147 998 1148 1093
rect 1264 964 1265 999
rect 1153 1000 1154 1093
rect 1168 964 1169 1001
rect 1159 1002 1160 1093
rect 1213 964 1214 1003
rect 1066 1004 1067 1093
rect 1213 1004 1214 1093
rect 1165 964 1166 1007
rect 1192 1006 1193 1093
rect 1156 964 1157 1009
rect 1165 1008 1166 1093
rect 1156 1010 1157 1093
rect 1204 964 1205 1011
rect 1174 964 1175 1013
rect 1216 1012 1217 1093
rect 1177 1014 1178 1093
rect 1436 964 1437 1015
rect 1183 964 1184 1017
rect 1240 1016 1241 1093
rect 1047 1018 1048 1093
rect 1183 1018 1184 1093
rect 1189 964 1190 1019
rect 1228 1018 1229 1093
rect 1150 964 1151 1021
rect 1189 1020 1190 1093
rect 1195 964 1196 1021
rect 1234 1020 1235 1093
rect 1195 1022 1196 1093
rect 1201 1022 1202 1093
rect 1198 1024 1199 1093
rect 1279 964 1280 1025
rect 1207 964 1208 1027
rect 1246 1026 1247 1093
rect 1243 964 1244 1029
rect 1294 1028 1295 1093
rect 1249 964 1250 1031
rect 1291 1030 1292 1093
rect 1258 964 1259 1033
rect 1264 1032 1265 1093
rect 1225 964 1226 1035
rect 1258 1034 1259 1093
rect 1270 964 1271 1035
rect 1312 1034 1313 1093
rect 1276 1036 1277 1093
rect 1458 1036 1459 1093
rect 1282 964 1283 1039
rect 1285 1038 1286 1093
rect 1300 1038 1301 1093
rect 1324 964 1325 1039
rect 1306 964 1307 1041
rect 1384 964 1385 1041
rect 1327 964 1328 1043
rect 1336 1042 1337 1093
rect 1333 964 1334 1045
rect 1342 1044 1343 1093
rect 1348 1044 1349 1093
rect 1396 964 1397 1045
rect 1354 964 1355 1047
rect 1476 964 1477 1047
rect 1318 964 1319 1049
rect 1354 1048 1355 1093
rect 1318 1050 1319 1093
rect 1363 964 1364 1051
rect 1357 1052 1358 1093
rect 1408 964 1409 1053
rect 1375 1054 1376 1093
rect 1414 964 1415 1055
rect 1387 964 1388 1057
rect 1449 1056 1450 1093
rect 1369 964 1370 1059
rect 1387 1058 1388 1093
rect 1369 1060 1370 1093
rect 1469 964 1470 1061
rect 1390 964 1391 1063
rect 1455 1062 1456 1093
rect 1372 964 1373 1065
rect 1390 1064 1391 1093
rect 1351 964 1352 1067
rect 1372 1066 1373 1093
rect 1321 964 1322 1069
rect 1351 1068 1352 1093
rect 1321 1070 1322 1093
rect 1366 964 1367 1071
rect 1402 964 1403 1071
rect 1418 1070 1419 1093
rect 1222 1072 1223 1093
rect 1403 1072 1404 1093
rect 1405 964 1406 1073
rect 1409 1072 1410 1093
rect 1399 964 1400 1075
rect 1406 1074 1407 1093
rect 1330 1076 1331 1093
rect 1400 1076 1401 1093
rect 1412 1076 1413 1093
rect 1432 964 1433 1077
rect 1423 964 1424 1079
rect 1443 1078 1444 1093
rect 1252 964 1253 1081
rect 1422 1080 1423 1093
rect 1252 1082 1253 1093
rect 1475 1082 1476 1093
rect 1426 964 1427 1085
rect 1428 1084 1429 1093
rect 1440 1084 1441 1093
rect 1460 964 1461 1085
rect 1219 964 1220 1087
rect 1461 1086 1462 1093
rect 1081 964 1082 1089
rect 1219 1088 1220 1093
rect 1452 1088 1453 1093
rect 1466 964 1467 1089
rect 1463 964 1464 1091
rect 1465 1090 1466 1093
rect 1006 1099 1007 1254
rect 1035 1099 1036 1254
rect 1012 1097 1013 1102
rect 1057 1101 1058 1254
rect 1013 1103 1014 1254
rect 1054 1103 1055 1254
rect 1033 1097 1034 1106
rect 1156 1097 1157 1106
rect 1037 1097 1038 1108
rect 1118 1107 1119 1254
rect 1040 1097 1041 1110
rect 1072 1097 1073 1110
rect 1041 1111 1042 1254
rect 1060 1111 1061 1254
rect 1047 1097 1048 1114
rect 1075 1097 1076 1114
rect 1048 1115 1049 1254
rect 1115 1115 1116 1254
rect 1050 1097 1051 1118
rect 1066 1117 1067 1254
rect 1062 1097 1063 1120
rect 1192 1097 1193 1120
rect 1069 1097 1070 1122
rect 1141 1097 1142 1122
rect 1038 1123 1039 1254
rect 1069 1123 1070 1254
rect 1076 1123 1077 1254
rect 1243 1097 1244 1124
rect 1078 1097 1079 1126
rect 1383 1125 1384 1254
rect 1081 1097 1082 1128
rect 1147 1097 1148 1128
rect 1094 1129 1095 1254
rect 1105 1097 1106 1130
rect 1100 1131 1101 1254
rect 1102 1097 1103 1132
rect 1019 1097 1020 1134
rect 1103 1133 1104 1254
rect 1020 1135 1021 1254
rect 1264 1097 1265 1136
rect 1106 1137 1107 1254
rect 1120 1097 1121 1138
rect 1026 1097 1027 1140
rect 1121 1139 1122 1254
rect 1109 1141 1110 1254
rect 1195 1097 1196 1142
rect 1129 1097 1130 1144
rect 1204 1097 1205 1144
rect 1135 1097 1136 1146
rect 1175 1145 1176 1254
rect 1148 1147 1149 1254
rect 1171 1097 1172 1148
rect 1153 1097 1154 1150
rect 1226 1149 1227 1254
rect 1154 1151 1155 1254
rect 1422 1097 1423 1152
rect 1165 1097 1166 1154
rect 1181 1153 1182 1254
rect 1166 1155 1167 1254
rect 1177 1097 1178 1156
rect 1172 1157 1173 1254
rect 1183 1097 1184 1158
rect 1090 1097 1091 1160
rect 1184 1159 1185 1254
rect 1178 1161 1179 1254
rect 1189 1097 1190 1162
rect 1159 1097 1160 1164
rect 1190 1163 1191 1254
rect 1063 1165 1064 1254
rect 1160 1165 1161 1254
rect 1186 1097 1187 1166
rect 1211 1165 1212 1254
rect 1193 1167 1194 1254
rect 1198 1097 1199 1168
rect 1201 1097 1202 1168
rect 1213 1097 1214 1168
rect 1044 1097 1045 1170
rect 1202 1169 1203 1254
rect 1044 1171 1045 1254
rect 1130 1171 1131 1254
rect 1205 1171 1206 1254
rect 1216 1097 1217 1172
rect 1214 1173 1215 1254
rect 1222 1097 1223 1174
rect 1219 1097 1220 1176
rect 1220 1175 1221 1254
rect 1228 1097 1229 1176
rect 1400 1097 1401 1176
rect 1229 1177 1230 1254
rect 1246 1097 1247 1178
rect 1234 1097 1235 1180
rect 1425 1097 1426 1180
rect 1235 1181 1236 1254
rect 1252 1097 1253 1182
rect 1247 1183 1248 1254
rect 1285 1097 1286 1184
rect 1253 1185 1254 1254
rect 1276 1097 1277 1186
rect 1256 1187 1257 1254
rect 1455 1097 1456 1188
rect 1262 1189 1263 1254
rect 1300 1097 1301 1190
rect 1268 1191 1269 1254
rect 1294 1097 1295 1192
rect 1274 1193 1275 1254
rect 1291 1097 1292 1194
rect 1289 1195 1290 1254
rect 1312 1097 1313 1196
rect 1301 1197 1302 1254
rect 1396 1097 1397 1198
rect 1304 1199 1305 1254
rect 1321 1097 1322 1200
rect 1307 1201 1308 1254
rect 1336 1097 1337 1202
rect 1313 1203 1314 1254
rect 1342 1097 1343 1204
rect 1318 1097 1319 1206
rect 1393 1097 1394 1206
rect 1319 1207 1320 1254
rect 1330 1097 1331 1208
rect 1325 1209 1326 1254
rect 1416 1209 1417 1254
rect 1331 1211 1332 1254
rect 1390 1097 1391 1212
rect 1337 1213 1338 1254
rect 1354 1097 1355 1214
rect 1346 1215 1347 1254
rect 1369 1097 1370 1216
rect 1351 1097 1352 1218
rect 1355 1217 1356 1254
rect 1348 1097 1349 1220
rect 1352 1219 1353 1254
rect 1349 1221 1350 1254
rect 1372 1097 1373 1222
rect 1357 1097 1358 1224
rect 1431 1223 1432 1254
rect 1358 1225 1359 1254
rect 1375 1097 1376 1226
rect 1258 1097 1259 1228
rect 1376 1227 1377 1254
rect 1389 1227 1390 1254
rect 1406 1097 1407 1228
rect 1392 1229 1393 1254
rect 1446 1097 1447 1230
rect 1395 1231 1396 1254
rect 1409 1097 1410 1232
rect 1387 1097 1388 1234
rect 1410 1233 1411 1254
rect 1386 1235 1387 1254
rect 1443 1097 1444 1236
rect 1398 1237 1399 1254
rect 1412 1097 1413 1238
rect 1401 1239 1402 1254
rect 1418 1097 1419 1240
rect 1404 1241 1405 1254
rect 1425 1241 1426 1254
rect 1407 1243 1408 1254
rect 1475 1097 1476 1244
rect 1413 1245 1414 1254
rect 1428 1097 1429 1246
rect 1422 1247 1423 1254
rect 1452 1097 1453 1248
rect 1438 1249 1439 1254
rect 1465 1097 1466 1250
rect 1440 1097 1441 1252
rect 1472 1097 1473 1252
rect 994 1260 995 1389
rect 998 1260 999 1389
rect 1006 1258 1007 1261
rect 1051 1258 1052 1261
rect 1013 1258 1014 1263
rect 1029 1262 1030 1389
rect 1020 1258 1021 1265
rect 1143 1264 1144 1389
rect 1008 1266 1009 1389
rect 1019 1266 1020 1389
rect 1022 1266 1023 1389
rect 1158 1266 1159 1389
rect 1026 1268 1027 1389
rect 1118 1258 1119 1269
rect 1035 1258 1036 1271
rect 1050 1270 1051 1389
rect 1066 1258 1067 1271
rect 1211 1258 1212 1271
rect 1069 1258 1070 1273
rect 1181 1258 1182 1273
rect 1010 1258 1011 1275
rect 1069 1274 1070 1389
rect 1076 1258 1077 1275
rect 1208 1258 1209 1275
rect 1054 1258 1055 1277
rect 1075 1276 1076 1389
rect 1038 1258 1039 1279
rect 1053 1278 1054 1389
rect 1091 1278 1092 1389
rect 1160 1258 1161 1279
rect 1094 1258 1095 1281
rect 1260 1280 1261 1389
rect 1106 1258 1107 1283
rect 1146 1282 1147 1389
rect 1100 1258 1101 1285
rect 1106 1284 1107 1389
rect 1115 1258 1116 1285
rect 1386 1258 1387 1285
rect 1125 1286 1126 1389
rect 1239 1286 1240 1389
rect 1128 1288 1129 1389
rect 1190 1258 1191 1289
rect 1072 1258 1073 1291
rect 1191 1290 1192 1389
rect 1154 1258 1155 1293
rect 1161 1292 1162 1389
rect 1044 1258 1045 1295
rect 1155 1294 1156 1389
rect 1005 1296 1006 1389
rect 1044 1296 1045 1389
rect 1172 1258 1173 1297
rect 1173 1296 1174 1389
rect 1184 1258 1185 1297
rect 1251 1296 1252 1389
rect 1178 1258 1179 1299
rect 1185 1298 1186 1389
rect 1166 1258 1167 1301
rect 1179 1300 1180 1389
rect 1214 1258 1215 1301
rect 1215 1300 1216 1389
rect 1220 1258 1221 1301
rect 1223 1258 1224 1301
rect 1202 1258 1203 1303
rect 1221 1302 1222 1389
rect 1203 1304 1204 1389
rect 1205 1258 1206 1305
rect 1224 1304 1225 1389
rect 1383 1258 1384 1305
rect 1226 1258 1227 1307
rect 1473 1306 1474 1389
rect 1088 1308 1089 1389
rect 1227 1308 1228 1389
rect 1229 1258 1230 1309
rect 1245 1308 1246 1389
rect 1121 1258 1122 1311
rect 1230 1310 1231 1389
rect 1121 1312 1122 1389
rect 1137 1312 1138 1389
rect 1235 1258 1236 1313
rect 1486 1312 1487 1389
rect 1247 1258 1248 1315
rect 1446 1314 1447 1389
rect 1253 1258 1254 1317
rect 1497 1316 1498 1389
rect 1193 1258 1194 1319
rect 1254 1318 1255 1389
rect 1148 1258 1149 1321
rect 1194 1320 1195 1389
rect 1130 1258 1131 1323
rect 1149 1322 1150 1389
rect 1131 1324 1132 1389
rect 1175 1258 1176 1325
rect 1081 1326 1082 1389
rect 1176 1326 1177 1389
rect 1262 1258 1263 1327
rect 1284 1326 1285 1389
rect 1256 1258 1257 1329
rect 1263 1328 1264 1389
rect 1268 1258 1269 1329
rect 1269 1328 1270 1389
rect 1274 1258 1275 1329
rect 1281 1328 1282 1389
rect 1289 1258 1290 1329
rect 1296 1328 1297 1389
rect 1079 1258 1080 1331
rect 1290 1330 1291 1389
rect 1057 1258 1058 1333
rect 1078 1332 1079 1389
rect 1056 1334 1057 1389
rect 1103 1258 1104 1335
rect 1307 1258 1308 1335
rect 1437 1334 1438 1389
rect 1308 1336 1309 1389
rect 1425 1258 1426 1337
rect 1313 1258 1314 1339
rect 1435 1258 1436 1339
rect 1325 1258 1326 1341
rect 1404 1258 1405 1341
rect 1301 1258 1302 1343
rect 1404 1342 1405 1389
rect 1302 1344 1303 1389
rect 1461 1344 1462 1389
rect 1331 1258 1332 1347
rect 1416 1258 1417 1347
rect 1319 1258 1320 1349
rect 1332 1348 1333 1389
rect 1320 1350 1321 1389
rect 1514 1350 1515 1389
rect 1337 1258 1338 1353
rect 1344 1352 1345 1389
rect 1346 1258 1347 1353
rect 1365 1352 1366 1389
rect 1347 1354 1348 1389
rect 1355 1258 1356 1355
rect 1349 1258 1350 1357
rect 1368 1356 1369 1389
rect 1356 1358 1357 1389
rect 1380 1358 1381 1389
rect 1358 1258 1359 1361
rect 1428 1258 1429 1361
rect 1383 1362 1384 1389
rect 1410 1258 1411 1363
rect 1352 1258 1353 1365
rect 1410 1364 1411 1389
rect 1353 1366 1354 1389
rect 1376 1258 1377 1367
rect 1389 1258 1390 1367
rect 1428 1366 1429 1389
rect 1389 1368 1390 1389
rect 1504 1368 1505 1389
rect 1395 1258 1396 1371
rect 1434 1370 1435 1389
rect 1398 1258 1399 1373
rect 1431 1258 1432 1373
rect 1392 1258 1393 1375
rect 1431 1374 1432 1389
rect 1401 1258 1402 1377
rect 1443 1376 1444 1389
rect 1407 1258 1408 1379
rect 1470 1378 1471 1389
rect 1304 1258 1305 1381
rect 1407 1380 1408 1389
rect 1416 1380 1417 1389
rect 1440 1380 1441 1389
rect 1422 1258 1423 1383
rect 1464 1382 1465 1389
rect 1452 1258 1453 1385
rect 1455 1384 1456 1389
rect 1413 1258 1414 1387
rect 1452 1386 1453 1389
rect 1467 1386 1468 1389
rect 1493 1386 1494 1389
rect 1008 1393 1009 1396
rect 1053 1393 1054 1396
rect 1015 1393 1016 1398
rect 1081 1397 1082 1536
rect 1019 1393 1020 1400
rect 1124 1399 1125 1536
rect 1019 1401 1020 1536
rect 1069 1393 1070 1402
rect 1038 1403 1039 1536
rect 1066 1393 1067 1404
rect 998 1393 999 1406
rect 1066 1405 1067 1536
rect 1041 1407 1042 1536
rect 1044 1393 1045 1408
rect 1053 1407 1054 1536
rect 1093 1407 1094 1536
rect 1059 1393 1060 1410
rect 1158 1393 1159 1410
rect 1063 1393 1064 1412
rect 1191 1393 1192 1412
rect 1001 1393 1002 1414
rect 1063 1413 1064 1536
rect 1000 1415 1001 1536
rect 1050 1393 1051 1416
rect 1075 1415 1076 1536
rect 1075 1393 1076 1416
rect 1084 1393 1085 1416
rect 1190 1415 1191 1536
rect 1088 1393 1089 1418
rect 1194 1393 1195 1418
rect 1087 1419 1088 1536
rect 1176 1393 1177 1420
rect 1106 1393 1107 1422
rect 1121 1393 1122 1422
rect 1100 1423 1101 1536
rect 1121 1423 1122 1536
rect 1118 1393 1119 1426
rect 1227 1393 1228 1426
rect 1118 1427 1119 1536
rect 1230 1393 1231 1428
rect 1143 1393 1144 1430
rect 1166 1429 1167 1536
rect 1016 1431 1017 1536
rect 1142 1431 1143 1536
rect 1146 1393 1147 1432
rect 1169 1431 1170 1536
rect 1057 1433 1058 1536
rect 1145 1433 1146 1536
rect 1160 1433 1161 1536
rect 1161 1393 1162 1434
rect 1173 1393 1174 1434
rect 1187 1433 1188 1536
rect 1155 1393 1156 1436
rect 1172 1435 1173 1536
rect 1149 1393 1150 1438
rect 1154 1437 1155 1536
rect 1137 1393 1138 1440
rect 1148 1439 1149 1536
rect 1131 1393 1132 1442
rect 1136 1441 1137 1536
rect 1179 1393 1180 1442
rect 1196 1441 1197 1536
rect 1178 1443 1179 1536
rect 1340 1443 1341 1536
rect 1185 1393 1186 1446
rect 1193 1445 1194 1536
rect 1199 1445 1200 1536
rect 1356 1393 1357 1446
rect 1215 1393 1216 1448
rect 1229 1447 1230 1536
rect 1217 1449 1218 1536
rect 1224 1393 1225 1450
rect 1223 1451 1224 1536
rect 1251 1393 1252 1452
rect 1226 1453 1227 1536
rect 1239 1393 1240 1454
rect 1235 1455 1236 1536
rect 1257 1393 1258 1456
rect 1128 1393 1129 1458
rect 1256 1457 1257 1536
rect 1078 1393 1079 1460
rect 1127 1459 1128 1536
rect 1241 1459 1242 1536
rect 1304 1459 1305 1536
rect 1245 1393 1246 1462
rect 1419 1393 1420 1462
rect 1254 1393 1255 1464
rect 1334 1463 1335 1536
rect 1253 1465 1254 1536
rect 1353 1393 1354 1466
rect 1260 1393 1261 1468
rect 1377 1393 1378 1468
rect 1259 1469 1260 1536
rect 1290 1393 1291 1470
rect 1263 1393 1264 1472
rect 1286 1471 1287 1536
rect 1265 1473 1266 1536
rect 1497 1393 1498 1474
rect 1284 1393 1285 1476
rect 1449 1393 1450 1476
rect 1281 1393 1282 1478
rect 1283 1477 1284 1536
rect 1308 1393 1309 1478
rect 1418 1477 1419 1536
rect 1302 1393 1303 1480
rect 1307 1479 1308 1536
rect 1310 1479 1311 1536
rect 1347 1393 1348 1480
rect 1316 1481 1317 1536
rect 1410 1393 1411 1482
rect 1320 1393 1321 1484
rect 1373 1483 1374 1536
rect 1328 1485 1329 1536
rect 1365 1393 1366 1486
rect 1332 1393 1333 1488
rect 1514 1393 1515 1488
rect 1269 1393 1270 1490
rect 1331 1489 1332 1536
rect 1337 1489 1338 1536
rect 1407 1393 1408 1490
rect 1344 1393 1345 1492
rect 1352 1491 1353 1536
rect 1346 1493 1347 1536
rect 1389 1393 1390 1494
rect 1349 1495 1350 1536
rect 1500 1393 1501 1496
rect 1355 1497 1356 1536
rect 1428 1393 1429 1498
rect 1262 1499 1263 1536
rect 1428 1499 1429 1536
rect 1358 1501 1359 1536
rect 1431 1393 1432 1502
rect 1368 1393 1369 1504
rect 1397 1503 1398 1536
rect 1370 1505 1371 1536
rect 1434 1393 1435 1506
rect 1376 1507 1377 1536
rect 1440 1393 1441 1508
rect 1296 1393 1297 1510
rect 1439 1509 1440 1536
rect 1380 1393 1381 1512
rect 1483 1393 1484 1512
rect 1379 1513 1380 1536
rect 1443 1393 1444 1514
rect 1367 1515 1368 1536
rect 1442 1515 1443 1536
rect 1388 1517 1389 1536
rect 1452 1393 1453 1518
rect 1391 1519 1392 1536
rect 1464 1393 1465 1520
rect 1394 1521 1395 1536
rect 1467 1393 1468 1522
rect 1400 1523 1401 1536
rect 1446 1393 1447 1524
rect 1404 1393 1405 1526
rect 1486 1393 1487 1526
rect 1383 1393 1384 1528
rect 1404 1527 1405 1536
rect 1407 1527 1408 1536
rect 1473 1393 1474 1528
rect 1437 1393 1438 1530
rect 1458 1393 1459 1530
rect 1455 1393 1456 1532
rect 1507 1393 1508 1532
rect 1470 1393 1471 1534
rect 1479 1393 1480 1534
rect 997 1540 998 1543
rect 1066 1540 1067 1543
rect 1016 1540 1017 1545
rect 1081 1540 1082 1545
rect 1024 1546 1025 1669
rect 1108 1546 1109 1669
rect 1031 1548 1032 1669
rect 1038 1540 1039 1549
rect 1035 1540 1036 1551
rect 1053 1540 1054 1551
rect 1026 1540 1027 1553
rect 1034 1552 1035 1669
rect 1027 1554 1028 1669
rect 1075 1540 1076 1555
rect 1041 1540 1042 1557
rect 1175 1540 1176 1557
rect 1043 1558 1044 1669
rect 1127 1540 1128 1559
rect 1052 1560 1053 1669
rect 1241 1540 1242 1561
rect 1057 1540 1058 1563
rect 1148 1540 1149 1563
rect 1056 1564 1057 1669
rect 1154 1540 1155 1565
rect 1063 1540 1064 1567
rect 1080 1566 1081 1669
rect 1068 1568 1069 1669
rect 1087 1540 1088 1569
rect 1086 1570 1087 1669
rect 1118 1540 1119 1571
rect 1019 1540 1020 1573
rect 1117 1572 1118 1669
rect 1020 1574 1021 1669
rect 1150 1574 1151 1669
rect 1100 1540 1101 1577
rect 1226 1540 1227 1577
rect 1102 1578 1103 1669
rect 1240 1578 1241 1669
rect 1120 1580 1121 1669
rect 1121 1540 1122 1581
rect 1124 1540 1125 1581
rect 1147 1580 1148 1669
rect 1136 1540 1137 1583
rect 1153 1582 1154 1669
rect 1160 1540 1161 1583
rect 1183 1582 1184 1669
rect 1012 1540 1013 1585
rect 1159 1584 1160 1669
rect 1169 1540 1170 1585
rect 1198 1584 1199 1669
rect 1145 1540 1146 1587
rect 1168 1586 1169 1669
rect 1172 1540 1173 1587
rect 1204 1586 1205 1669
rect 1060 1540 1061 1589
rect 1171 1588 1172 1669
rect 1059 1590 1060 1669
rect 1135 1590 1136 1669
rect 1177 1590 1178 1669
rect 1304 1540 1305 1591
rect 1187 1540 1188 1593
rect 1246 1592 1247 1669
rect 1186 1594 1187 1669
rect 1190 1540 1191 1595
rect 1074 1596 1075 1669
rect 1189 1596 1190 1669
rect 1196 1540 1197 1597
rect 1207 1596 1208 1669
rect 1166 1540 1167 1599
rect 1195 1598 1196 1669
rect 1142 1540 1143 1601
rect 1165 1600 1166 1669
rect 1201 1600 1202 1669
rect 1223 1540 1224 1601
rect 1050 1540 1051 1603
rect 1222 1602 1223 1669
rect 1217 1540 1218 1605
rect 1231 1604 1232 1669
rect 1220 1540 1221 1607
rect 1237 1606 1238 1669
rect 1193 1540 1194 1609
rect 1219 1608 1220 1669
rect 1225 1608 1226 1669
rect 1253 1540 1254 1609
rect 1229 1540 1230 1611
rect 1252 1610 1253 1669
rect 1228 1612 1229 1669
rect 1256 1540 1257 1613
rect 1235 1540 1236 1615
rect 1336 1614 1337 1669
rect 1249 1616 1250 1669
rect 1259 1540 1260 1617
rect 1262 1540 1263 1617
rect 1312 1616 1313 1669
rect 1265 1540 1266 1619
rect 1300 1618 1301 1669
rect 1243 1620 1244 1669
rect 1264 1620 1265 1669
rect 1283 1540 1284 1621
rect 1318 1620 1319 1669
rect 1286 1540 1287 1623
rect 1294 1622 1295 1669
rect 1310 1540 1311 1623
rect 1385 1540 1386 1623
rect 1316 1540 1317 1625
rect 1334 1540 1335 1625
rect 1315 1626 1316 1669
rect 1418 1540 1419 1627
rect 1333 1628 1334 1669
rect 1376 1540 1377 1629
rect 1346 1540 1347 1631
rect 1384 1630 1385 1669
rect 1345 1632 1346 1669
rect 1355 1540 1356 1633
rect 1349 1540 1350 1635
rect 1415 1634 1416 1669
rect 1348 1636 1349 1669
rect 1358 1540 1359 1637
rect 1352 1540 1353 1639
rect 1381 1638 1382 1669
rect 1340 1540 1341 1641
rect 1351 1640 1352 1669
rect 1339 1642 1340 1669
rect 1373 1540 1374 1643
rect 1331 1540 1332 1645
rect 1372 1644 1373 1669
rect 1354 1646 1355 1669
rect 1379 1540 1380 1647
rect 1367 1540 1368 1649
rect 1396 1648 1397 1669
rect 1370 1540 1371 1651
rect 1400 1540 1401 1651
rect 1328 1540 1329 1653
rect 1369 1652 1370 1669
rect 1327 1654 1328 1669
rect 1421 1540 1422 1655
rect 1388 1540 1389 1657
rect 1405 1656 1406 1669
rect 1387 1658 1388 1669
rect 1425 1658 1426 1669
rect 1391 1540 1392 1661
rect 1399 1660 1400 1669
rect 1270 1662 1271 1669
rect 1390 1662 1391 1669
rect 1394 1540 1395 1663
rect 1402 1662 1403 1669
rect 1288 1664 1289 1669
rect 1393 1664 1394 1669
rect 1407 1540 1408 1665
rect 1422 1664 1423 1669
rect 1342 1666 1343 1669
rect 1408 1666 1409 1669
rect 1006 1673 1007 1676
rect 1195 1673 1196 1676
rect 1010 1673 1011 1678
rect 1043 1673 1044 1678
rect 1013 1673 1014 1680
rect 1150 1673 1151 1680
rect 1003 1673 1004 1682
rect 1151 1681 1152 1822
rect 1017 1673 1018 1684
rect 1049 1673 1050 1684
rect 1020 1673 1021 1686
rect 1034 1673 1035 1686
rect 1009 1687 1010 1822
rect 1019 1687 1020 1822
rect 1024 1673 1025 1688
rect 1100 1687 1101 1822
rect 1030 1689 1031 1822
rect 1204 1673 1205 1690
rect 1037 1691 1038 1822
rect 1168 1673 1169 1692
rect 1059 1673 1060 1694
rect 1068 1673 1069 1694
rect 1059 1695 1060 1822
rect 1177 1673 1178 1696
rect 1062 1697 1063 1822
rect 1080 1673 1081 1698
rect 1068 1699 1069 1822
rect 1196 1699 1197 1822
rect 1077 1673 1078 1702
rect 1178 1701 1179 1822
rect 1079 1703 1080 1822
rect 1189 1673 1190 1704
rect 1083 1673 1084 1706
rect 1120 1673 1121 1706
rect 1082 1707 1083 1822
rect 1237 1673 1238 1708
rect 1097 1709 1098 1822
rect 1108 1673 1109 1710
rect 1102 1673 1103 1712
rect 1231 1673 1232 1712
rect 1105 1673 1106 1714
rect 1307 1713 1308 1822
rect 1106 1715 1107 1822
rect 1228 1673 1229 1716
rect 1115 1717 1116 1822
rect 1117 1673 1118 1718
rect 1118 1719 1119 1822
rect 1198 1673 1199 1720
rect 1127 1721 1128 1822
rect 1135 1673 1136 1722
rect 1133 1723 1134 1822
rect 1153 1673 1154 1724
rect 1139 1725 1140 1822
rect 1147 1673 1148 1726
rect 1142 1727 1143 1822
rect 1159 1673 1160 1728
rect 1056 1673 1057 1730
rect 1160 1729 1161 1822
rect 1148 1731 1149 1822
rect 1165 1673 1166 1732
rect 1154 1733 1155 1822
rect 1171 1673 1172 1734
rect 1172 1735 1173 1822
rect 1183 1673 1184 1736
rect 1175 1737 1176 1822
rect 1186 1673 1187 1738
rect 1184 1739 1185 1822
rect 1207 1673 1208 1740
rect 1187 1741 1188 1822
rect 1222 1673 1223 1742
rect 1199 1743 1200 1822
rect 1201 1673 1202 1744
rect 1202 1745 1203 1822
rect 1225 1673 1226 1746
rect 1205 1747 1206 1822
rect 1363 1673 1364 1748
rect 1208 1749 1209 1822
rect 1246 1673 1247 1750
rect 1211 1751 1212 1822
rect 1240 1673 1241 1752
rect 1219 1673 1220 1754
rect 1235 1753 1236 1822
rect 1220 1755 1221 1822
rect 1249 1673 1250 1756
rect 1229 1757 1230 1822
rect 1336 1673 1337 1758
rect 1232 1759 1233 1822
rect 1252 1673 1253 1760
rect 1265 1759 1266 1822
rect 1345 1673 1346 1760
rect 1267 1673 1268 1762
rect 1270 1673 1271 1762
rect 1268 1763 1269 1822
rect 1298 1763 1299 1822
rect 1283 1765 1284 1822
rect 1318 1673 1319 1766
rect 1288 1673 1289 1768
rect 1292 1767 1293 1822
rect 1289 1769 1290 1822
rect 1339 1673 1340 1770
rect 1294 1673 1295 1772
rect 1304 1771 1305 1822
rect 1295 1773 1296 1822
rect 1322 1773 1323 1822
rect 1300 1673 1301 1776
rect 1390 1673 1391 1776
rect 1301 1777 1302 1822
rect 1402 1673 1403 1778
rect 1310 1779 1311 1822
rect 1312 1673 1313 1780
rect 1313 1781 1314 1822
rect 1422 1673 1423 1782
rect 1315 1673 1316 1784
rect 1325 1783 1326 1822
rect 1316 1785 1317 1822
rect 1369 1673 1370 1786
rect 1319 1787 1320 1822
rect 1372 1673 1373 1788
rect 1327 1673 1328 1790
rect 1418 1673 1419 1790
rect 1328 1791 1329 1822
rect 1405 1673 1406 1792
rect 1331 1793 1332 1822
rect 1428 1673 1429 1794
rect 1333 1673 1334 1796
rect 1354 1673 1355 1796
rect 1337 1797 1338 1822
rect 1381 1673 1382 1798
rect 1334 1799 1335 1822
rect 1381 1799 1382 1822
rect 1342 1673 1343 1802
rect 1393 1673 1394 1802
rect 1348 1673 1349 1804
rect 1366 1673 1367 1804
rect 1347 1805 1348 1822
rect 1399 1673 1400 1806
rect 1354 1807 1355 1822
rect 1387 1673 1388 1808
rect 1360 1809 1361 1822
rect 1403 1809 1404 1822
rect 1363 1811 1364 1822
rect 1388 1811 1389 1822
rect 1375 1813 1376 1822
rect 1435 1673 1436 1814
rect 1378 1815 1379 1822
rect 1442 1673 1443 1816
rect 1384 1673 1385 1818
rect 1425 1673 1426 1818
rect 1396 1673 1397 1820
rect 1438 1673 1439 1820
rect 1012 1826 1013 1829
rect 1139 1826 1140 1829
rect 1012 1830 1013 1937
rect 1019 1830 1020 1937
rect 1016 1826 1017 1833
rect 1120 1832 1121 1937
rect 1023 1834 1024 1937
rect 1030 1834 1031 1937
rect 1033 1826 1034 1835
rect 1189 1834 1190 1937
rect 1040 1826 1041 1837
rect 1129 1836 1130 1937
rect 1044 1826 1045 1839
rect 1133 1826 1134 1839
rect 1047 1826 1048 1841
rect 1127 1826 1128 1841
rect 1056 1826 1057 1843
rect 1144 1842 1145 1937
rect 1059 1826 1060 1845
rect 1187 1826 1188 1845
rect 1060 1846 1061 1937
rect 1062 1826 1063 1847
rect 1063 1848 1064 1937
rect 1160 1826 1161 1849
rect 1065 1826 1066 1851
rect 1175 1826 1176 1851
rect 1066 1852 1067 1937
rect 1213 1852 1214 1937
rect 1070 1854 1071 1937
rect 1304 1826 1305 1855
rect 1080 1856 1081 1937
rect 1301 1826 1302 1857
rect 1084 1858 1085 1937
rect 1208 1826 1209 1859
rect 1103 1826 1104 1861
rect 1126 1860 1127 1937
rect 1097 1826 1098 1863
rect 1102 1862 1103 1937
rect 1096 1864 1097 1937
rect 1100 1826 1101 1865
rect 1114 1864 1115 1937
rect 1115 1826 1116 1865
rect 1117 1864 1118 1937
rect 1118 1826 1119 1865
rect 1151 1826 1152 1865
rect 1156 1864 1157 1937
rect 1154 1826 1155 1867
rect 1174 1866 1175 1937
rect 1148 1826 1149 1869
rect 1153 1868 1154 1937
rect 1142 1826 1143 1871
rect 1147 1870 1148 1937
rect 1026 1826 1027 1873
rect 1141 1872 1142 1937
rect 1165 1872 1166 1937
rect 1202 1826 1203 1873
rect 1171 1874 1172 1937
rect 1172 1826 1173 1875
rect 1184 1826 1185 1875
rect 1192 1874 1193 1937
rect 1183 1876 1184 1937
rect 1207 1876 1208 1937
rect 1205 1826 1206 1879
rect 1222 1878 1223 1937
rect 1217 1826 1218 1881
rect 1232 1826 1233 1881
rect 1211 1826 1212 1883
rect 1216 1882 1217 1937
rect 1210 1884 1211 1937
rect 1220 1826 1221 1885
rect 1123 1886 1124 1937
rect 1219 1886 1220 1937
rect 1229 1826 1230 1887
rect 1235 1826 1236 1887
rect 1228 1888 1229 1937
rect 1240 1888 1241 1937
rect 1237 1890 1238 1937
rect 1238 1826 1239 1891
rect 1249 1890 1250 1937
rect 1295 1826 1296 1891
rect 1252 1892 1253 1937
rect 1268 1826 1269 1893
rect 1255 1894 1256 1937
rect 1289 1826 1290 1895
rect 1265 1826 1266 1897
rect 1298 1826 1299 1897
rect 1264 1898 1265 1937
rect 1279 1898 1280 1937
rect 1273 1900 1274 1937
rect 1313 1826 1314 1901
rect 1276 1902 1277 1937
rect 1307 1826 1308 1903
rect 1288 1904 1289 1937
rect 1328 1826 1329 1905
rect 1292 1826 1293 1907
rect 1340 1826 1341 1907
rect 1291 1908 1292 1937
rect 1331 1826 1332 1909
rect 1294 1910 1295 1937
rect 1357 1910 1358 1937
rect 1297 1912 1298 1937
rect 1331 1912 1332 1937
rect 1303 1914 1304 1937
rect 1319 1826 1320 1915
rect 1310 1826 1311 1917
rect 1325 1826 1326 1917
rect 1199 1826 1200 1919
rect 1324 1918 1325 1937
rect 1196 1826 1197 1921
rect 1198 1920 1199 1937
rect 1178 1826 1179 1923
rect 1195 1922 1196 1937
rect 1314 1922 1315 1937
rect 1316 1826 1317 1923
rect 1334 1826 1335 1923
rect 1340 1922 1341 1937
rect 1334 1924 1335 1937
rect 1363 1826 1364 1925
rect 1337 1826 1338 1927
rect 1403 1826 1404 1927
rect 1283 1826 1284 1929
rect 1337 1928 1338 1937
rect 1347 1928 1348 1937
rect 1381 1826 1382 1929
rect 1364 1930 1365 1937
rect 1397 1826 1398 1931
rect 1375 1826 1376 1933
rect 1391 1826 1392 1933
rect 1360 1826 1361 1935
rect 1374 1934 1375 1937
rect 1378 1826 1379 1935
rect 1388 1826 1389 1935
rect 997 1943 998 2048
rect 1009 1943 1010 2048
rect 1019 1941 1020 1944
rect 1174 1941 1175 1944
rect 1012 1945 1013 2048
rect 1019 1945 1020 2048
rect 1023 1941 1024 1946
rect 1099 1945 1100 2048
rect 1023 1947 1024 2048
rect 1120 1941 1121 1948
rect 1030 1941 1031 1950
rect 1141 1941 1142 1950
rect 1033 1941 1034 1952
rect 1129 1941 1130 1952
rect 1035 1953 1036 2048
rect 1060 1941 1061 1954
rect 1052 1955 1053 2048
rect 1096 1941 1097 1956
rect 1057 1941 1058 1958
rect 1162 1957 1163 2048
rect 1059 1959 1060 2048
rect 1192 1941 1193 1960
rect 1066 1941 1067 1962
rect 1132 1961 1133 2048
rect 1087 1941 1088 1964
rect 1213 1941 1214 1964
rect 1090 1965 1091 2048
rect 1102 1941 1103 1966
rect 1093 1967 1094 2048
rect 1144 1941 1145 1968
rect 1096 1969 1097 2048
rect 1117 1941 1118 1970
rect 1102 1971 1103 2048
rect 1198 1941 1199 1972
rect 1105 1973 1106 2048
rect 1159 1973 1160 2048
rect 1114 1941 1115 1976
rect 1174 1975 1175 2048
rect 1120 1977 1121 2048
rect 1147 1941 1148 1978
rect 1126 1979 1127 2048
rect 1153 1941 1154 1980
rect 1129 1981 1130 2048
rect 1156 1941 1157 1982
rect 1141 1983 1142 2048
rect 1216 1941 1217 1984
rect 1150 1985 1151 2048
rect 1171 1941 1172 1986
rect 1070 1941 1071 1988
rect 1171 1987 1172 2048
rect 1063 1941 1064 1990
rect 1069 1989 1070 2048
rect 1153 1989 1154 2048
rect 1195 1941 1196 1990
rect 1156 1991 1157 2048
rect 1189 1941 1190 1992
rect 1183 1941 1184 1994
rect 1210 1941 1211 1994
rect 1183 1995 1184 2048
rect 1207 1941 1208 1996
rect 1186 1995 1187 2048
rect 1186 1941 1187 1996
rect 1195 1997 1196 2048
rect 1219 1941 1220 1998
rect 1084 1941 1085 2000
rect 1219 1999 1220 2048
rect 1045 1941 1046 2002
rect 1084 2001 1085 2048
rect 1198 2001 1199 2048
rect 1222 1941 1223 2002
rect 1165 1941 1166 2004
rect 1222 2003 1223 2048
rect 1073 1941 1074 2006
rect 1165 2005 1166 2048
rect 1201 2005 1202 2048
rect 1240 1941 1241 2006
rect 1204 2007 1205 2048
rect 1241 2007 1242 2048
rect 1213 2009 1214 2048
rect 1258 1941 1259 2010
rect 1228 1941 1229 2012
rect 1249 1941 1250 2012
rect 1232 2013 1233 2048
rect 1255 1941 1256 2014
rect 1237 1941 1238 2016
rect 1317 2015 1318 2048
rect 1247 2017 1248 2048
rect 1291 1941 1292 2018
rect 1252 1941 1253 2020
rect 1256 2019 1257 2048
rect 1229 2021 1230 2048
rect 1253 2021 1254 2048
rect 1259 2021 1260 2048
rect 1261 1941 1262 2022
rect 1226 2023 1227 2048
rect 1262 2023 1263 2048
rect 1273 1941 1274 2024
rect 1274 2023 1275 2048
rect 1279 1941 1280 2024
rect 1292 2023 1293 2048
rect 1264 1941 1265 2026
rect 1280 2025 1281 2048
rect 1288 1941 1289 2026
rect 1304 2025 1305 2048
rect 1294 1941 1295 2028
rect 1361 1941 1362 2028
rect 1276 1941 1277 2030
rect 1295 2029 1296 2048
rect 1277 2031 1278 2048
rect 1314 1941 1315 2032
rect 1297 1941 1298 2034
rect 1301 2033 1302 2048
rect 1298 2035 1299 2048
rect 1357 1941 1358 2036
rect 1307 1941 1308 2038
rect 1337 1941 1338 2038
rect 1323 2039 1324 2048
rect 1353 2039 1354 2048
rect 1328 1941 1329 2042
rect 1340 1941 1341 2042
rect 1334 1941 1335 2044
rect 1343 1941 1344 2044
rect 1307 2045 1308 2048
rect 1343 2045 1344 2048
rect 1367 1941 1368 2046
rect 1377 1941 1378 2046
rect 1000 2052 1001 2055
rect 1035 2052 1036 2055
rect 1016 2052 1017 2057
rect 1096 2052 1097 2057
rect 1026 2052 1027 2059
rect 1066 2058 1067 2129
rect 1034 2060 1035 2129
rect 1093 2052 1094 2061
rect 1041 2052 1042 2063
rect 1079 2062 1080 2129
rect 1043 2064 1044 2129
rect 1156 2052 1157 2065
rect 1045 2052 1046 2067
rect 1142 2066 1143 2129
rect 1048 2052 1049 2069
rect 1084 2052 1085 2069
rect 1050 2070 1051 2129
rect 1129 2052 1130 2071
rect 1052 2052 1053 2073
rect 1171 2052 1172 2073
rect 1059 2052 1060 2075
rect 1106 2074 1107 2129
rect 1082 2076 1083 2129
rect 1145 2076 1146 2129
rect 1085 2078 1086 2129
rect 1109 2078 1110 2129
rect 1094 2080 1095 2129
rect 1099 2052 1100 2081
rect 1102 2052 1103 2081
rect 1229 2052 1230 2081
rect 1090 2052 1091 2083
rect 1103 2082 1104 2129
rect 1126 2052 1127 2083
rect 1139 2082 1140 2129
rect 1073 2084 1074 2129
rect 1127 2084 1128 2129
rect 1150 2052 1151 2085
rect 1157 2084 1158 2129
rect 1162 2052 1163 2085
rect 1169 2084 1170 2129
rect 1055 2052 1056 2087
rect 1163 2086 1164 2129
rect 1165 2052 1166 2087
rect 1172 2086 1173 2129
rect 1159 2052 1160 2089
rect 1166 2088 1167 2129
rect 1153 2052 1154 2091
rect 1160 2090 1161 2129
rect 1174 2052 1175 2091
rect 1175 2090 1176 2129
rect 1178 2090 1179 2129
rect 1280 2052 1281 2091
rect 1183 2052 1184 2093
rect 1226 2052 1227 2093
rect 1195 2052 1196 2095
rect 1196 2094 1197 2129
rect 1198 2052 1199 2095
rect 1222 2052 1223 2095
rect 1201 2052 1202 2097
rect 1223 2096 1224 2129
rect 1186 2052 1187 2099
rect 1202 2098 1203 2129
rect 1204 2052 1205 2099
rect 1226 2098 1227 2129
rect 1205 2100 1206 2129
rect 1250 2100 1251 2129
rect 1232 2052 1233 2103
rect 1235 2102 1236 2129
rect 1190 2104 1191 2129
rect 1232 2104 1233 2129
rect 1244 2052 1245 2105
rect 1310 2104 1311 2129
rect 1244 2106 1245 2129
rect 1247 2052 1248 2107
rect 1253 2052 1254 2107
rect 1268 2106 1269 2129
rect 1256 2106 1257 2129
rect 1256 2052 1257 2107
rect 1259 2106 1260 2129
rect 1259 2052 1260 2107
rect 1271 2106 1272 2129
rect 1332 2106 1333 2129
rect 1274 2052 1275 2109
rect 1343 2052 1344 2109
rect 1277 2052 1278 2111
rect 1325 2110 1326 2129
rect 1199 2112 1200 2129
rect 1277 2112 1278 2129
rect 1286 2112 1287 2129
rect 1307 2052 1308 2113
rect 1213 2052 1214 2115
rect 1307 2114 1308 2129
rect 1298 2052 1299 2117
rect 1356 2052 1357 2117
rect 1292 2052 1293 2119
rect 1298 2118 1299 2129
rect 1301 2052 1302 2119
rect 1313 2118 1314 2129
rect 1295 2052 1296 2121
rect 1301 2120 1302 2129
rect 1304 2052 1305 2121
rect 1316 2120 1317 2129
rect 1319 2120 1320 2129
rect 1340 2052 1341 2121
rect 1304 2122 1305 2129
rect 1339 2122 1340 2129
rect 1323 2052 1324 2125
rect 1346 2052 1347 2125
rect 1238 2126 1239 2129
rect 1346 2126 1347 2129
rect 1015 2133 1016 2136
rect 1094 2133 1095 2136
rect 1022 2133 1023 2138
rect 1079 2133 1080 2138
rect 1025 2133 1026 2140
rect 1103 2133 1104 2140
rect 1024 2141 1025 2236
rect 1034 2133 1035 2142
rect 1031 2143 1032 2236
rect 1040 2133 1041 2144
rect 1034 2145 1035 2236
rect 1106 2133 1107 2146
rect 1037 2147 1038 2236
rect 1139 2133 1140 2148
rect 1040 2149 1041 2236
rect 1133 2133 1134 2150
rect 1044 2151 1045 2236
rect 1157 2133 1158 2152
rect 1047 2133 1048 2154
rect 1089 2153 1090 2236
rect 1062 2133 1063 2156
rect 1095 2155 1096 2236
rect 1066 2133 1067 2158
rect 1163 2133 1164 2158
rect 1065 2159 1066 2236
rect 1131 2159 1132 2236
rect 1069 2133 1070 2162
rect 1098 2161 1099 2236
rect 1056 2163 1057 2236
rect 1069 2163 1070 2236
rect 1073 2133 1074 2164
rect 1121 2133 1122 2164
rect 1079 2165 1080 2236
rect 1212 2165 1213 2236
rect 1085 2133 1086 2168
rect 1169 2133 1170 2168
rect 1092 2169 1093 2236
rect 1142 2133 1143 2170
rect 1107 2171 1108 2236
rect 1127 2133 1128 2172
rect 1109 2133 1110 2174
rect 1140 2173 1141 2236
rect 1119 2175 1120 2236
rect 1166 2133 1167 2176
rect 1125 2177 1126 2236
rect 1172 2133 1173 2178
rect 1128 2179 1129 2236
rect 1175 2133 1176 2180
rect 1137 2181 1138 2236
rect 1145 2133 1146 2182
rect 1149 2181 1150 2236
rect 1196 2133 1197 2182
rect 1154 2133 1155 2184
rect 1215 2183 1216 2236
rect 1160 2133 1161 2186
rect 1253 2133 1254 2186
rect 1164 2187 1165 2236
rect 1199 2133 1200 2188
rect 1170 2189 1171 2236
rect 1205 2133 1206 2190
rect 1176 2191 1177 2236
rect 1202 2133 1203 2192
rect 1179 2193 1180 2236
rect 1190 2133 1191 2194
rect 1188 2195 1189 2236
rect 1226 2133 1227 2196
rect 1191 2197 1192 2236
rect 1223 2133 1224 2198
rect 1200 2199 1201 2236
rect 1350 2133 1351 2200
rect 1221 2201 1222 2236
rect 1298 2133 1299 2202
rect 1225 2203 1226 2236
rect 1265 2203 1266 2236
rect 1231 2205 1232 2236
rect 1271 2133 1272 2206
rect 1241 2207 1242 2236
rect 1250 2207 1251 2236
rect 1244 2133 1245 2210
rect 1274 2209 1275 2236
rect 1247 2211 1248 2236
rect 1301 2133 1302 2212
rect 1256 2133 1257 2214
rect 1310 2133 1311 2214
rect 1259 2133 1260 2216
rect 1322 2133 1323 2216
rect 1259 2217 1260 2236
rect 1280 2217 1281 2236
rect 1262 2219 1263 2236
rect 1304 2133 1305 2220
rect 1268 2133 1269 2222
rect 1329 2133 1330 2222
rect 1235 2133 1236 2224
rect 1268 2223 1269 2236
rect 1152 2225 1153 2236
rect 1234 2225 1235 2236
rect 1271 2225 1272 2236
rect 1316 2133 1317 2226
rect 1286 2133 1287 2228
rect 1339 2133 1340 2228
rect 1238 2133 1239 2230
rect 1287 2229 1288 2236
rect 1313 2133 1314 2230
rect 1343 2133 1344 2230
rect 1319 2133 1320 2232
rect 1346 2133 1347 2232
rect 1332 2133 1333 2234
rect 1336 2133 1337 2234
rect 1021 2240 1022 2243
rect 1034 2240 1035 2243
rect 1037 2242 1038 2301
rect 1056 2240 1057 2243
rect 1044 2240 1045 2245
rect 1095 2240 1096 2245
rect 1044 2246 1045 2301
rect 1047 2240 1048 2247
rect 1051 2246 1052 2301
rect 1271 2240 1272 2247
rect 1062 2240 1063 2249
rect 1066 2248 1067 2301
rect 1069 2240 1070 2249
rect 1128 2240 1129 2249
rect 1073 2250 1074 2301
rect 1083 2240 1084 2251
rect 1086 2240 1087 2251
rect 1188 2240 1189 2251
rect 1086 2252 1087 2301
rect 1089 2240 1090 2253
rect 1089 2254 1090 2301
rect 1092 2240 1093 2255
rect 1028 2240 1029 2257
rect 1092 2256 1093 2301
rect 1027 2258 1028 2301
rect 1137 2240 1138 2259
rect 1095 2260 1096 2301
rect 1098 2240 1099 2261
rect 1079 2240 1080 2263
rect 1098 2262 1099 2301
rect 1122 2262 1123 2301
rect 1212 2240 1213 2263
rect 1131 2240 1132 2265
rect 1155 2264 1156 2301
rect 1140 2240 1141 2267
rect 1158 2266 1159 2301
rect 1143 2268 1144 2301
rect 1179 2240 1180 2269
rect 1149 2240 1150 2271
rect 1173 2270 1174 2301
rect 1125 2240 1126 2273
rect 1149 2272 1150 2301
rect 1119 2240 1120 2275
rect 1125 2274 1126 2301
rect 1080 2276 1081 2301
rect 1119 2276 1120 2301
rect 1152 2240 1153 2277
rect 1225 2240 1226 2277
rect 1107 2240 1108 2279
rect 1152 2278 1153 2301
rect 1161 2278 1162 2301
rect 1164 2240 1165 2279
rect 1170 2240 1171 2279
rect 1204 2278 1205 2301
rect 1170 2280 1171 2301
rect 1176 2240 1177 2281
rect 1176 2282 1177 2301
rect 1226 2282 1227 2301
rect 1182 2284 1183 2301
rect 1215 2240 1216 2285
rect 1191 2284 1192 2301
rect 1191 2240 1192 2285
rect 1194 2286 1195 2301
rect 1207 2286 1208 2301
rect 1200 2240 1201 2289
rect 1284 2240 1285 2289
rect 1167 2290 1168 2301
rect 1200 2290 1201 2301
rect 1210 2290 1211 2301
rect 1247 2240 1248 2291
rect 1213 2292 1214 2301
rect 1231 2240 1232 2293
rect 1223 2294 1224 2301
rect 1250 2240 1251 2295
rect 1259 2240 1260 2295
rect 1277 2240 1278 2295
rect 1262 2240 1263 2297
rect 1280 2240 1281 2297
rect 1274 2240 1275 2299
rect 1287 2240 1288 2299
rect 1027 2305 1028 2308
rect 1149 2305 1150 2308
rect 1037 2305 1038 2310
rect 1089 2305 1090 2310
rect 1041 2311 1042 2364
rect 1092 2305 1093 2312
rect 1027 2313 1028 2364
rect 1092 2313 1093 2364
rect 1044 2305 1045 2316
rect 1125 2305 1126 2316
rect 1051 2305 1052 2318
rect 1073 2305 1074 2318
rect 1034 2305 1035 2320
rect 1074 2319 1075 2364
rect 1034 2321 1035 2364
rect 1152 2305 1153 2322
rect 1056 2323 1057 2364
rect 1076 2305 1077 2324
rect 1044 2325 1045 2364
rect 1077 2325 1078 2364
rect 1071 2327 1072 2364
rect 1086 2305 1087 2328
rect 1080 2329 1081 2364
rect 1095 2305 1096 2330
rect 1089 2331 1090 2364
rect 1113 2331 1114 2364
rect 1095 2333 1096 2364
rect 1098 2305 1099 2334
rect 1104 2333 1105 2364
rect 1155 2305 1156 2334
rect 1110 2335 1111 2364
rect 1158 2305 1159 2336
rect 1116 2337 1117 2364
rect 1179 2305 1180 2338
rect 1119 2305 1120 2340
rect 1164 2339 1165 2364
rect 1134 2341 1135 2364
rect 1167 2305 1168 2342
rect 1143 2305 1144 2344
rect 1155 2343 1156 2364
rect 1152 2345 1153 2364
rect 1170 2305 1171 2346
rect 1158 2347 1159 2364
rect 1191 2305 1192 2348
rect 1161 2305 1162 2350
rect 1197 2305 1198 2350
rect 1122 2305 1123 2352
rect 1161 2351 1162 2364
rect 1122 2353 1123 2364
rect 1170 2353 1171 2364
rect 1173 2305 1174 2354
rect 1182 2305 1183 2354
rect 1173 2355 1174 2364
rect 1176 2305 1177 2356
rect 1176 2357 1177 2364
rect 1182 2357 1183 2364
rect 1185 2357 1186 2364
rect 1213 2305 1214 2358
rect 1194 2305 1195 2360
rect 1195 2359 1196 2364
rect 1200 2305 1201 2360
rect 1210 2305 1211 2360
rect 1204 2305 1205 2362
rect 1216 2305 1217 2362
rect 1232 2305 1233 2362
rect 1239 2305 1240 2362
rect 1245 2305 1246 2362
rect 1252 2305 1253 2362
rect 1030 2368 1031 2371
rect 1083 2370 1084 2409
rect 1033 2372 1034 2409
rect 1074 2368 1075 2373
rect 1041 2368 1042 2375
rect 1062 2374 1063 2409
rect 1050 2376 1051 2409
rect 1071 2368 1072 2377
rect 1053 2368 1054 2379
rect 1095 2368 1096 2379
rect 1040 2380 1041 2409
rect 1095 2380 1096 2409
rect 1059 2382 1060 2409
rect 1077 2368 1078 2383
rect 1065 2368 1066 2385
rect 1155 2368 1156 2385
rect 1068 2368 1069 2387
rect 1089 2386 1090 2409
rect 1080 2368 1081 2389
rect 1086 2368 1087 2389
rect 1037 2368 1038 2391
rect 1086 2390 1087 2409
rect 1036 2392 1037 2409
rect 1077 2392 1078 2409
rect 1092 2368 1093 2393
rect 1101 2392 1102 2409
rect 1110 2368 1111 2393
rect 1188 2368 1189 2393
rect 1116 2368 1117 2395
rect 1149 2394 1150 2409
rect 1113 2368 1114 2397
rect 1116 2396 1117 2409
rect 1104 2368 1105 2399
rect 1113 2398 1114 2409
rect 1056 2368 1057 2401
rect 1104 2400 1105 2409
rect 1122 2368 1123 2401
rect 1125 2400 1126 2409
rect 1128 2400 1129 2409
rect 1134 2368 1135 2401
rect 1137 2400 1138 2409
rect 1173 2368 1174 2401
rect 1140 2402 1141 2409
rect 1158 2368 1159 2403
rect 1152 2402 1153 2409
rect 1152 2368 1153 2403
rect 1161 2368 1162 2403
rect 1170 2368 1171 2403
rect 1164 2368 1165 2405
rect 1167 2368 1168 2405
rect 1176 2368 1177 2405
rect 1191 2368 1192 2405
rect 1182 2368 1183 2407
rect 1185 2368 1186 2407
rect 1033 2413 1034 2416
rect 1083 2413 1084 2416
rect 1040 2413 1041 2418
rect 1062 2413 1063 2418
rect 1039 2419 1040 2450
rect 1059 2413 1060 2420
rect 1042 2421 1043 2450
rect 1089 2413 1090 2422
rect 1045 2423 1046 2450
rect 1077 2413 1078 2424
rect 1047 2413 1048 2426
rect 1104 2413 1105 2426
rect 1048 2427 1049 2450
rect 1054 2427 1055 2450
rect 1050 2413 1051 2430
rect 1101 2413 1102 2430
rect 1058 2431 1059 2450
rect 1113 2413 1114 2432
rect 1065 2433 1066 2450
rect 1116 2413 1117 2434
rect 1072 2435 1073 2450
rect 1137 2413 1138 2436
rect 1078 2437 1079 2450
rect 1128 2413 1129 2438
rect 1086 2413 1087 2440
rect 1119 2413 1120 2440
rect 1098 2413 1099 2442
rect 1131 2413 1132 2442
rect 1122 2413 1123 2444
rect 1140 2413 1141 2444
rect 1125 2413 1126 2446
rect 1146 2413 1147 2446
rect 1143 2413 1144 2448
rect 1149 2413 1150 2448
rect 1039 2454 1040 2457
rect 1061 2454 1062 2457
rect 1045 2454 1046 2459
rect 1048 2454 1049 2459
rect 1054 2454 1055 2459
rect 1072 2454 1073 2459
rect 1058 2454 1059 2461
rect 1078 2454 1079 2461
<< via >>
rect 1028 497 1029 498
rect 1047 497 1048 498
rect 1038 499 1039 500
rect 1068 499 1069 500
rect 1041 501 1042 502
rect 1062 501 1063 502
rect 1050 503 1051 504
rect 1071 503 1072 504
rect 1074 503 1075 504
rect 1077 503 1078 504
rect 1084 503 1085 504
rect 1090 503 1091 504
rect 1099 503 1100 504
rect 1102 503 1103 504
rect 1132 503 1133 504
rect 1139 503 1140 504
rect 1021 513 1022 514
rect 1034 513 1035 514
rect 1031 515 1032 516
rect 1056 515 1057 516
rect 1044 517 1045 518
rect 1068 517 1069 518
rect 1047 519 1048 520
rect 1068 519 1069 520
rect 1046 521 1047 522
rect 1071 521 1072 522
rect 1050 523 1051 524
rect 1062 523 1063 524
rect 1028 525 1029 526
rect 1062 525 1063 526
rect 1053 527 1054 528
rect 1074 527 1075 528
rect 1028 529 1029 530
rect 1074 529 1075 530
rect 1031 531 1032 532
rect 1053 531 1054 532
rect 1077 531 1078 532
rect 1157 531 1158 532
rect 1021 533 1022 534
rect 1077 533 1078 534
rect 1080 533 1081 534
rect 1127 533 1128 534
rect 1087 535 1088 536
rect 1170 535 1171 536
rect 1090 537 1091 538
rect 1130 537 1131 538
rect 1090 539 1091 540
rect 1102 539 1103 540
rect 1093 541 1094 542
rect 1154 541 1155 542
rect 1099 543 1100 544
rect 1182 543 1183 544
rect 1087 545 1088 546
rect 1099 545 1100 546
rect 1105 545 1106 546
rect 1226 545 1227 546
rect 1112 547 1113 548
rect 1124 547 1125 548
rect 1115 549 1116 550
rect 1145 549 1146 550
rect 1142 551 1143 552
rect 1151 551 1152 552
rect 1164 551 1165 552
rect 1197 551 1198 552
rect 1167 553 1168 554
rect 1188 553 1189 554
rect 1200 553 1201 554
rect 1220 553 1221 554
rect 1203 555 1204 556
rect 1216 555 1217 556
rect 1229 555 1230 556
rect 1235 555 1236 556
rect 1009 564 1010 565
rect 1015 564 1016 565
rect 1024 564 1025 565
rect 1028 564 1029 565
rect 1028 566 1029 567
rect 1077 566 1078 567
rect 1032 568 1033 569
rect 1099 568 1100 569
rect 1034 570 1035 571
rect 1045 570 1046 571
rect 1039 572 1040 573
rect 1068 572 1069 573
rect 1043 574 1044 575
rect 1074 574 1075 575
rect 1042 576 1043 577
rect 1215 576 1216 577
rect 1056 578 1057 579
rect 1074 578 1075 579
rect 1057 580 1058 581
rect 1113 580 1114 581
rect 1062 582 1063 583
rect 1080 582 1081 583
rect 1061 584 1062 585
rect 1098 584 1099 585
rect 1064 586 1065 587
rect 1122 586 1123 587
rect 1071 588 1072 589
rect 1110 588 1111 589
rect 1083 590 1084 591
rect 1119 590 1120 591
rect 1025 592 1026 593
rect 1083 592 1084 593
rect 1086 592 1087 593
rect 1127 592 1128 593
rect 1102 594 1103 595
rect 1104 594 1105 595
rect 1115 594 1116 595
rect 1152 594 1153 595
rect 1130 596 1131 597
rect 1137 596 1138 597
rect 1124 598 1125 599
rect 1131 598 1132 599
rect 1154 598 1155 599
rect 1194 598 1195 599
rect 1145 600 1146 601
rect 1155 600 1156 601
rect 1170 600 1171 601
rect 1176 600 1177 601
rect 1173 602 1174 603
rect 1209 602 1210 603
rect 1182 604 1183 605
rect 1185 604 1186 605
rect 1182 606 1183 607
rect 1200 606 1201 607
rect 1203 606 1204 607
rect 1242 606 1243 607
rect 1148 608 1149 609
rect 1203 608 1204 609
rect 1089 610 1090 611
rect 1149 610 1150 611
rect 1206 610 1207 611
rect 1218 610 1219 611
rect 1142 612 1143 613
rect 1206 612 1207 613
rect 1223 612 1224 613
rect 1233 612 1234 613
rect 1226 614 1227 615
rect 1279 614 1280 615
rect 1220 616 1221 617
rect 1227 616 1228 617
rect 1229 616 1230 617
rect 1282 616 1283 617
rect 1197 618 1198 619
rect 1230 618 1231 619
rect 1021 627 1022 628
rect 1096 627 1097 628
rect 1035 629 1036 630
rect 1083 629 1084 630
rect 1015 631 1016 632
rect 1034 631 1035 632
rect 1039 631 1040 632
rect 1135 631 1136 632
rect 1049 633 1050 634
rect 1122 633 1123 634
rect 1052 635 1053 636
rect 1077 635 1078 636
rect 1054 637 1055 638
rect 1171 637 1172 638
rect 1057 639 1058 640
rect 1083 639 1084 640
rect 1061 641 1062 642
rect 1141 641 1142 642
rect 1045 643 1046 644
rect 1062 643 1063 644
rect 1064 643 1065 644
rect 1168 643 1169 644
rect 1071 645 1072 646
rect 1119 645 1120 646
rect 1074 647 1075 648
rect 1102 647 1103 648
rect 1080 649 1081 650
rect 1108 649 1109 650
rect 1040 651 1041 652
rect 1080 651 1081 652
rect 1089 651 1090 652
rect 1267 651 1268 652
rect 1090 653 1091 654
rect 1104 653 1105 654
rect 1098 655 1099 656
rect 1147 655 1148 656
rect 1113 657 1114 658
rect 1165 657 1166 658
rect 1114 659 1115 660
rect 1186 659 1187 660
rect 1117 661 1118 662
rect 1155 661 1156 662
rect 1125 663 1126 664
rect 1152 663 1153 664
rect 1110 665 1111 666
rect 1153 665 1154 666
rect 1025 667 1026 668
rect 1111 667 1112 668
rect 1024 669 1025 670
rect 1037 669 1038 670
rect 1126 669 1127 670
rect 1224 669 1225 670
rect 1128 671 1129 672
rect 1137 671 1138 672
rect 1042 673 1043 674
rect 1138 673 1139 674
rect 1149 673 1150 674
rect 1162 673 1163 674
rect 1173 673 1174 674
rect 1201 673 1202 674
rect 1174 675 1175 676
rect 1206 675 1207 676
rect 1176 677 1177 678
rect 1225 677 1226 678
rect 1189 679 1190 680
rect 1203 679 1204 680
rect 1192 681 1193 682
rect 1212 681 1213 682
rect 1194 683 1195 684
rect 1246 683 1247 684
rect 1204 685 1205 686
rect 1221 685 1222 686
rect 1207 687 1208 688
rect 1209 687 1210 688
rect 1131 689 1132 690
rect 1210 689 1211 690
rect 1213 689 1214 690
rect 1218 689 1219 690
rect 1215 691 1216 692
rect 1270 691 1271 692
rect 1219 693 1220 694
rect 1300 693 1301 694
rect 1227 695 1228 696
rect 1273 695 1274 696
rect 1233 697 1234 698
rect 1291 697 1292 698
rect 1242 699 1243 700
rect 1294 699 1295 700
rect 1259 701 1260 702
rect 1285 701 1286 702
rect 1276 703 1277 704
rect 1288 703 1289 704
rect 1230 705 1231 706
rect 1288 705 1289 706
rect 1182 707 1183 708
rect 1231 707 1232 708
rect 1279 707 1280 708
rect 1337 707 1338 708
rect 1279 709 1280 710
rect 1282 709 1283 710
rect 1198 711 1199 712
rect 1282 711 1283 712
rect 1297 711 1298 712
rect 1307 711 1308 712
rect 1334 711 1335 712
rect 1344 711 1345 712
rect 1015 720 1016 721
rect 1183 720 1184 721
rect 1018 722 1019 723
rect 1111 722 1112 723
rect 1021 724 1022 725
rect 1064 724 1065 725
rect 1031 726 1032 727
rect 1096 726 1097 727
rect 1028 728 1029 729
rect 1032 728 1033 729
rect 1049 728 1050 729
rect 1171 728 1172 729
rect 1048 730 1049 731
rect 1177 730 1178 731
rect 1059 732 1060 733
rect 1080 732 1081 733
rect 1062 734 1063 735
rect 1067 734 1068 735
rect 1071 734 1072 735
rect 1165 734 1166 735
rect 1070 736 1071 737
rect 1195 736 1196 737
rect 1074 738 1075 739
rect 1159 738 1160 739
rect 1090 740 1091 741
rect 1165 740 1166 741
rect 1077 742 1078 743
rect 1089 742 1090 743
rect 1102 742 1103 743
rect 1120 742 1121 743
rect 1105 744 1106 745
rect 1153 744 1154 745
rect 1041 746 1042 747
rect 1153 746 1154 747
rect 1108 748 1109 749
rect 1117 748 1118 749
rect 1114 750 1115 751
rect 1162 750 1163 751
rect 1129 752 1130 753
rect 1141 752 1142 753
rect 1138 754 1139 755
rect 1156 754 1157 755
rect 1186 754 1187 755
rect 1243 754 1244 755
rect 1126 756 1127 757
rect 1186 756 1187 757
rect 1192 756 1193 757
rect 1249 756 1250 757
rect 1198 758 1199 759
rect 1228 758 1229 759
rect 1168 760 1169 761
rect 1198 760 1199 761
rect 1083 762 1084 763
rect 1168 762 1169 763
rect 1201 762 1202 763
rect 1252 762 1253 763
rect 1204 764 1205 765
rect 1261 764 1262 765
rect 1213 766 1214 767
rect 1285 766 1286 767
rect 1225 768 1226 769
rect 1285 768 1286 769
rect 1052 770 1053 771
rect 1225 770 1226 771
rect 1240 770 1241 771
rect 1433 770 1434 771
rect 1255 772 1256 773
rect 1366 772 1367 773
rect 1267 774 1268 775
rect 1357 774 1358 775
rect 1246 776 1247 777
rect 1267 776 1268 777
rect 1189 778 1190 779
rect 1246 778 1247 779
rect 1073 780 1074 781
rect 1189 780 1190 781
rect 1270 780 1271 781
rect 1360 780 1361 781
rect 1273 782 1274 783
rect 1375 782 1376 783
rect 1207 784 1208 785
rect 1273 784 1274 785
rect 1174 786 1175 787
rect 1207 786 1208 787
rect 1276 786 1277 787
rect 1339 786 1340 787
rect 1279 788 1280 789
rect 1342 788 1343 789
rect 1219 790 1220 791
rect 1279 790 1280 791
rect 1288 790 1289 791
rect 1410 790 1411 791
rect 1294 792 1295 793
rect 1387 792 1388 793
rect 1297 794 1298 795
rect 1327 794 1328 795
rect 1303 796 1304 797
rect 1321 796 1322 797
rect 1291 798 1292 799
rect 1303 798 1304 799
rect 1234 800 1235 801
rect 1291 800 1292 801
rect 1307 800 1308 801
rect 1390 800 1391 801
rect 1231 802 1232 803
rect 1306 802 1307 803
rect 1324 802 1325 803
rect 1348 802 1349 803
rect 1334 804 1335 805
rect 1427 804 1428 805
rect 1310 806 1311 807
rect 1333 806 1334 807
rect 1344 806 1345 807
rect 1350 806 1351 807
rect 1345 808 1346 809
rect 1407 808 1408 809
rect 1378 810 1379 811
rect 1384 810 1385 811
rect 955 819 956 820
rect 962 819 963 820
rect 993 819 994 820
rect 1035 819 1036 820
rect 1012 821 1013 822
rect 1026 821 1027 822
rect 1016 823 1017 824
rect 1064 823 1065 824
rect 1029 825 1030 826
rect 1132 825 1133 826
rect 1019 827 1020 828
rect 1030 827 1031 828
rect 1038 827 1039 828
rect 1052 827 1053 828
rect 1033 829 1034 830
rect 1037 829 1038 830
rect 1052 829 1053 830
rect 1067 829 1068 830
rect 1055 831 1056 832
rect 1306 831 1307 832
rect 1058 833 1059 834
rect 1135 833 1136 834
rect 1065 835 1066 836
rect 1162 835 1163 836
rect 1068 837 1069 838
rect 1089 837 1090 838
rect 1070 839 1071 840
rect 1177 839 1178 840
rect 1071 841 1072 842
rect 1393 841 1394 842
rect 1077 843 1078 844
rect 1189 843 1190 844
rect 1078 845 1079 846
rect 1324 845 1325 846
rect 1080 847 1081 848
rect 1095 847 1096 848
rect 1090 849 1091 850
rect 1117 849 1118 850
rect 1105 851 1106 852
rect 1276 851 1277 852
rect 1108 853 1109 854
rect 1183 853 1184 854
rect 1120 855 1121 856
rect 1135 855 1136 856
rect 1009 857 1010 858
rect 1120 857 1121 858
rect 1123 857 1124 858
rect 1186 857 1187 858
rect 1129 859 1130 860
rect 1201 859 1202 860
rect 1138 861 1139 862
rect 1147 861 1148 862
rect 1144 863 1145 864
rect 1153 863 1154 864
rect 1147 865 1148 866
rect 1156 865 1157 866
rect 1074 867 1075 868
rect 1156 867 1157 868
rect 1150 869 1151 870
rect 1225 869 1226 870
rect 1159 871 1160 872
rect 1264 871 1265 872
rect 1165 873 1166 874
rect 1213 873 1214 874
rect 1048 875 1049 876
rect 1165 875 1166 876
rect 1022 877 1023 878
rect 1049 877 1050 878
rect 1174 877 1175 878
rect 1240 877 1241 878
rect 1183 879 1184 880
rect 1381 879 1382 880
rect 1189 881 1190 882
rect 1261 881 1262 882
rect 1198 883 1199 884
rect 1204 883 1205 884
rect 1207 883 1208 884
rect 1306 883 1307 884
rect 1219 885 1220 886
rect 1285 885 1286 886
rect 1225 887 1226 888
rect 1249 887 1250 888
rect 1228 889 1229 890
rect 1294 889 1295 890
rect 1234 891 1235 892
rect 1258 891 1259 892
rect 1243 893 1244 894
rect 1309 893 1310 894
rect 1243 895 1244 896
rect 1342 895 1343 896
rect 1246 897 1247 898
rect 1363 897 1364 898
rect 1249 899 1250 900
rect 1447 899 1448 900
rect 1252 901 1253 902
rect 1366 901 1367 902
rect 1252 903 1253 904
rect 1279 903 1280 904
rect 1168 905 1169 906
rect 1279 905 1280 906
rect 1168 907 1169 908
rect 1195 907 1196 908
rect 1195 909 1196 910
rect 1439 909 1440 910
rect 1255 911 1256 912
rect 1384 911 1385 912
rect 1267 913 1268 914
rect 1414 913 1415 914
rect 1270 915 1271 916
rect 1473 915 1474 916
rect 1282 917 1283 918
rect 1300 917 1301 918
rect 1318 917 1319 918
rect 1417 917 1418 918
rect 1321 919 1322 920
rect 1400 919 1401 920
rect 1321 921 1322 922
rect 1348 921 1349 922
rect 1207 923 1208 924
rect 1348 923 1349 924
rect 1339 925 1340 926
rect 1354 925 1355 926
rect 1351 927 1352 928
rect 1469 927 1470 928
rect 1357 929 1358 930
rect 1369 929 1370 930
rect 1360 931 1361 932
rect 1372 931 1373 932
rect 1363 933 1364 934
rect 1384 933 1385 934
rect 1375 935 1376 936
rect 1399 935 1400 936
rect 1378 937 1379 938
rect 1402 937 1403 938
rect 1387 939 1388 940
rect 1405 939 1406 940
rect 1387 941 1388 942
rect 1410 941 1411 942
rect 1273 943 1274 944
rect 1411 943 1412 944
rect 1390 945 1391 946
rect 1408 945 1409 946
rect 1303 947 1304 948
rect 1390 947 1391 948
rect 1396 947 1397 948
rect 1432 947 1433 948
rect 1345 949 1346 950
rect 1396 949 1397 950
rect 1102 951 1103 952
rect 1345 951 1346 952
rect 1423 951 1424 952
rect 1460 951 1461 952
rect 1427 953 1428 954
rect 1463 953 1464 954
rect 1426 955 1427 956
rect 1457 955 1458 956
rect 1437 957 1438 958
rect 1444 957 1445 958
rect 979 966 980 967
rect 986 966 987 967
rect 989 966 990 967
rect 993 966 994 967
rect 1012 966 1013 967
rect 1108 966 1109 967
rect 1019 968 1020 969
rect 1120 968 1121 969
rect 1023 970 1024 971
rect 1049 970 1050 971
rect 1026 972 1027 973
rect 1132 972 1133 973
rect 1030 974 1031 975
rect 1055 974 1056 975
rect 1030 976 1031 977
rect 1162 976 1163 977
rect 1033 978 1034 979
rect 1171 978 1172 979
rect 1050 980 1051 981
rect 1052 980 1053 981
rect 1068 980 1069 981
rect 1072 980 1073 981
rect 1074 980 1075 981
rect 1309 980 1310 981
rect 1037 982 1038 983
rect 1075 982 1076 983
rect 1037 984 1038 985
rect 1078 984 1079 985
rect 1090 984 1091 985
rect 1102 984 1103 985
rect 1090 986 1091 987
rect 1276 986 1277 987
rect 1105 988 1106 989
rect 1135 988 1136 989
rect 1120 990 1121 991
rect 1123 990 1124 991
rect 1129 990 1130 991
rect 1138 990 1139 991
rect 1135 992 1136 993
rect 1144 992 1145 993
rect 1141 994 1142 995
rect 1201 994 1202 995
rect 1147 996 1148 997
rect 1186 996 1187 997
rect 1147 998 1148 999
rect 1264 998 1265 999
rect 1153 1000 1154 1001
rect 1168 1000 1169 1001
rect 1159 1002 1160 1003
rect 1213 1002 1214 1003
rect 1066 1004 1067 1005
rect 1213 1004 1214 1005
rect 1165 1006 1166 1007
rect 1192 1006 1193 1007
rect 1156 1008 1157 1009
rect 1165 1008 1166 1009
rect 1156 1010 1157 1011
rect 1204 1010 1205 1011
rect 1174 1012 1175 1013
rect 1216 1012 1217 1013
rect 1177 1014 1178 1015
rect 1436 1014 1437 1015
rect 1183 1016 1184 1017
rect 1240 1016 1241 1017
rect 1047 1018 1048 1019
rect 1183 1018 1184 1019
rect 1189 1018 1190 1019
rect 1228 1018 1229 1019
rect 1150 1020 1151 1021
rect 1189 1020 1190 1021
rect 1195 1020 1196 1021
rect 1234 1020 1235 1021
rect 1195 1022 1196 1023
rect 1201 1022 1202 1023
rect 1198 1024 1199 1025
rect 1279 1024 1280 1025
rect 1207 1026 1208 1027
rect 1246 1026 1247 1027
rect 1243 1028 1244 1029
rect 1294 1028 1295 1029
rect 1249 1030 1250 1031
rect 1291 1030 1292 1031
rect 1258 1032 1259 1033
rect 1264 1032 1265 1033
rect 1225 1034 1226 1035
rect 1258 1034 1259 1035
rect 1270 1034 1271 1035
rect 1312 1034 1313 1035
rect 1276 1036 1277 1037
rect 1458 1036 1459 1037
rect 1282 1038 1283 1039
rect 1285 1038 1286 1039
rect 1300 1038 1301 1039
rect 1324 1038 1325 1039
rect 1306 1040 1307 1041
rect 1384 1040 1385 1041
rect 1327 1042 1328 1043
rect 1336 1042 1337 1043
rect 1333 1044 1334 1045
rect 1342 1044 1343 1045
rect 1348 1044 1349 1045
rect 1396 1044 1397 1045
rect 1354 1046 1355 1047
rect 1476 1046 1477 1047
rect 1318 1048 1319 1049
rect 1354 1048 1355 1049
rect 1318 1050 1319 1051
rect 1363 1050 1364 1051
rect 1357 1052 1358 1053
rect 1408 1052 1409 1053
rect 1375 1054 1376 1055
rect 1414 1054 1415 1055
rect 1387 1056 1388 1057
rect 1449 1056 1450 1057
rect 1369 1058 1370 1059
rect 1387 1058 1388 1059
rect 1369 1060 1370 1061
rect 1469 1060 1470 1061
rect 1390 1062 1391 1063
rect 1455 1062 1456 1063
rect 1372 1064 1373 1065
rect 1390 1064 1391 1065
rect 1351 1066 1352 1067
rect 1372 1066 1373 1067
rect 1321 1068 1322 1069
rect 1351 1068 1352 1069
rect 1321 1070 1322 1071
rect 1366 1070 1367 1071
rect 1402 1070 1403 1071
rect 1418 1070 1419 1071
rect 1222 1072 1223 1073
rect 1403 1072 1404 1073
rect 1405 1072 1406 1073
rect 1409 1072 1410 1073
rect 1399 1074 1400 1075
rect 1406 1074 1407 1075
rect 1330 1076 1331 1077
rect 1400 1076 1401 1077
rect 1412 1076 1413 1077
rect 1432 1076 1433 1077
rect 1423 1078 1424 1079
rect 1443 1078 1444 1079
rect 1252 1080 1253 1081
rect 1422 1080 1423 1081
rect 1252 1082 1253 1083
rect 1475 1082 1476 1083
rect 1426 1084 1427 1085
rect 1428 1084 1429 1085
rect 1440 1084 1441 1085
rect 1460 1084 1461 1085
rect 1219 1086 1220 1087
rect 1461 1086 1462 1087
rect 1081 1088 1082 1089
rect 1219 1088 1220 1089
rect 1452 1088 1453 1089
rect 1466 1088 1467 1089
rect 1463 1090 1464 1091
rect 1465 1090 1466 1091
rect 1006 1099 1007 1100
rect 1035 1099 1036 1100
rect 1012 1101 1013 1102
rect 1057 1101 1058 1102
rect 1013 1103 1014 1104
rect 1054 1103 1055 1104
rect 1033 1105 1034 1106
rect 1156 1105 1157 1106
rect 1037 1107 1038 1108
rect 1118 1107 1119 1108
rect 1040 1109 1041 1110
rect 1072 1109 1073 1110
rect 1041 1111 1042 1112
rect 1060 1111 1061 1112
rect 1047 1113 1048 1114
rect 1075 1113 1076 1114
rect 1048 1115 1049 1116
rect 1115 1115 1116 1116
rect 1050 1117 1051 1118
rect 1066 1117 1067 1118
rect 1062 1119 1063 1120
rect 1192 1119 1193 1120
rect 1069 1121 1070 1122
rect 1141 1121 1142 1122
rect 1038 1123 1039 1124
rect 1069 1123 1070 1124
rect 1076 1123 1077 1124
rect 1243 1123 1244 1124
rect 1078 1125 1079 1126
rect 1383 1125 1384 1126
rect 1081 1127 1082 1128
rect 1147 1127 1148 1128
rect 1094 1129 1095 1130
rect 1105 1129 1106 1130
rect 1100 1131 1101 1132
rect 1102 1131 1103 1132
rect 1019 1133 1020 1134
rect 1103 1133 1104 1134
rect 1020 1135 1021 1136
rect 1264 1135 1265 1136
rect 1106 1137 1107 1138
rect 1120 1137 1121 1138
rect 1026 1139 1027 1140
rect 1121 1139 1122 1140
rect 1109 1141 1110 1142
rect 1195 1141 1196 1142
rect 1129 1143 1130 1144
rect 1204 1143 1205 1144
rect 1135 1145 1136 1146
rect 1175 1145 1176 1146
rect 1148 1147 1149 1148
rect 1171 1147 1172 1148
rect 1153 1149 1154 1150
rect 1226 1149 1227 1150
rect 1154 1151 1155 1152
rect 1422 1151 1423 1152
rect 1165 1153 1166 1154
rect 1181 1153 1182 1154
rect 1166 1155 1167 1156
rect 1177 1155 1178 1156
rect 1172 1157 1173 1158
rect 1183 1157 1184 1158
rect 1090 1159 1091 1160
rect 1184 1159 1185 1160
rect 1178 1161 1179 1162
rect 1189 1161 1190 1162
rect 1159 1163 1160 1164
rect 1190 1163 1191 1164
rect 1063 1165 1064 1166
rect 1160 1165 1161 1166
rect 1186 1165 1187 1166
rect 1211 1165 1212 1166
rect 1193 1167 1194 1168
rect 1198 1167 1199 1168
rect 1201 1167 1202 1168
rect 1213 1167 1214 1168
rect 1044 1169 1045 1170
rect 1202 1169 1203 1170
rect 1044 1171 1045 1172
rect 1130 1171 1131 1172
rect 1205 1171 1206 1172
rect 1216 1171 1217 1172
rect 1214 1173 1215 1174
rect 1222 1173 1223 1174
rect 1228 1175 1229 1176
rect 1400 1175 1401 1176
rect 1229 1177 1230 1178
rect 1246 1177 1247 1178
rect 1234 1179 1235 1180
rect 1425 1179 1426 1180
rect 1235 1181 1236 1182
rect 1252 1181 1253 1182
rect 1247 1183 1248 1184
rect 1285 1183 1286 1184
rect 1253 1185 1254 1186
rect 1276 1185 1277 1186
rect 1256 1187 1257 1188
rect 1455 1187 1456 1188
rect 1262 1189 1263 1190
rect 1300 1189 1301 1190
rect 1268 1191 1269 1192
rect 1294 1191 1295 1192
rect 1274 1193 1275 1194
rect 1291 1193 1292 1194
rect 1289 1195 1290 1196
rect 1312 1195 1313 1196
rect 1301 1197 1302 1198
rect 1396 1197 1397 1198
rect 1304 1199 1305 1200
rect 1321 1199 1322 1200
rect 1307 1201 1308 1202
rect 1336 1201 1337 1202
rect 1313 1203 1314 1204
rect 1342 1203 1343 1204
rect 1318 1205 1319 1206
rect 1393 1205 1394 1206
rect 1319 1207 1320 1208
rect 1330 1207 1331 1208
rect 1325 1209 1326 1210
rect 1416 1209 1417 1210
rect 1331 1211 1332 1212
rect 1390 1211 1391 1212
rect 1337 1213 1338 1214
rect 1354 1213 1355 1214
rect 1346 1215 1347 1216
rect 1369 1215 1370 1216
rect 1351 1217 1352 1218
rect 1355 1217 1356 1218
rect 1348 1219 1349 1220
rect 1352 1219 1353 1220
rect 1349 1221 1350 1222
rect 1372 1221 1373 1222
rect 1357 1223 1358 1224
rect 1431 1223 1432 1224
rect 1358 1225 1359 1226
rect 1375 1225 1376 1226
rect 1258 1227 1259 1228
rect 1376 1227 1377 1228
rect 1389 1227 1390 1228
rect 1406 1227 1407 1228
rect 1392 1229 1393 1230
rect 1446 1229 1447 1230
rect 1395 1231 1396 1232
rect 1409 1231 1410 1232
rect 1387 1233 1388 1234
rect 1410 1233 1411 1234
rect 1386 1235 1387 1236
rect 1443 1235 1444 1236
rect 1398 1237 1399 1238
rect 1412 1237 1413 1238
rect 1401 1239 1402 1240
rect 1418 1239 1419 1240
rect 1404 1241 1405 1242
rect 1425 1241 1426 1242
rect 1407 1243 1408 1244
rect 1475 1243 1476 1244
rect 1413 1245 1414 1246
rect 1428 1245 1429 1246
rect 1422 1247 1423 1248
rect 1452 1247 1453 1248
rect 1438 1249 1439 1250
rect 1465 1249 1466 1250
rect 1440 1251 1441 1252
rect 1472 1251 1473 1252
rect 994 1260 995 1261
rect 998 1260 999 1261
rect 1006 1260 1007 1261
rect 1051 1260 1052 1261
rect 1013 1262 1014 1263
rect 1029 1262 1030 1263
rect 1020 1264 1021 1265
rect 1143 1264 1144 1265
rect 1008 1266 1009 1267
rect 1019 1266 1020 1267
rect 1022 1266 1023 1267
rect 1158 1266 1159 1267
rect 1026 1268 1027 1269
rect 1118 1268 1119 1269
rect 1035 1270 1036 1271
rect 1050 1270 1051 1271
rect 1066 1270 1067 1271
rect 1211 1270 1212 1271
rect 1069 1272 1070 1273
rect 1181 1272 1182 1273
rect 1010 1274 1011 1275
rect 1069 1274 1070 1275
rect 1076 1274 1077 1275
rect 1208 1274 1209 1275
rect 1054 1276 1055 1277
rect 1075 1276 1076 1277
rect 1038 1278 1039 1279
rect 1053 1278 1054 1279
rect 1091 1278 1092 1279
rect 1160 1278 1161 1279
rect 1094 1280 1095 1281
rect 1260 1280 1261 1281
rect 1106 1282 1107 1283
rect 1146 1282 1147 1283
rect 1100 1284 1101 1285
rect 1106 1284 1107 1285
rect 1115 1284 1116 1285
rect 1386 1284 1387 1285
rect 1125 1286 1126 1287
rect 1239 1286 1240 1287
rect 1128 1288 1129 1289
rect 1190 1288 1191 1289
rect 1072 1290 1073 1291
rect 1191 1290 1192 1291
rect 1154 1292 1155 1293
rect 1161 1292 1162 1293
rect 1044 1294 1045 1295
rect 1155 1294 1156 1295
rect 1005 1296 1006 1297
rect 1044 1296 1045 1297
rect 1184 1296 1185 1297
rect 1251 1296 1252 1297
rect 1178 1298 1179 1299
rect 1185 1298 1186 1299
rect 1166 1300 1167 1301
rect 1179 1300 1180 1301
rect 1220 1300 1221 1301
rect 1223 1300 1224 1301
rect 1202 1302 1203 1303
rect 1221 1302 1222 1303
rect 1203 1304 1204 1305
rect 1205 1304 1206 1305
rect 1224 1304 1225 1305
rect 1383 1304 1384 1305
rect 1226 1306 1227 1307
rect 1473 1306 1474 1307
rect 1088 1308 1089 1309
rect 1227 1308 1228 1309
rect 1229 1308 1230 1309
rect 1245 1308 1246 1309
rect 1121 1310 1122 1311
rect 1230 1310 1231 1311
rect 1121 1312 1122 1313
rect 1137 1312 1138 1313
rect 1235 1312 1236 1313
rect 1486 1312 1487 1313
rect 1247 1314 1248 1315
rect 1446 1314 1447 1315
rect 1253 1316 1254 1317
rect 1497 1316 1498 1317
rect 1193 1318 1194 1319
rect 1254 1318 1255 1319
rect 1148 1320 1149 1321
rect 1194 1320 1195 1321
rect 1130 1322 1131 1323
rect 1149 1322 1150 1323
rect 1131 1324 1132 1325
rect 1175 1324 1176 1325
rect 1081 1326 1082 1327
rect 1176 1326 1177 1327
rect 1262 1326 1263 1327
rect 1284 1326 1285 1327
rect 1256 1328 1257 1329
rect 1263 1328 1264 1329
rect 1274 1328 1275 1329
rect 1281 1328 1282 1329
rect 1289 1328 1290 1329
rect 1296 1328 1297 1329
rect 1079 1330 1080 1331
rect 1290 1330 1291 1331
rect 1057 1332 1058 1333
rect 1078 1332 1079 1333
rect 1056 1334 1057 1335
rect 1103 1334 1104 1335
rect 1307 1334 1308 1335
rect 1437 1334 1438 1335
rect 1308 1336 1309 1337
rect 1425 1336 1426 1337
rect 1313 1338 1314 1339
rect 1435 1338 1436 1339
rect 1325 1340 1326 1341
rect 1404 1340 1405 1341
rect 1301 1342 1302 1343
rect 1404 1342 1405 1343
rect 1302 1344 1303 1345
rect 1461 1344 1462 1345
rect 1331 1346 1332 1347
rect 1416 1346 1417 1347
rect 1319 1348 1320 1349
rect 1332 1348 1333 1349
rect 1320 1350 1321 1351
rect 1514 1350 1515 1351
rect 1337 1352 1338 1353
rect 1344 1352 1345 1353
rect 1346 1352 1347 1353
rect 1365 1352 1366 1353
rect 1347 1354 1348 1355
rect 1355 1354 1356 1355
rect 1349 1356 1350 1357
rect 1368 1356 1369 1357
rect 1356 1358 1357 1359
rect 1380 1358 1381 1359
rect 1358 1360 1359 1361
rect 1428 1360 1429 1361
rect 1383 1362 1384 1363
rect 1410 1362 1411 1363
rect 1352 1364 1353 1365
rect 1410 1364 1411 1365
rect 1353 1366 1354 1367
rect 1376 1366 1377 1367
rect 1389 1366 1390 1367
rect 1428 1366 1429 1367
rect 1389 1368 1390 1369
rect 1504 1368 1505 1369
rect 1395 1370 1396 1371
rect 1434 1370 1435 1371
rect 1398 1372 1399 1373
rect 1431 1372 1432 1373
rect 1392 1374 1393 1375
rect 1431 1374 1432 1375
rect 1401 1376 1402 1377
rect 1443 1376 1444 1377
rect 1407 1378 1408 1379
rect 1470 1378 1471 1379
rect 1304 1380 1305 1381
rect 1407 1380 1408 1381
rect 1416 1380 1417 1381
rect 1440 1380 1441 1381
rect 1422 1382 1423 1383
rect 1464 1382 1465 1383
rect 1452 1384 1453 1385
rect 1455 1384 1456 1385
rect 1413 1386 1414 1387
rect 1452 1386 1453 1387
rect 1467 1386 1468 1387
rect 1493 1386 1494 1387
rect 1008 1395 1009 1396
rect 1053 1395 1054 1396
rect 1015 1397 1016 1398
rect 1081 1397 1082 1398
rect 1019 1399 1020 1400
rect 1124 1399 1125 1400
rect 1019 1401 1020 1402
rect 1069 1401 1070 1402
rect 1038 1403 1039 1404
rect 1066 1403 1067 1404
rect 998 1405 999 1406
rect 1066 1405 1067 1406
rect 1041 1407 1042 1408
rect 1044 1407 1045 1408
rect 1053 1407 1054 1408
rect 1093 1407 1094 1408
rect 1059 1409 1060 1410
rect 1158 1409 1159 1410
rect 1063 1411 1064 1412
rect 1191 1411 1192 1412
rect 1001 1413 1002 1414
rect 1063 1413 1064 1414
rect 1000 1415 1001 1416
rect 1050 1415 1051 1416
rect 1084 1415 1085 1416
rect 1190 1415 1191 1416
rect 1088 1417 1089 1418
rect 1194 1417 1195 1418
rect 1087 1419 1088 1420
rect 1176 1419 1177 1420
rect 1106 1421 1107 1422
rect 1121 1421 1122 1422
rect 1100 1423 1101 1424
rect 1121 1423 1122 1424
rect 1118 1425 1119 1426
rect 1227 1425 1228 1426
rect 1118 1427 1119 1428
rect 1230 1427 1231 1428
rect 1143 1429 1144 1430
rect 1166 1429 1167 1430
rect 1016 1431 1017 1432
rect 1142 1431 1143 1432
rect 1146 1431 1147 1432
rect 1169 1431 1170 1432
rect 1057 1433 1058 1434
rect 1145 1433 1146 1434
rect 1173 1433 1174 1434
rect 1187 1433 1188 1434
rect 1155 1435 1156 1436
rect 1172 1435 1173 1436
rect 1149 1437 1150 1438
rect 1154 1437 1155 1438
rect 1137 1439 1138 1440
rect 1148 1439 1149 1440
rect 1131 1441 1132 1442
rect 1136 1441 1137 1442
rect 1179 1441 1180 1442
rect 1196 1441 1197 1442
rect 1178 1443 1179 1444
rect 1340 1443 1341 1444
rect 1185 1445 1186 1446
rect 1193 1445 1194 1446
rect 1199 1445 1200 1446
rect 1356 1445 1357 1446
rect 1215 1447 1216 1448
rect 1229 1447 1230 1448
rect 1217 1449 1218 1450
rect 1224 1449 1225 1450
rect 1223 1451 1224 1452
rect 1251 1451 1252 1452
rect 1226 1453 1227 1454
rect 1239 1453 1240 1454
rect 1235 1455 1236 1456
rect 1257 1455 1258 1456
rect 1128 1457 1129 1458
rect 1256 1457 1257 1458
rect 1078 1459 1079 1460
rect 1127 1459 1128 1460
rect 1241 1459 1242 1460
rect 1304 1459 1305 1460
rect 1245 1461 1246 1462
rect 1419 1461 1420 1462
rect 1254 1463 1255 1464
rect 1334 1463 1335 1464
rect 1253 1465 1254 1466
rect 1353 1465 1354 1466
rect 1260 1467 1261 1468
rect 1377 1467 1378 1468
rect 1259 1469 1260 1470
rect 1290 1469 1291 1470
rect 1263 1471 1264 1472
rect 1286 1471 1287 1472
rect 1265 1473 1266 1474
rect 1497 1473 1498 1474
rect 1284 1475 1285 1476
rect 1449 1475 1450 1476
rect 1281 1477 1282 1478
rect 1283 1477 1284 1478
rect 1308 1477 1309 1478
rect 1418 1477 1419 1478
rect 1302 1479 1303 1480
rect 1307 1479 1308 1480
rect 1310 1479 1311 1480
rect 1347 1479 1348 1480
rect 1316 1481 1317 1482
rect 1410 1481 1411 1482
rect 1320 1483 1321 1484
rect 1373 1483 1374 1484
rect 1328 1485 1329 1486
rect 1365 1485 1366 1486
rect 1332 1487 1333 1488
rect 1514 1487 1515 1488
rect 1269 1489 1270 1490
rect 1331 1489 1332 1490
rect 1337 1489 1338 1490
rect 1407 1489 1408 1490
rect 1344 1491 1345 1492
rect 1352 1491 1353 1492
rect 1346 1493 1347 1494
rect 1389 1493 1390 1494
rect 1349 1495 1350 1496
rect 1500 1495 1501 1496
rect 1355 1497 1356 1498
rect 1428 1497 1429 1498
rect 1262 1499 1263 1500
rect 1428 1499 1429 1500
rect 1358 1501 1359 1502
rect 1431 1501 1432 1502
rect 1368 1503 1369 1504
rect 1397 1503 1398 1504
rect 1370 1505 1371 1506
rect 1434 1505 1435 1506
rect 1376 1507 1377 1508
rect 1440 1507 1441 1508
rect 1296 1509 1297 1510
rect 1439 1509 1440 1510
rect 1380 1511 1381 1512
rect 1483 1511 1484 1512
rect 1379 1513 1380 1514
rect 1443 1513 1444 1514
rect 1367 1515 1368 1516
rect 1442 1515 1443 1516
rect 1388 1517 1389 1518
rect 1452 1517 1453 1518
rect 1391 1519 1392 1520
rect 1464 1519 1465 1520
rect 1394 1521 1395 1522
rect 1467 1521 1468 1522
rect 1400 1523 1401 1524
rect 1446 1523 1447 1524
rect 1404 1525 1405 1526
rect 1486 1525 1487 1526
rect 1383 1527 1384 1528
rect 1404 1527 1405 1528
rect 1407 1527 1408 1528
rect 1473 1527 1474 1528
rect 1437 1529 1438 1530
rect 1458 1529 1459 1530
rect 1455 1531 1456 1532
rect 1507 1531 1508 1532
rect 1470 1533 1471 1534
rect 1479 1533 1480 1534
rect 997 1542 998 1543
rect 1066 1542 1067 1543
rect 1016 1544 1017 1545
rect 1081 1544 1082 1545
rect 1024 1546 1025 1547
rect 1108 1546 1109 1547
rect 1031 1548 1032 1549
rect 1038 1548 1039 1549
rect 1035 1550 1036 1551
rect 1053 1550 1054 1551
rect 1026 1552 1027 1553
rect 1034 1552 1035 1553
rect 1027 1554 1028 1555
rect 1075 1554 1076 1555
rect 1041 1556 1042 1557
rect 1175 1556 1176 1557
rect 1043 1558 1044 1559
rect 1127 1558 1128 1559
rect 1052 1560 1053 1561
rect 1241 1560 1242 1561
rect 1057 1562 1058 1563
rect 1148 1562 1149 1563
rect 1056 1564 1057 1565
rect 1154 1564 1155 1565
rect 1063 1566 1064 1567
rect 1080 1566 1081 1567
rect 1068 1568 1069 1569
rect 1087 1568 1088 1569
rect 1086 1570 1087 1571
rect 1118 1570 1119 1571
rect 1019 1572 1020 1573
rect 1117 1572 1118 1573
rect 1020 1574 1021 1575
rect 1150 1574 1151 1575
rect 1100 1576 1101 1577
rect 1226 1576 1227 1577
rect 1102 1578 1103 1579
rect 1240 1578 1241 1579
rect 1124 1580 1125 1581
rect 1147 1580 1148 1581
rect 1136 1582 1137 1583
rect 1153 1582 1154 1583
rect 1160 1582 1161 1583
rect 1183 1582 1184 1583
rect 1012 1584 1013 1585
rect 1159 1584 1160 1585
rect 1169 1584 1170 1585
rect 1198 1584 1199 1585
rect 1145 1586 1146 1587
rect 1168 1586 1169 1587
rect 1172 1586 1173 1587
rect 1204 1586 1205 1587
rect 1060 1588 1061 1589
rect 1171 1588 1172 1589
rect 1059 1590 1060 1591
rect 1135 1590 1136 1591
rect 1177 1590 1178 1591
rect 1304 1590 1305 1591
rect 1187 1592 1188 1593
rect 1246 1592 1247 1593
rect 1186 1594 1187 1595
rect 1190 1594 1191 1595
rect 1074 1596 1075 1597
rect 1189 1596 1190 1597
rect 1196 1596 1197 1597
rect 1207 1596 1208 1597
rect 1166 1598 1167 1599
rect 1195 1598 1196 1599
rect 1142 1600 1143 1601
rect 1165 1600 1166 1601
rect 1201 1600 1202 1601
rect 1223 1600 1224 1601
rect 1050 1602 1051 1603
rect 1222 1602 1223 1603
rect 1217 1604 1218 1605
rect 1231 1604 1232 1605
rect 1220 1606 1221 1607
rect 1237 1606 1238 1607
rect 1193 1608 1194 1609
rect 1219 1608 1220 1609
rect 1225 1608 1226 1609
rect 1253 1608 1254 1609
rect 1229 1610 1230 1611
rect 1252 1610 1253 1611
rect 1228 1612 1229 1613
rect 1256 1612 1257 1613
rect 1235 1614 1236 1615
rect 1336 1614 1337 1615
rect 1249 1616 1250 1617
rect 1259 1616 1260 1617
rect 1262 1616 1263 1617
rect 1312 1616 1313 1617
rect 1265 1618 1266 1619
rect 1300 1618 1301 1619
rect 1243 1620 1244 1621
rect 1264 1620 1265 1621
rect 1283 1620 1284 1621
rect 1318 1620 1319 1621
rect 1286 1622 1287 1623
rect 1294 1622 1295 1623
rect 1310 1622 1311 1623
rect 1385 1622 1386 1623
rect 1316 1624 1317 1625
rect 1334 1624 1335 1625
rect 1315 1626 1316 1627
rect 1418 1626 1419 1627
rect 1333 1628 1334 1629
rect 1376 1628 1377 1629
rect 1346 1630 1347 1631
rect 1384 1630 1385 1631
rect 1345 1632 1346 1633
rect 1355 1632 1356 1633
rect 1349 1634 1350 1635
rect 1415 1634 1416 1635
rect 1348 1636 1349 1637
rect 1358 1636 1359 1637
rect 1352 1638 1353 1639
rect 1381 1638 1382 1639
rect 1340 1640 1341 1641
rect 1351 1640 1352 1641
rect 1339 1642 1340 1643
rect 1373 1642 1374 1643
rect 1331 1644 1332 1645
rect 1372 1644 1373 1645
rect 1354 1646 1355 1647
rect 1379 1646 1380 1647
rect 1367 1648 1368 1649
rect 1396 1648 1397 1649
rect 1370 1650 1371 1651
rect 1400 1650 1401 1651
rect 1328 1652 1329 1653
rect 1369 1652 1370 1653
rect 1327 1654 1328 1655
rect 1421 1654 1422 1655
rect 1388 1656 1389 1657
rect 1405 1656 1406 1657
rect 1387 1658 1388 1659
rect 1425 1658 1426 1659
rect 1391 1660 1392 1661
rect 1399 1660 1400 1661
rect 1270 1662 1271 1663
rect 1390 1662 1391 1663
rect 1394 1662 1395 1663
rect 1402 1662 1403 1663
rect 1288 1664 1289 1665
rect 1393 1664 1394 1665
rect 1407 1664 1408 1665
rect 1422 1664 1423 1665
rect 1342 1666 1343 1667
rect 1408 1666 1409 1667
rect 1006 1675 1007 1676
rect 1195 1675 1196 1676
rect 1010 1677 1011 1678
rect 1043 1677 1044 1678
rect 1013 1679 1014 1680
rect 1150 1679 1151 1680
rect 1003 1681 1004 1682
rect 1151 1681 1152 1682
rect 1017 1683 1018 1684
rect 1049 1683 1050 1684
rect 1020 1685 1021 1686
rect 1034 1685 1035 1686
rect 1009 1687 1010 1688
rect 1019 1687 1020 1688
rect 1024 1687 1025 1688
rect 1100 1687 1101 1688
rect 1030 1689 1031 1690
rect 1204 1689 1205 1690
rect 1037 1691 1038 1692
rect 1168 1691 1169 1692
rect 1059 1693 1060 1694
rect 1068 1693 1069 1694
rect 1059 1695 1060 1696
rect 1177 1695 1178 1696
rect 1062 1697 1063 1698
rect 1080 1697 1081 1698
rect 1068 1699 1069 1700
rect 1196 1699 1197 1700
rect 1077 1701 1078 1702
rect 1178 1701 1179 1702
rect 1079 1703 1080 1704
rect 1189 1703 1190 1704
rect 1083 1705 1084 1706
rect 1120 1705 1121 1706
rect 1082 1707 1083 1708
rect 1237 1707 1238 1708
rect 1097 1709 1098 1710
rect 1108 1709 1109 1710
rect 1102 1711 1103 1712
rect 1231 1711 1232 1712
rect 1105 1713 1106 1714
rect 1307 1713 1308 1714
rect 1106 1715 1107 1716
rect 1228 1715 1229 1716
rect 1115 1717 1116 1718
rect 1117 1717 1118 1718
rect 1118 1719 1119 1720
rect 1198 1719 1199 1720
rect 1127 1721 1128 1722
rect 1135 1721 1136 1722
rect 1133 1723 1134 1724
rect 1153 1723 1154 1724
rect 1139 1725 1140 1726
rect 1147 1725 1148 1726
rect 1142 1727 1143 1728
rect 1159 1727 1160 1728
rect 1056 1729 1057 1730
rect 1160 1729 1161 1730
rect 1148 1731 1149 1732
rect 1165 1731 1166 1732
rect 1154 1733 1155 1734
rect 1171 1733 1172 1734
rect 1172 1735 1173 1736
rect 1183 1735 1184 1736
rect 1175 1737 1176 1738
rect 1186 1737 1187 1738
rect 1184 1739 1185 1740
rect 1207 1739 1208 1740
rect 1187 1741 1188 1742
rect 1222 1741 1223 1742
rect 1199 1743 1200 1744
rect 1201 1743 1202 1744
rect 1202 1745 1203 1746
rect 1225 1745 1226 1746
rect 1205 1747 1206 1748
rect 1363 1747 1364 1748
rect 1208 1749 1209 1750
rect 1246 1749 1247 1750
rect 1211 1751 1212 1752
rect 1240 1751 1241 1752
rect 1219 1753 1220 1754
rect 1235 1753 1236 1754
rect 1220 1755 1221 1756
rect 1249 1755 1250 1756
rect 1229 1757 1230 1758
rect 1336 1757 1337 1758
rect 1232 1759 1233 1760
rect 1252 1759 1253 1760
rect 1265 1759 1266 1760
rect 1345 1759 1346 1760
rect 1267 1761 1268 1762
rect 1270 1761 1271 1762
rect 1268 1763 1269 1764
rect 1298 1763 1299 1764
rect 1283 1765 1284 1766
rect 1318 1765 1319 1766
rect 1288 1767 1289 1768
rect 1292 1767 1293 1768
rect 1289 1769 1290 1770
rect 1339 1769 1340 1770
rect 1294 1771 1295 1772
rect 1304 1771 1305 1772
rect 1295 1773 1296 1774
rect 1322 1773 1323 1774
rect 1300 1775 1301 1776
rect 1390 1775 1391 1776
rect 1301 1777 1302 1778
rect 1402 1777 1403 1778
rect 1310 1779 1311 1780
rect 1312 1779 1313 1780
rect 1313 1781 1314 1782
rect 1422 1781 1423 1782
rect 1315 1783 1316 1784
rect 1325 1783 1326 1784
rect 1316 1785 1317 1786
rect 1369 1785 1370 1786
rect 1319 1787 1320 1788
rect 1372 1787 1373 1788
rect 1327 1789 1328 1790
rect 1418 1789 1419 1790
rect 1328 1791 1329 1792
rect 1405 1791 1406 1792
rect 1331 1793 1332 1794
rect 1428 1793 1429 1794
rect 1333 1795 1334 1796
rect 1354 1795 1355 1796
rect 1337 1797 1338 1798
rect 1381 1797 1382 1798
rect 1334 1799 1335 1800
rect 1381 1799 1382 1800
rect 1342 1801 1343 1802
rect 1393 1801 1394 1802
rect 1348 1803 1349 1804
rect 1366 1803 1367 1804
rect 1347 1805 1348 1806
rect 1399 1805 1400 1806
rect 1354 1807 1355 1808
rect 1387 1807 1388 1808
rect 1360 1809 1361 1810
rect 1403 1809 1404 1810
rect 1363 1811 1364 1812
rect 1388 1811 1389 1812
rect 1375 1813 1376 1814
rect 1435 1813 1436 1814
rect 1378 1815 1379 1816
rect 1442 1815 1443 1816
rect 1384 1817 1385 1818
rect 1425 1817 1426 1818
rect 1396 1819 1397 1820
rect 1438 1819 1439 1820
rect 1012 1828 1013 1829
rect 1139 1828 1140 1829
rect 1012 1830 1013 1831
rect 1019 1830 1020 1831
rect 1016 1832 1017 1833
rect 1120 1832 1121 1833
rect 1023 1834 1024 1835
rect 1030 1834 1031 1835
rect 1033 1834 1034 1835
rect 1189 1834 1190 1835
rect 1040 1836 1041 1837
rect 1129 1836 1130 1837
rect 1044 1838 1045 1839
rect 1133 1838 1134 1839
rect 1047 1840 1048 1841
rect 1127 1840 1128 1841
rect 1056 1842 1057 1843
rect 1144 1842 1145 1843
rect 1059 1844 1060 1845
rect 1187 1844 1188 1845
rect 1060 1846 1061 1847
rect 1062 1846 1063 1847
rect 1063 1848 1064 1849
rect 1160 1848 1161 1849
rect 1065 1850 1066 1851
rect 1175 1850 1176 1851
rect 1066 1852 1067 1853
rect 1213 1852 1214 1853
rect 1070 1854 1071 1855
rect 1304 1854 1305 1855
rect 1080 1856 1081 1857
rect 1301 1856 1302 1857
rect 1084 1858 1085 1859
rect 1208 1858 1209 1859
rect 1103 1860 1104 1861
rect 1126 1860 1127 1861
rect 1097 1862 1098 1863
rect 1102 1862 1103 1863
rect 1096 1864 1097 1865
rect 1100 1864 1101 1865
rect 1151 1864 1152 1865
rect 1156 1864 1157 1865
rect 1154 1866 1155 1867
rect 1174 1866 1175 1867
rect 1148 1868 1149 1869
rect 1153 1868 1154 1869
rect 1142 1870 1143 1871
rect 1147 1870 1148 1871
rect 1026 1872 1027 1873
rect 1141 1872 1142 1873
rect 1165 1872 1166 1873
rect 1202 1872 1203 1873
rect 1184 1874 1185 1875
rect 1192 1874 1193 1875
rect 1183 1876 1184 1877
rect 1207 1876 1208 1877
rect 1205 1878 1206 1879
rect 1222 1878 1223 1879
rect 1217 1880 1218 1881
rect 1232 1880 1233 1881
rect 1211 1882 1212 1883
rect 1216 1882 1217 1883
rect 1210 1884 1211 1885
rect 1220 1884 1221 1885
rect 1123 1886 1124 1887
rect 1219 1886 1220 1887
rect 1229 1886 1230 1887
rect 1235 1886 1236 1887
rect 1228 1888 1229 1889
rect 1240 1888 1241 1889
rect 1249 1890 1250 1891
rect 1295 1890 1296 1891
rect 1252 1892 1253 1893
rect 1268 1892 1269 1893
rect 1255 1894 1256 1895
rect 1289 1894 1290 1895
rect 1265 1896 1266 1897
rect 1298 1896 1299 1897
rect 1264 1898 1265 1899
rect 1279 1898 1280 1899
rect 1273 1900 1274 1901
rect 1313 1900 1314 1901
rect 1276 1902 1277 1903
rect 1307 1902 1308 1903
rect 1288 1904 1289 1905
rect 1328 1904 1329 1905
rect 1292 1906 1293 1907
rect 1340 1906 1341 1907
rect 1291 1908 1292 1909
rect 1331 1908 1332 1909
rect 1294 1910 1295 1911
rect 1357 1910 1358 1911
rect 1297 1912 1298 1913
rect 1331 1912 1332 1913
rect 1303 1914 1304 1915
rect 1319 1914 1320 1915
rect 1310 1916 1311 1917
rect 1325 1916 1326 1917
rect 1199 1918 1200 1919
rect 1324 1918 1325 1919
rect 1196 1920 1197 1921
rect 1198 1920 1199 1921
rect 1178 1922 1179 1923
rect 1195 1922 1196 1923
rect 1314 1922 1315 1923
rect 1316 1922 1317 1923
rect 1334 1922 1335 1923
rect 1340 1922 1341 1923
rect 1334 1924 1335 1925
rect 1363 1924 1364 1925
rect 1337 1926 1338 1927
rect 1403 1926 1404 1927
rect 1283 1928 1284 1929
rect 1337 1928 1338 1929
rect 1347 1928 1348 1929
rect 1381 1928 1382 1929
rect 1364 1930 1365 1931
rect 1397 1930 1398 1931
rect 1375 1932 1376 1933
rect 1391 1932 1392 1933
rect 1360 1934 1361 1935
rect 1374 1934 1375 1935
rect 1378 1934 1379 1935
rect 1388 1934 1389 1935
rect 997 1943 998 1944
rect 1009 1943 1010 1944
rect 1019 1943 1020 1944
rect 1174 1943 1175 1944
rect 1012 1945 1013 1946
rect 1019 1945 1020 1946
rect 1023 1945 1024 1946
rect 1099 1945 1100 1946
rect 1023 1947 1024 1948
rect 1120 1947 1121 1948
rect 1030 1949 1031 1950
rect 1141 1949 1142 1950
rect 1033 1951 1034 1952
rect 1129 1951 1130 1952
rect 1035 1953 1036 1954
rect 1060 1953 1061 1954
rect 1052 1955 1053 1956
rect 1096 1955 1097 1956
rect 1057 1957 1058 1958
rect 1162 1957 1163 1958
rect 1059 1959 1060 1960
rect 1192 1959 1193 1960
rect 1066 1961 1067 1962
rect 1132 1961 1133 1962
rect 1087 1963 1088 1964
rect 1213 1963 1214 1964
rect 1090 1965 1091 1966
rect 1102 1965 1103 1966
rect 1093 1967 1094 1968
rect 1144 1967 1145 1968
rect 1096 1969 1097 1970
rect 1117 1969 1118 1970
rect 1102 1971 1103 1972
rect 1198 1971 1199 1972
rect 1105 1973 1106 1974
rect 1159 1973 1160 1974
rect 1114 1975 1115 1976
rect 1174 1975 1175 1976
rect 1120 1977 1121 1978
rect 1147 1977 1148 1978
rect 1126 1979 1127 1980
rect 1153 1979 1154 1980
rect 1129 1981 1130 1982
rect 1156 1981 1157 1982
rect 1141 1983 1142 1984
rect 1216 1983 1217 1984
rect 1150 1985 1151 1986
rect 1171 1985 1172 1986
rect 1070 1987 1071 1988
rect 1171 1987 1172 1988
rect 1063 1989 1064 1990
rect 1069 1989 1070 1990
rect 1153 1989 1154 1990
rect 1195 1989 1196 1990
rect 1156 1991 1157 1992
rect 1189 1991 1190 1992
rect 1183 1993 1184 1994
rect 1210 1993 1211 1994
rect 1183 1995 1184 1996
rect 1207 1995 1208 1996
rect 1195 1997 1196 1998
rect 1219 1997 1220 1998
rect 1084 1999 1085 2000
rect 1219 1999 1220 2000
rect 1045 2001 1046 2002
rect 1084 2001 1085 2002
rect 1198 2001 1199 2002
rect 1222 2001 1223 2002
rect 1165 2003 1166 2004
rect 1222 2003 1223 2004
rect 1073 2005 1074 2006
rect 1165 2005 1166 2006
rect 1201 2005 1202 2006
rect 1240 2005 1241 2006
rect 1204 2007 1205 2008
rect 1241 2007 1242 2008
rect 1213 2009 1214 2010
rect 1258 2009 1259 2010
rect 1228 2011 1229 2012
rect 1249 2011 1250 2012
rect 1232 2013 1233 2014
rect 1255 2013 1256 2014
rect 1237 2015 1238 2016
rect 1317 2015 1318 2016
rect 1247 2017 1248 2018
rect 1291 2017 1292 2018
rect 1252 2019 1253 2020
rect 1256 2019 1257 2020
rect 1229 2021 1230 2022
rect 1253 2021 1254 2022
rect 1259 2021 1260 2022
rect 1261 2021 1262 2022
rect 1226 2023 1227 2024
rect 1262 2023 1263 2024
rect 1279 2023 1280 2024
rect 1292 2023 1293 2024
rect 1264 2025 1265 2026
rect 1280 2025 1281 2026
rect 1288 2025 1289 2026
rect 1304 2025 1305 2026
rect 1294 2027 1295 2028
rect 1361 2027 1362 2028
rect 1276 2029 1277 2030
rect 1295 2029 1296 2030
rect 1277 2031 1278 2032
rect 1314 2031 1315 2032
rect 1297 2033 1298 2034
rect 1301 2033 1302 2034
rect 1298 2035 1299 2036
rect 1357 2035 1358 2036
rect 1307 2037 1308 2038
rect 1337 2037 1338 2038
rect 1323 2039 1324 2040
rect 1353 2039 1354 2040
rect 1328 2041 1329 2042
rect 1340 2041 1341 2042
rect 1334 2043 1335 2044
rect 1343 2043 1344 2044
rect 1307 2045 1308 2046
rect 1343 2045 1344 2046
rect 1367 2045 1368 2046
rect 1377 2045 1378 2046
rect 1000 2054 1001 2055
rect 1035 2054 1036 2055
rect 1016 2056 1017 2057
rect 1096 2056 1097 2057
rect 1026 2058 1027 2059
rect 1066 2058 1067 2059
rect 1034 2060 1035 2061
rect 1093 2060 1094 2061
rect 1041 2062 1042 2063
rect 1079 2062 1080 2063
rect 1043 2064 1044 2065
rect 1156 2064 1157 2065
rect 1045 2066 1046 2067
rect 1142 2066 1143 2067
rect 1048 2068 1049 2069
rect 1084 2068 1085 2069
rect 1050 2070 1051 2071
rect 1129 2070 1130 2071
rect 1052 2072 1053 2073
rect 1171 2072 1172 2073
rect 1059 2074 1060 2075
rect 1106 2074 1107 2075
rect 1082 2076 1083 2077
rect 1145 2076 1146 2077
rect 1085 2078 1086 2079
rect 1109 2078 1110 2079
rect 1094 2080 1095 2081
rect 1099 2080 1100 2081
rect 1102 2080 1103 2081
rect 1229 2080 1230 2081
rect 1090 2082 1091 2083
rect 1103 2082 1104 2083
rect 1126 2082 1127 2083
rect 1139 2082 1140 2083
rect 1073 2084 1074 2085
rect 1127 2084 1128 2085
rect 1150 2084 1151 2085
rect 1157 2084 1158 2085
rect 1162 2084 1163 2085
rect 1169 2084 1170 2085
rect 1055 2086 1056 2087
rect 1163 2086 1164 2087
rect 1165 2086 1166 2087
rect 1172 2086 1173 2087
rect 1159 2088 1160 2089
rect 1166 2088 1167 2089
rect 1153 2090 1154 2091
rect 1160 2090 1161 2091
rect 1178 2090 1179 2091
rect 1280 2090 1281 2091
rect 1183 2092 1184 2093
rect 1226 2092 1227 2093
rect 1198 2094 1199 2095
rect 1222 2094 1223 2095
rect 1201 2096 1202 2097
rect 1223 2096 1224 2097
rect 1186 2098 1187 2099
rect 1202 2098 1203 2099
rect 1204 2098 1205 2099
rect 1226 2098 1227 2099
rect 1205 2100 1206 2101
rect 1250 2100 1251 2101
rect 1232 2102 1233 2103
rect 1235 2102 1236 2103
rect 1190 2104 1191 2105
rect 1232 2104 1233 2105
rect 1244 2104 1245 2105
rect 1310 2104 1311 2105
rect 1244 2106 1245 2107
rect 1247 2106 1248 2107
rect 1253 2106 1254 2107
rect 1268 2106 1269 2107
rect 1271 2106 1272 2107
rect 1332 2106 1333 2107
rect 1274 2108 1275 2109
rect 1343 2108 1344 2109
rect 1277 2110 1278 2111
rect 1325 2110 1326 2111
rect 1199 2112 1200 2113
rect 1277 2112 1278 2113
rect 1286 2112 1287 2113
rect 1307 2112 1308 2113
rect 1213 2114 1214 2115
rect 1307 2114 1308 2115
rect 1298 2116 1299 2117
rect 1356 2116 1357 2117
rect 1292 2118 1293 2119
rect 1298 2118 1299 2119
rect 1301 2118 1302 2119
rect 1313 2118 1314 2119
rect 1295 2120 1296 2121
rect 1301 2120 1302 2121
rect 1304 2120 1305 2121
rect 1316 2120 1317 2121
rect 1319 2120 1320 2121
rect 1340 2120 1341 2121
rect 1304 2122 1305 2123
rect 1339 2122 1340 2123
rect 1323 2124 1324 2125
rect 1346 2124 1347 2125
rect 1238 2126 1239 2127
rect 1346 2126 1347 2127
rect 1015 2135 1016 2136
rect 1094 2135 1095 2136
rect 1022 2137 1023 2138
rect 1079 2137 1080 2138
rect 1025 2139 1026 2140
rect 1103 2139 1104 2140
rect 1024 2141 1025 2142
rect 1034 2141 1035 2142
rect 1031 2143 1032 2144
rect 1040 2143 1041 2144
rect 1034 2145 1035 2146
rect 1106 2145 1107 2146
rect 1037 2147 1038 2148
rect 1139 2147 1140 2148
rect 1040 2149 1041 2150
rect 1133 2149 1134 2150
rect 1044 2151 1045 2152
rect 1157 2151 1158 2152
rect 1047 2153 1048 2154
rect 1089 2153 1090 2154
rect 1062 2155 1063 2156
rect 1095 2155 1096 2156
rect 1066 2157 1067 2158
rect 1163 2157 1164 2158
rect 1065 2159 1066 2160
rect 1131 2159 1132 2160
rect 1069 2161 1070 2162
rect 1098 2161 1099 2162
rect 1056 2163 1057 2164
rect 1069 2163 1070 2164
rect 1073 2163 1074 2164
rect 1121 2163 1122 2164
rect 1079 2165 1080 2166
rect 1212 2165 1213 2166
rect 1085 2167 1086 2168
rect 1169 2167 1170 2168
rect 1092 2169 1093 2170
rect 1142 2169 1143 2170
rect 1107 2171 1108 2172
rect 1127 2171 1128 2172
rect 1109 2173 1110 2174
rect 1140 2173 1141 2174
rect 1119 2175 1120 2176
rect 1166 2175 1167 2176
rect 1125 2177 1126 2178
rect 1172 2177 1173 2178
rect 1128 2179 1129 2180
rect 1175 2179 1176 2180
rect 1137 2181 1138 2182
rect 1145 2181 1146 2182
rect 1149 2181 1150 2182
rect 1196 2181 1197 2182
rect 1154 2183 1155 2184
rect 1215 2183 1216 2184
rect 1160 2185 1161 2186
rect 1253 2185 1254 2186
rect 1164 2187 1165 2188
rect 1199 2187 1200 2188
rect 1170 2189 1171 2190
rect 1205 2189 1206 2190
rect 1176 2191 1177 2192
rect 1202 2191 1203 2192
rect 1179 2193 1180 2194
rect 1190 2193 1191 2194
rect 1188 2195 1189 2196
rect 1226 2195 1227 2196
rect 1191 2197 1192 2198
rect 1223 2197 1224 2198
rect 1200 2199 1201 2200
rect 1350 2199 1351 2200
rect 1221 2201 1222 2202
rect 1298 2201 1299 2202
rect 1225 2203 1226 2204
rect 1265 2203 1266 2204
rect 1231 2205 1232 2206
rect 1271 2205 1272 2206
rect 1241 2207 1242 2208
rect 1250 2207 1251 2208
rect 1244 2209 1245 2210
rect 1274 2209 1275 2210
rect 1247 2211 1248 2212
rect 1301 2211 1302 2212
rect 1256 2213 1257 2214
rect 1310 2213 1311 2214
rect 1259 2215 1260 2216
rect 1322 2215 1323 2216
rect 1259 2217 1260 2218
rect 1280 2217 1281 2218
rect 1262 2219 1263 2220
rect 1304 2219 1305 2220
rect 1268 2221 1269 2222
rect 1329 2221 1330 2222
rect 1235 2223 1236 2224
rect 1268 2223 1269 2224
rect 1152 2225 1153 2226
rect 1234 2225 1235 2226
rect 1271 2225 1272 2226
rect 1316 2225 1317 2226
rect 1286 2227 1287 2228
rect 1339 2227 1340 2228
rect 1238 2229 1239 2230
rect 1287 2229 1288 2230
rect 1313 2229 1314 2230
rect 1343 2229 1344 2230
rect 1319 2231 1320 2232
rect 1346 2231 1347 2232
rect 1332 2233 1333 2234
rect 1336 2233 1337 2234
rect 1021 2242 1022 2243
rect 1034 2242 1035 2243
rect 1037 2242 1038 2243
rect 1056 2242 1057 2243
rect 1044 2244 1045 2245
rect 1095 2244 1096 2245
rect 1044 2246 1045 2247
rect 1047 2246 1048 2247
rect 1051 2246 1052 2247
rect 1271 2246 1272 2247
rect 1062 2248 1063 2249
rect 1066 2248 1067 2249
rect 1069 2248 1070 2249
rect 1128 2248 1129 2249
rect 1073 2250 1074 2251
rect 1083 2250 1084 2251
rect 1086 2250 1087 2251
rect 1188 2250 1189 2251
rect 1086 2252 1087 2253
rect 1089 2252 1090 2253
rect 1089 2254 1090 2255
rect 1092 2254 1093 2255
rect 1028 2256 1029 2257
rect 1092 2256 1093 2257
rect 1027 2258 1028 2259
rect 1137 2258 1138 2259
rect 1095 2260 1096 2261
rect 1098 2260 1099 2261
rect 1079 2262 1080 2263
rect 1098 2262 1099 2263
rect 1122 2262 1123 2263
rect 1212 2262 1213 2263
rect 1131 2264 1132 2265
rect 1155 2264 1156 2265
rect 1140 2266 1141 2267
rect 1158 2266 1159 2267
rect 1143 2268 1144 2269
rect 1179 2268 1180 2269
rect 1149 2270 1150 2271
rect 1173 2270 1174 2271
rect 1125 2272 1126 2273
rect 1149 2272 1150 2273
rect 1119 2274 1120 2275
rect 1125 2274 1126 2275
rect 1080 2276 1081 2277
rect 1119 2276 1120 2277
rect 1152 2276 1153 2277
rect 1225 2276 1226 2277
rect 1107 2278 1108 2279
rect 1152 2278 1153 2279
rect 1161 2278 1162 2279
rect 1164 2278 1165 2279
rect 1170 2278 1171 2279
rect 1204 2278 1205 2279
rect 1170 2280 1171 2281
rect 1176 2280 1177 2281
rect 1176 2282 1177 2283
rect 1226 2282 1227 2283
rect 1182 2284 1183 2285
rect 1215 2284 1216 2285
rect 1194 2286 1195 2287
rect 1207 2286 1208 2287
rect 1200 2288 1201 2289
rect 1284 2288 1285 2289
rect 1167 2290 1168 2291
rect 1200 2290 1201 2291
rect 1210 2290 1211 2291
rect 1247 2290 1248 2291
rect 1213 2292 1214 2293
rect 1231 2292 1232 2293
rect 1223 2294 1224 2295
rect 1250 2294 1251 2295
rect 1259 2294 1260 2295
rect 1277 2294 1278 2295
rect 1262 2296 1263 2297
rect 1280 2296 1281 2297
rect 1274 2298 1275 2299
rect 1287 2298 1288 2299
rect 1027 2307 1028 2308
rect 1149 2307 1150 2308
rect 1037 2309 1038 2310
rect 1089 2309 1090 2310
rect 1041 2311 1042 2312
rect 1092 2311 1093 2312
rect 1027 2313 1028 2314
rect 1092 2313 1093 2314
rect 1044 2315 1045 2316
rect 1125 2315 1126 2316
rect 1051 2317 1052 2318
rect 1073 2317 1074 2318
rect 1034 2319 1035 2320
rect 1074 2319 1075 2320
rect 1034 2321 1035 2322
rect 1152 2321 1153 2322
rect 1056 2323 1057 2324
rect 1076 2323 1077 2324
rect 1044 2325 1045 2326
rect 1077 2325 1078 2326
rect 1071 2327 1072 2328
rect 1086 2327 1087 2328
rect 1080 2329 1081 2330
rect 1095 2329 1096 2330
rect 1089 2331 1090 2332
rect 1113 2331 1114 2332
rect 1095 2333 1096 2334
rect 1098 2333 1099 2334
rect 1104 2333 1105 2334
rect 1155 2333 1156 2334
rect 1110 2335 1111 2336
rect 1158 2335 1159 2336
rect 1116 2337 1117 2338
rect 1179 2337 1180 2338
rect 1119 2339 1120 2340
rect 1164 2339 1165 2340
rect 1134 2341 1135 2342
rect 1167 2341 1168 2342
rect 1143 2343 1144 2344
rect 1155 2343 1156 2344
rect 1152 2345 1153 2346
rect 1170 2345 1171 2346
rect 1158 2347 1159 2348
rect 1191 2347 1192 2348
rect 1161 2349 1162 2350
rect 1197 2349 1198 2350
rect 1122 2351 1123 2352
rect 1161 2351 1162 2352
rect 1122 2353 1123 2354
rect 1170 2353 1171 2354
rect 1173 2353 1174 2354
rect 1182 2353 1183 2354
rect 1173 2355 1174 2356
rect 1176 2355 1177 2356
rect 1176 2357 1177 2358
rect 1182 2357 1183 2358
rect 1185 2357 1186 2358
rect 1213 2357 1214 2358
rect 1200 2359 1201 2360
rect 1210 2359 1211 2360
rect 1204 2361 1205 2362
rect 1216 2361 1217 2362
rect 1232 2361 1233 2362
rect 1239 2361 1240 2362
rect 1245 2361 1246 2362
rect 1252 2361 1253 2362
rect 1030 2370 1031 2371
rect 1083 2370 1084 2371
rect 1033 2372 1034 2373
rect 1074 2372 1075 2373
rect 1041 2374 1042 2375
rect 1062 2374 1063 2375
rect 1050 2376 1051 2377
rect 1071 2376 1072 2377
rect 1053 2378 1054 2379
rect 1095 2378 1096 2379
rect 1040 2380 1041 2381
rect 1095 2380 1096 2381
rect 1059 2382 1060 2383
rect 1077 2382 1078 2383
rect 1065 2384 1066 2385
rect 1155 2384 1156 2385
rect 1068 2386 1069 2387
rect 1089 2386 1090 2387
rect 1080 2388 1081 2389
rect 1086 2388 1087 2389
rect 1037 2390 1038 2391
rect 1086 2390 1087 2391
rect 1036 2392 1037 2393
rect 1077 2392 1078 2393
rect 1092 2392 1093 2393
rect 1101 2392 1102 2393
rect 1110 2392 1111 2393
rect 1188 2392 1189 2393
rect 1116 2394 1117 2395
rect 1149 2394 1150 2395
rect 1113 2396 1114 2397
rect 1116 2396 1117 2397
rect 1104 2398 1105 2399
rect 1113 2398 1114 2399
rect 1056 2400 1057 2401
rect 1104 2400 1105 2401
rect 1122 2400 1123 2401
rect 1125 2400 1126 2401
rect 1128 2400 1129 2401
rect 1134 2400 1135 2401
rect 1137 2400 1138 2401
rect 1173 2400 1174 2401
rect 1140 2402 1141 2403
rect 1158 2402 1159 2403
rect 1161 2402 1162 2403
rect 1170 2402 1171 2403
rect 1164 2404 1165 2405
rect 1167 2404 1168 2405
rect 1176 2404 1177 2405
rect 1191 2404 1192 2405
rect 1182 2406 1183 2407
rect 1185 2406 1186 2407
rect 1033 2415 1034 2416
rect 1083 2415 1084 2416
rect 1040 2417 1041 2418
rect 1062 2417 1063 2418
rect 1039 2419 1040 2420
rect 1059 2419 1060 2420
rect 1042 2421 1043 2422
rect 1089 2421 1090 2422
rect 1045 2423 1046 2424
rect 1077 2423 1078 2424
rect 1047 2425 1048 2426
rect 1104 2425 1105 2426
rect 1048 2427 1049 2428
rect 1054 2427 1055 2428
rect 1050 2429 1051 2430
rect 1101 2429 1102 2430
rect 1058 2431 1059 2432
rect 1113 2431 1114 2432
rect 1065 2433 1066 2434
rect 1116 2433 1117 2434
rect 1072 2435 1073 2436
rect 1137 2435 1138 2436
rect 1078 2437 1079 2438
rect 1128 2437 1129 2438
rect 1086 2439 1087 2440
rect 1119 2439 1120 2440
rect 1098 2441 1099 2442
rect 1131 2441 1132 2442
rect 1122 2443 1123 2444
rect 1140 2443 1141 2444
rect 1125 2445 1126 2446
rect 1146 2445 1147 2446
rect 1143 2447 1144 2448
rect 1149 2447 1150 2448
rect 1039 2456 1040 2457
rect 1061 2456 1062 2457
rect 1045 2458 1046 2459
rect 1048 2458 1049 2459
rect 1054 2458 1055 2459
rect 1072 2458 1073 2459
rect 1058 2460 1059 2461
rect 1078 2460 1079 2461
<< end >>
