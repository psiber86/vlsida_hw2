magic
tech scmos
timestamp 1395729179
<< m1p >>
use CELL  1
transform 1 0 154 0 1 102
box 0 0 6 6
use CELL  2
transform -1 0 121 0 1 66
box 0 0 6 6
use CELL  3
transform -1 0 109 0 -1 102
box 0 0 6 6
use CELL  4
transform -1 0 115 0 1 108
box 0 0 6 6
use CELL  5
transform -1 0 114 0 1 72
box 0 0 6 6
use CELL  6
transform 1 0 139 0 -1 78
box 0 0 6 6
use CELL  7
transform -1 0 124 0 1 108
box 0 0 6 6
use CELL  8
transform -1 0 159 0 1 90
box 0 0 6 6
use CELL  9
transform -1 0 141 0 -1 66
box 0 0 6 6
use CELL  10
transform 1 0 158 0 1 72
box 0 0 6 6
use CELL  11
transform -1 0 108 0 1 78
box 0 0 6 6
use CELL  12
transform 1 0 181 0 1 66
box 0 0 6 6
use CELL  13
transform -1 0 131 0 1 108
box 0 0 6 6
use CELL  14
transform -1 0 114 0 1 60
box 0 0 6 6
use CELL  15
transform -1 0 120 0 1 54
box 0 0 6 6
use CELL  16
transform -1 0 115 0 1 78
box 0 0 6 6
use CELL  17
transform 1 0 154 0 1 78
box 0 0 6 6
use CELL  18
transform 1 0 102 0 1 108
box 0 0 6 6
use CELL  19
transform 1 0 165 0 1 72
box 0 0 6 6
use CELL  20
transform -1 0 96 0 -1 96
box 0 0 6 6
use CELL  21
transform 1 0 146 0 1 84
box 0 0 6 6
use CELL  22
transform 1 0 151 0 1 72
box 0 0 6 6
use CELL  23
transform -1 0 121 0 1 72
box 0 0 6 6
use CELL  24
transform -1 0 145 0 1 78
box 0 0 6 6
use CELL  25
transform -1 0 114 0 1 102
box 0 0 6 6
use CELL  26
transform 1 0 99 0 -1 96
box 0 0 6 6
use CELL  27
transform 1 0 126 0 -1 66
box 0 0 6 6
use CELL  28
transform -1 0 180 0 1 66
box 0 0 6 6
use CELL  29
transform -1 0 121 0 1 102
box 0 0 6 6
use CELL  30
transform -1 0 158 0 -1 102
box 0 0 6 6
use CELL  31
transform -1 0 142 0 1 96
box 0 0 6 6
use CELL  32
transform -1 0 145 0 1 84
box 0 0 6 6
use CELL  33
transform -1 0 102 0 1 84
box 0 0 6 6
use CELL  34
transform -1 0 118 0 1 84
box 0 0 6 6
use CELL  35
transform 1 0 145 0 -1 102
box 0 0 6 6
use CELL  36
transform -1 0 154 0 1 78
box 0 0 6 6
use CELL  37
transform -1 0 102 0 1 96
box 0 0 6 6
use CELL  38
transform -1 0 167 0 1 102
box 0 0 6 6
use CELL  39
transform -1 0 132 0 1 90
box 0 0 6 6
use CELL  40
transform -1 0 123 0 1 90
box 0 0 6 6
use CELL  41
transform -1 0 109 0 1 84
box 0 0 6 6
use CELL  42
transform -1 0 114 0 1 66
box 0 0 6 6
use CELL  43
transform -1 0 166 0 1 66
box 0 0 6 6
use CELL  44
transform -1 0 166 0 1 90
box 0 0 6 6
use CELL  45
transform -1 0 173 0 1 66
box 0 0 6 6
<< metal1 >>
rect 171 73 172 75
rect 122 73 171 74
rect 122 73 123 82
rect 109 82 122 83
rect 107 100 108 102
rect 107 100 116 101
rect 116 91 117 100
rect 109 91 116 92
rect 100 125 101 127
rect 100 127 110 128
rect 110 118 111 127
rect 104 118 110 119
rect 165 127 166 129
rect 140 127 165 128
rect 162 134 163 136
rect 155 136 162 137
rect 100 116 101 118
rect 97 118 100 119
rect 97 109 98 118
rect 91 109 97 110
rect 140 109 141 120
rect 140 109 154 110
rect 161 116 162 118
rect 161 118 167 119
rect 167 100 168 118
rect 130 100 167 101
rect 118 116 119 118
rect 118 118 130 119
rect 119 89 120 109
rect 115 109 119 110
rect 115 109 116 127
rect 115 127 122 128
rect 122 127 123 136
rect 88 136 122 137
rect 88 91 89 136
rect 88 91 103 92
rect 122 143 123 145
rect 110 145 122 146
rect 118 55 119 57
rect 112 55 118 56
rect 161 80 162 82
rect 161 82 188 83
rect 188 64 189 82
rect 139 64 188 65
rect 149 91 150 93
rect 149 91 190 92
rect 190 53 191 91
rect 106 53 190 54
<< metal2 >>
rect 130 64 131 66
rect 122 64 130 65
rect 122 64 123 91
rect 112 91 122 92
rect 116 82 117 84
rect 100 82 116 83
rect 100 82 101 100
rect 100 100 113 101
rect 127 109 128 111
rect 106 109 127 110
rect 106 109 107 118
rect 103 118 106 119
rect 146 125 147 136
rect 129 136 146 137
rect 127 71 128 73
rect 127 73 133 74
rect 133 55 134 73
rect 112 55 133 56
rect 112 55 113 64
rect 112 64 115 65
rect 126 143 127 145
rect 116 145 126 146
rect 116 136 117 145
rect 116 136 122 137
rect 107 118 108 120
rect 107 118 110 119
rect 110 118 111 127
rect 104 127 110 128
rect 161 100 162 111
rect 149 100 161 101
rect 149 125 150 127
rect 149 127 159 128
rect 159 118 160 127
rect 156 118 159 119
rect 106 143 107 145
rect 106 145 113 146
rect 152 82 153 84
rect 149 82 152 83
rect 149 82 150 91
rect 149 91 155 92
rect 164 91 165 111
rect 164 91 172 92
rect 172 82 173 91
rect 153 82 172 83
rect 153 80 154 82
rect 134 80 153 81
rect 134 80 135 127
rect 134 127 137 128
rect 140 98 141 100
rect 137 100 140 101
rect 137 82 138 100
rect 137 82 140 83
<< end >>
