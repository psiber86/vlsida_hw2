magic
tech scmos
timestamp 1394680313
<< m1p >>
use CELL  1
transform 1 0 2668 0 1 2544
box 0 0 6 6
use CELL  2
transform -1 0 2650 0 1 2652
box 0 0 6 6
use CELL  3
transform -1 0 2630 0 1 2796
box 0 0 6 6
use CELL  4
transform -1 0 2656 0 1 2532
box 0 0 6 6
use CELL  5
transform 1 0 3056 0 1 2724
box 0 0 6 6
use CELL  6
transform -1 0 2604 0 1 2712
box 0 0 6 6
use CELL  7
transform -1 0 2840 0 1 2724
box 0 0 6 6
use CELL  8
transform -1 0 2669 0 1 2832
box 0 0 6 6
use CELL  9
transform -1 0 2595 0 1 2640
box 0 0 6 6
use CELL  10
transform -1 0 2761 0 1 2844
box 0 0 6 6
use CELL  11
transform -1 0 2789 0 1 2856
box 0 0 6 6
use CELL  12
transform -1 0 3155 0 1 2688
box 0 0 6 6
use CELL  13
transform -1 0 2598 0 1 2736
box 0 0 6 6
use CELL  14
transform -1 0 2575 0 1 2832
box 0 0 6 6
use CELL  15
transform -1 0 2962 0 1 2748
box 0 0 6 6
use CELL  16
transform -1 0 2702 0 1 2712
box 0 0 6 6
use CELL  17
transform -1 0 2690 0 -1 2538
box 0 0 6 6
use CELL  18
transform -1 0 2694 0 1 2808
box 0 0 6 6
use CELL  19
transform -1 0 2711 0 1 2532
box 0 0 6 6
use CELL  20
transform -1 0 3094 0 1 2748
box 0 0 6 6
use CELL  21
transform 1 0 2948 0 1 2736
box 0 0 6 6
use CELL  22
transform -1 0 2790 0 1 2604
box 0 0 6 6
use CELL  23
transform -1 0 2635 0 1 2748
box 0 0 6 6
use CELL  24
transform -1 0 2895 0 -1 2766
box 0 0 6 6
use CELL  25
transform -1 0 2710 0 1 2856
box 0 0 6 6
use CELL  26
transform -1 0 2556 0 1 2796
box 0 0 6 6
use CELL  27
transform -1 0 2801 0 1 2580
box 0 0 6 6
use CELL  28
transform 1 0 2941 0 1 2808
box 0 0 6 6
use CELL  29
transform -1 0 2617 0 1 2832
box 0 0 6 6
use CELL  30
transform -1 0 2545 0 1 2628
box 0 0 6 6
use CELL  31
transform -1 0 2569 0 1 2820
box 0 0 6 6
use CELL  32
transform -1 0 2928 0 1 2724
box 0 0 6 6
use CELL  33
transform -1 0 2574 0 1 2640
box 0 0 6 6
use CELL  34
transform 1 0 2586 0 1 2724
box 0 0 6 6
use CELL  35
transform 1 0 2955 0 1 2808
box 0 0 6 6
use CELL  36
transform -1 0 3230 0 -1 2658
box 0 0 6 6
use CELL  37
transform 1 0 2701 0 1 2664
box 0 0 6 6
use CELL  38
transform -1 0 2721 0 1 2664
box 0 0 6 6
use CELL  39
transform -1 0 2688 0 1 2736
box 0 0 6 6
use CELL  40
transform 1 0 3199 0 1 2628
box 0 0 6 6
use CELL  41
transform -1 0 2995 0 1 2664
box 0 0 6 6
use CELL  42
transform -1 0 2714 0 1 2616
box 0 0 6 6
use CELL  43
transform -1 0 2832 0 1 2556
box 0 0 6 6
use CELL  44
transform -1 0 2808 0 1 2544
box 0 0 6 6
use CELL  45
transform -1 0 2728 0 -1 2562
box 0 0 6 6
use CELL  46
transform 1 0 2636 0 -1 2598
box 0 0 6 6
use CELL  47
transform 1 0 2943 0 1 2772
box 0 0 6 6
use CELL  48
transform -1 0 2667 0 1 2724
box 0 0 6 6
use CELL  49
transform 1 0 2791 0 1 2772
box 0 0 6 6
use CELL  50
transform -1 0 3065 0 1 2604
box 0 0 6 6
use CELL  51
transform -1 0 3044 0 -1 2730
box 0 0 6 6
use CELL  52
transform -1 0 3249 0 -1 2646
box 0 0 6 6
use CELL  53
transform 1 0 3133 0 1 2676
box 0 0 6 6
use CELL  54
transform -1 0 2847 0 1 2796
box 0 0 6 6
use CELL  55
transform -1 0 2719 0 1 2700
box 0 0 6 6
use CELL  56
transform 1 0 2647 0 -1 2766
box 0 0 6 6
use CELL  57
transform -1 0 2797 0 1 2844
box 0 0 6 6
use CELL  58
transform -1 0 3113 0 1 2652
box 0 0 6 6
use CELL  59
transform -1 0 3124 0 -1 2634
box 0 0 6 6
use CELL  60
transform 1 0 2690 0 1 2604
box 0 0 6 6
use CELL  61
transform -1 0 3223 0 -1 2670
box 0 0 6 6
use CELL  62
transform -1 0 2771 0 1 2580
box 0 0 6 6
use CELL  63
transform 1 0 2974 0 -1 2802
box 0 0 6 6
use CELL  64
transform 1 0 3031 0 1 2592
box 0 0 6 6
use CELL  65
transform -1 0 2871 0 1 2580
box 0 0 6 6
use CELL  66
transform -1 0 2697 0 1 2532
box 0 0 6 6
use CELL  67
transform -1 0 2654 0 1 2676
box 0 0 6 6
use CELL  68
transform 1 0 3020 0 1 2748
box 0 0 6 6
use CELL  69
transform -1 0 2622 0 1 2724
box 0 0 6 6
use CELL  70
transform -1 0 2626 0 1 2784
box 0 0 6 6
use CELL  71
transform -1 0 2676 0 1 2580
box 0 0 6 6
use CELL  72
transform -1 0 2606 0 1 2700
box 0 0 6 6
use CELL  73
transform 1 0 3084 0 1 2724
box 0 0 6 6
use CELL  74
transform -1 0 2680 0 1 2616
box 0 0 6 6
use CELL  75
transform -1 0 2902 0 1 2736
box 0 0 6 6
use CELL  76
transform -1 0 2930 0 1 2784
box 0 0 6 6
use CELL  77
transform -1 0 3077 0 1 2700
box 0 0 6 6
use CELL  78
transform -1 0 2633 0 1 2616
box 0 0 6 6
use CELL  79
transform -1 0 2616 0 1 2856
box 0 0 6 6
use CELL  80
transform 1 0 3074 0 1 2664
box 0 0 6 6
use CELL  81
transform -1 0 2950 0 1 2796
box 0 0 6 6
use CELL  82
transform -1 0 3183 0 1 2664
box 0 0 6 6
use CELL  83
transform -1 0 2641 0 1 2700
box 0 0 6 6
use CELL  84
transform -1 0 2611 0 1 2712
box 0 0 6 6
use CELL  85
transform -1 0 2856 0 -1 2574
box 0 0 6 6
use CELL  86
transform -1 0 2627 0 1 2700
box 0 0 6 6
use CELL  87
transform 1 0 2905 0 -1 2598
box 0 0 6 6
use CELL  88
transform -1 0 2911 0 1 2784
box 0 0 6 6
use CELL  89
transform -1 0 2624 0 1 2832
box 0 0 6 6
use CELL  90
transform 1 0 2833 0 1 2556
box 0 0 6 6
use CELL  91
transform 1 0 3173 0 1 2688
box 0 0 6 6
use CELL  92
transform -1 0 3074 0 1 2652
box 0 0 6 6
use CELL  93
transform -1 0 2816 0 1 2556
box 0 0 6 6
use CELL  94
transform 1 0 3050 0 1 2736
box 0 0 6 6
use CELL  95
transform -1 0 2668 0 1 2640
box 0 0 6 6
use CELL  96
transform -1 0 2631 0 1 2820
box 0 0 6 6
use CELL  97
transform 1 0 3095 0 1 2748
box 0 0 6 6
use CELL  98
transform -1 0 2917 0 1 2712
box 0 0 6 6
use CELL  99
transform 1 0 2661 0 1 2808
box 0 0 6 6
use CELL  100
transform -1 0 2764 0 1 2580
box 0 0 6 6
use CELL  101
transform -1 0 2993 0 1 2712
box 0 0 6 6
use CELL  102
transform -1 0 2625 0 1 2760
box 0 0 6 6
use CELL  103
transform 1 0 2678 0 -1 2838
box 0 0 6 6
use CELL  104
transform -1 0 3085 0 1 2736
box 0 0 6 6
use CELL  105
transform 1 0 2580 0 -1 2634
box 0 0 6 6
use CELL  106
transform -1 0 2805 0 -1 2742
box 0 0 6 6
use CELL  107
transform -1 0 2726 0 1 2868
box 0 0 6 6
use CELL  108
transform -1 0 2928 0 1 2700
box 0 0 6 6
use CELL  109
transform 1 0 3025 0 1 2760
box 0 0 6 6
use CELL  110
transform -1 0 3044 0 1 2604
box 0 0 6 6
use CELL  111
transform -1 0 2730 0 1 2736
box 0 0 6 6
use CELL  112
transform -1 0 2720 0 1 2544
box 0 0 6 6
use CELL  113
transform -1 0 2720 0 1 2712
box 0 0 6 6
use CELL  114
transform -1 0 2922 0 1 2604
box 0 0 6 6
use CELL  115
transform -1 0 2637 0 1 2856
box 0 0 6 6
use CELL  116
transform 1 0 2999 0 -1 2718
box 0 0 6 6
use CELL  117
transform 1 0 2965 0 1 2772
box 0 0 6 6
use CELL  118
transform 1 0 3081 0 -1 2670
box 0 0 6 6
use CELL  119
transform -1 0 3010 0 1 2604
box 0 0 6 6
use CELL  120
transform -1 0 2756 0 1 2700
box 0 0 6 6
use CELL  121
transform 1 0 2995 0 1 2796
box 0 0 6 6
use CELL  122
transform -1 0 2907 0 1 2724
box 0 0 6 6
use CELL  123
transform -1 0 3131 0 1 2616
box 0 0 6 6
use CELL  124
transform -1 0 2668 0 1 2676
box 0 0 6 6
use CELL  125
transform -1 0 2912 0 1 2772
box 0 0 6 6
use CELL  126
transform -1 0 2628 0 1 2748
box 0 0 6 6
use CELL  127
transform 1 0 2657 0 -1 2790
box 0 0 6 6
use CELL  128
transform -1 0 2812 0 1 2736
box 0 0 6 6
use CELL  129
transform -1 0 2646 0 1 2832
box 0 0 6 6
use CELL  130
transform 1 0 3094 0 -1 2610
box 0 0 6 6
use CELL  131
transform 1 0 2617 0 1 2772
box 0 0 6 6
use CELL  132
transform -1 0 2628 0 1 2844
box 0 0 6 6
use CELL  133
transform -1 0 3107 0 1 2712
box 0 0 6 6
use CELL  134
transform -1 0 2629 0 1 2724
box 0 0 6 6
use CELL  135
transform -1 0 2939 0 1 2784
box 0 0 6 6
use CELL  136
transform -1 0 3195 0 1 2664
box 0 0 6 6
use CELL  137
transform -1 0 2796 0 1 2760
box 0 0 6 6
use CELL  138
transform -1 0 2630 0 1 2640
box 0 0 6 6
use CELL  139
transform 1 0 2649 0 -1 2634
box 0 0 6 6
use CELL  140
transform -1 0 2616 0 1 2640
box 0 0 6 6
use CELL  141
transform 1 0 3139 0 1 2616
box 0 0 6 6
use CELL  142
transform -1 0 2890 0 1 2580
box 0 0 6 6
use CELL  143
transform -1 0 2642 0 -1 2646
box 0 0 6 6
use CELL  144
transform 1 0 3139 0 1 2664
box 0 0 6 6
use CELL  145
transform -1 0 2699 0 1 2616
box 0 0 6 6
use CELL  146
transform -1 0 2974 0 1 2604
box 0 0 6 6
use CELL  147
transform -1 0 3146 0 1 2688
box 0 0 6 6
use CELL  148
transform 1 0 3115 0 1 2700
box 0 0 6 6
use CELL  149
transform -1 0 2676 0 1 2808
box 0 0 6 6
use CELL  150
transform -1 0 2653 0 1 2868
box 0 0 6 6
use CELL  151
transform 1 0 3076 0 -1 2754
box 0 0 6 6
use CELL  152
transform 1 0 2809 0 -1 2550
box 0 0 6 6
use CELL  153
transform -1 0 2790 0 1 2748
box 0 0 6 6
use CELL  154
transform -1 0 2622 0 1 2808
box 0 0 6 6
use CELL  155
transform -1 0 3138 0 1 2664
box 0 0 6 6
use CELL  156
transform 1 0 2843 0 1 2568
box 0 0 6 6
use CELL  157
transform 1 0 2977 0 1 2784
box 0 0 6 6
use CELL  158
transform -1 0 2708 0 1 2592
box 0 0 6 6
use CELL  159
transform 1 0 2580 0 -1 2766
box 0 0 6 6
use CELL  160
transform -1 0 2739 0 1 2784
box 0 0 6 6
use CELL  161
transform 1 0 2643 0 -1 2562
box 0 0 6 6
use CELL  162
transform -1 0 2672 0 1 2568
box 0 0 6 6
use CELL  163
transform -1 0 2642 0 1 2844
box 0 0 6 6
use CELL  164
transform -1 0 2623 0 1 2664
box 0 0 6 6
use CELL  165
transform 1 0 2875 0 -1 2562
box 0 0 6 6
use CELL  166
transform -1 0 2709 0 1 2724
box 0 0 6 6
use CELL  167
transform 1 0 2742 0 1 2736
box 0 0 6 6
use CELL  168
transform -1 0 2608 0 1 2724
box 0 0 6 6
use CELL  169
transform -1 0 2800 0 -1 2562
box 0 0 6 6
use CELL  170
transform -1 0 2649 0 1 2844
box 0 0 6 6
use CELL  171
transform -1 0 2712 0 1 2820
box 0 0 6 6
use CELL  172
transform 1 0 3126 0 1 2712
box 0 0 6 6
use CELL  173
transform -1 0 2770 0 1 2664
box 0 0 6 6
use CELL  174
transform -1 0 2882 0 -1 2850
box 0 0 6 6
use CELL  175
transform -1 0 3017 0 -1 2766
box 0 0 6 6
use CELL  176
transform 1 0 2694 0 -1 2838
box 0 0 6 6
use CELL  177
transform -1 0 2546 0 -1 2730
box 0 0 6 6
use CELL  178
transform 1 0 2569 0 1 2844
box 0 0 6 6
use CELL  179
transform -1 0 2845 0 -1 2850
box 0 0 6 6
use CELL  180
transform -1 0 3146 0 1 2652
box 0 0 6 6
use CELL  181
transform -1 0 2720 0 1 2592
box 0 0 6 6
use CELL  182
transform 1 0 3031 0 -1 2610
box 0 0 6 6
use CELL  183
transform -1 0 2610 0 1 2832
box 0 0 6 6
use CELL  184
transform -1 0 2727 0 1 2748
box 0 0 6 6
use CELL  185
transform -1 0 2623 0 1 2796
box 0 0 6 6
use CELL  186
transform -1 0 2667 0 1 2868
box 0 0 6 6
use CELL  187
transform -1 0 3026 0 1 2652
box 0 0 6 6
use CELL  188
transform -1 0 3078 0 1 2724
box 0 0 6 6
use CELL  189
transform -1 0 2884 0 1 2568
box 0 0 6 6
use CELL  190
transform -1 0 2759 0 1 2592
box 0 0 6 6
use CELL  191
transform 1 0 2520 0 -1 2610
box 0 0 6 6
use CELL  192
transform -1 0 2702 0 1 2556
box 0 0 6 6
use CELL  193
transform -1 0 2702 0 1 2688
box 0 0 6 6
use CELL  194
transform -1 0 3050 0 1 2712
box 0 0 6 6
use CELL  195
transform 1 0 3009 0 1 2796
box 0 0 6 6
use CELL  196
transform 1 0 3120 0 -1 2670
box 0 0 6 6
use CELL  197
transform 1 0 2853 0 -1 2610
box 0 0 6 6
use CELL  198
transform 1 0 3132 0 -1 2622
box 0 0 6 6
use CELL  199
transform -1 0 2766 0 1 2592
box 0 0 6 6
use CELL  200
transform 1 0 2993 0 1 2784
box 0 0 6 6
use CELL  201
transform -1 0 2676 0 1 2868
box 0 0 6 6
use CELL  202
transform 1 0 2626 0 1 2712
box 0 0 6 6
use CELL  203
transform -1 0 2640 0 1 2736
box 0 0 6 6
use CELL  204
transform -1 0 2826 0 1 2760
box 0 0 6 6
use CELL  205
transform -1 0 3139 0 1 2688
box 0 0 6 6
use CELL  206
transform -1 0 2749 0 1 2700
box 0 0 6 6
use CELL  207
transform -1 0 2638 0 1 2820
box 0 0 6 6
use CELL  208
transform -1 0 3255 0 -1 2646
box 0 0 6 6
use CELL  209
transform -1 0 2556 0 1 2784
box 0 0 6 6
use CELL  210
transform -1 0 2706 0 1 2868
box 0 0 6 6
use CELL  211
transform 1 0 2716 0 1 2832
box 0 0 6 6
use CELL  212
transform 1 0 3133 0 1 2712
box 0 0 6 6
use CELL  213
transform -1 0 3078 0 1 2736
box 0 0 6 6
use CELL  214
transform -1 0 2935 0 1 2700
box 0 0 6 6
use CELL  215
transform 1 0 2572 0 1 2820
box 0 0 6 6
use CELL  216
transform 1 0 2868 0 -1 2562
box 0 0 6 6
use CELL  217
transform 1 0 2728 0 -1 2718
box 0 0 6 6
use CELL  218
transform -1 0 3198 0 -1 2634
box 0 0 6 6
use CELL  219
transform 1 0 2725 0 1 2628
box 0 0 6 6
use CELL  220
transform 1 0 2902 0 1 2808
box 0 0 6 6
use CELL  221
transform -1 0 2662 0 1 2628
box 0 0 6 6
use CELL  222
transform 1 0 2607 0 1 2760
box 0 0 6 6
use CELL  223
transform -1 0 2661 0 1 2676
box 0 0 6 6
use CELL  224
transform -1 0 2553 0 1 2724
box 0 0 6 6
use CELL  225
transform -1 0 2704 0 1 2532
box 0 0 6 6
use CELL  226
transform -1 0 2641 0 1 2712
box 0 0 6 6
use CELL  227
transform -1 0 2955 0 1 2784
box 0 0 6 6
use CELL  228
transform 1 0 2948 0 1 2808
box 0 0 6 6
use CELL  229
transform 1 0 3030 0 -1 2622
box 0 0 6 6
use CELL  230
transform -1 0 3114 0 1 2700
box 0 0 6 6
use CELL  231
transform -1 0 2724 0 1 2844
box 0 0 6 6
use CELL  232
transform -1 0 2643 0 1 2628
box 0 0 6 6
use CELL  233
transform 1 0 2894 0 1 2832
box 0 0 6 6
use CELL  234
transform -1 0 2602 0 1 2676
box 0 0 6 6
use CELL  235
transform 1 0 2731 0 -1 2646
box 0 0 6 6
use CELL  236
transform -1 0 2683 0 1 2868
box 0 0 6 6
use CELL  237
transform 1 0 2622 0 -1 2562
box 0 0 6 6
use CELL  238
transform 1 0 3051 0 1 2772
box 0 0 6 6
use CELL  239
transform 1 0 2710 0 -1 2562
box 0 0 6 6
use CELL  240
transform -1 0 2695 0 1 2544
box 0 0 6 6
use CELL  241
transform -1 0 2676 0 -1 2730
box 0 0 6 6
use CELL  242
transform -1 0 2827 0 1 2772
box 0 0 6 6
use CELL  243
transform 1 0 3038 0 -1 2778
box 0 0 6 6
use CELL  244
transform -1 0 2693 0 -1 2838
box 0 0 6 6
use CELL  245
transform 1 0 2984 0 1 2592
box 0 0 6 6
use CELL  246
transform -1 0 2655 0 1 2616
box 0 0 6 6
use CELL  247
transform 1 0 2956 0 1 2784
box 0 0 6 6
use CELL  248
transform -1 0 2875 0 1 2832
box 0 0 6 6
use CELL  249
transform -1 0 2626 0 1 2736
box 0 0 6 6
use CELL  250
transform 1 0 2654 0 -1 2874
box 0 0 6 6
use CELL  251
transform 1 0 2818 0 1 2856
box 0 0 6 6
use CELL  252
transform 1 0 3237 0 -1 2658
box 0 0 6 6
use CELL  253
transform -1 0 3237 0 1 2652
box 0 0 6 6
use CELL  254
transform 1 0 3088 0 -1 2694
box 0 0 6 6
use CELL  255
transform 1 0 3006 0 1 2784
box 0 0 6 6
use CELL  256
transform -1 0 2613 0 1 2700
box 0 0 6 6
use CELL  257
transform 1 0 2804 0 -1 2862
box 0 0 6 6
use CELL  258
transform 1 0 2675 0 -1 2562
box 0 0 6 6
use CELL  259
transform -1 0 2669 0 1 2880
box 0 0 6 6
use CELL  260
transform -1 0 3116 0 1 2640
box 0 0 6 6
use CELL  261
transform -1 0 2677 0 1 2712
box 0 0 6 6
use CELL  262
transform 1 0 2806 0 1 2568
box 0 0 6 6
use CELL  263
transform -1 0 2742 0 1 2748
box 0 0 6 6
use CELL  264
transform -1 0 2693 0 1 2640
box 0 0 6 6
use CELL  265
transform 1 0 2963 0 -1 2754
box 0 0 6 6
use CELL  266
transform -1 0 3051 0 1 2592
box 0 0 6 6
use CELL  267
transform 1 0 2746 0 1 2724
box 0 0 6 6
use CELL  268
transform -1 0 2644 0 1 2856
box 0 0 6 6
use CELL  269
transform -1 0 2659 0 1 2664
box 0 0 6 6
use CELL  270
transform -1 0 2984 0 1 2736
box 0 0 6 6
use CELL  271
transform 1 0 2646 0 1 2820
box 0 0 6 6
use CELL  272
transform -1 0 2610 0 1 2628
box 0 0 6 6
use CELL  273
transform -1 0 2604 0 1 2652
box 0 0 6 6
use CELL  274
transform -1 0 2655 0 1 2736
box 0 0 6 6
use CELL  275
transform -1 0 2989 0 1 2760
box 0 0 6 6
use CELL  276
transform -1 0 3054 0 1 2760
box 0 0 6 6
use CELL  277
transform 1 0 2655 0 1 2592
box 0 0 6 6
use CELL  278
transform 1 0 2769 0 1 2784
box 0 0 6 6
use CELL  279
transform -1 0 2648 0 1 2880
box 0 0 6 6
use CELL  280
transform -1 0 2835 0 1 2808
box 0 0 6 6
use CELL  281
transform 1 0 2930 0 1 2712
box 0 0 6 6
use CELL  282
transform 1 0 2647 0 -1 2838
box 0 0 6 6
use CELL  283
transform -1 0 3059 0 1 2700
box 0 0 6 6
use CELL  284
transform -1 0 2642 0 -1 2574
box 0 0 6 6
use CELL  285
transform 1 0 3083 0 1 2640
box 0 0 6 6
use CELL  286
transform -1 0 2615 0 1 2724
box 0 0 6 6
use CELL  287
transform -1 0 2811 0 1 2784
box 0 0 6 6
use CELL  288
transform 1 0 2643 0 -1 2538
box 0 0 6 6
use CELL  289
transform -1 0 3030 0 1 2592
box 0 0 6 6
use CELL  290
transform 1 0 3043 0 1 2736
box 0 0 6 6
use CELL  291
transform -1 0 2689 0 1 2676
box 0 0 6 6
use CELL  292
transform 1 0 3003 0 1 2592
box 0 0 6 6
use CELL  293
transform 1 0 2877 0 1 2580
box 0 0 6 6
use CELL  294
transform 1 0 3045 0 1 2772
box 0 0 6 6
use CELL  295
transform 1 0 2859 0 -1 2826
box 0 0 6 6
use CELL  296
transform 1 0 2860 0 1 2844
box 0 0 6 6
use CELL  297
transform 1 0 2857 0 1 2832
box 0 0 6 6
use CELL  298
transform -1 0 3022 0 -1 2778
box 0 0 6 6
use CELL  299
transform -1 0 2904 0 1 2592
box 0 0 6 6
use CELL  300
transform 1 0 3210 0 -1 2658
box 0 0 6 6
use CELL  301
transform -1 0 2877 0 1 2820
box 0 0 6 6
use CELL  302
transform 1 0 2734 0 -1 2562
box 0 0 6 6
use CELL  303
transform -1 0 2651 0 1 2856
box 0 0 6 6
use CELL  304
transform -1 0 3209 0 1 2664
box 0 0 6 6
use CELL  305
transform 1 0 2940 0 1 2784
box 0 0 6 6
use CELL  306
transform 1 0 2950 0 1 2820
box 0 0 6 6
use CELL  307
transform -1 0 2649 0 1 2772
box 0 0 6 6
use CELL  308
transform -1 0 2728 0 1 2664
box 0 0 6 6
use CELL  309
transform -1 0 2616 0 1 2580
box 0 0 6 6
use CELL  310
transform -1 0 2720 0 1 2784
box 0 0 6 6
use CELL  311
transform -1 0 3262 0 -1 2646
box 0 0 6 6
use CELL  312
transform 1 0 2586 0 1 2700
box 0 0 6 6
use CELL  313
transform -1 0 2721 0 1 2616
box 0 0 6 6
use CELL  314
transform -1 0 2691 0 1 2568
box 0 0 6 6
use CELL  315
transform -1 0 2717 0 1 2796
box 0 0 6 6
use CELL  316
transform 1 0 2918 0 1 2712
box 0 0 6 6
use CELL  317
transform -1 0 3086 0 1 2604
box 0 0 6 6
use CELL  318
transform 1 0 3153 0 -1 2622
box 0 0 6 6
use CELL  319
transform -1 0 2838 0 1 2592
box 0 0 6 6
use CELL  320
transform -1 0 2695 0 -1 2670
box 0 0 6 6
use CELL  321
transform -1 0 2660 0 1 2544
box 0 0 6 6
use CELL  322
transform 1 0 2822 0 1 2568
box 0 0 6 6
use CELL  323
transform -1 0 2616 0 1 2796
box 0 0 6 6
use CELL  324
transform 1 0 2776 0 -1 2862
box 0 0 6 6
use CELL  325
transform -1 0 3041 0 1 2676
box 0 0 6 6
use CELL  326
transform -1 0 2623 0 1 2592
box 0 0 6 6
use CELL  327
transform 1 0 3031 0 -1 2730
box 0 0 6 6
use CELL  328
transform 1 0 3210 0 1 2664
box 0 0 6 6
use CELL  329
transform -1 0 2648 0 1 2700
box 0 0 6 6
use CELL  330
transform -1 0 2599 0 1 2760
box 0 0 6 6
use CELL  331
transform -1 0 2688 0 1 2544
box 0 0 6 6
use CELL  332
transform -1 0 3088 0 1 2748
box 0 0 6 6
use CELL  333
transform -1 0 2688 0 1 2688
box 0 0 6 6
use CELL  334
transform -1 0 2673 0 1 2700
box 0 0 6 6
use CELL  335
transform 1 0 2864 0 1 2568
box 0 0 6 6
use CELL  336
transform -1 0 2623 0 1 2676
box 0 0 6 6
use CELL  337
transform -1 0 2956 0 1 2604
box 0 0 6 6
use CELL  338
transform -1 0 2767 0 -1 2550
box 0 0 6 6
use CELL  339
transform -1 0 2846 0 -1 2562
box 0 0 6 6
use CELL  340
transform -1 0 2903 0 1 2568
box 0 0 6 6
use CELL  341
transform 1 0 2661 0 1 2772
box 0 0 6 6
use CELL  342
transform 1 0 2941 0 1 2736
box 0 0 6 6
use CELL  343
transform -1 0 2562 0 1 2820
box 0 0 6 6
use CELL  344
transform -1 0 2929 0 1 2736
box 0 0 6 6
use CELL  345
transform 1 0 3117 0 1 2676
box 0 0 6 6
use CELL  346
transform -1 0 2610 0 1 2808
box 0 0 6 6
use CELL  347
transform 1 0 3004 0 1 2736
box 0 0 6 6
use CELL  348
transform -1 0 3216 0 -1 2646
box 0 0 6 6
use CELL  349
transform 1 0 2647 0 1 2580
box 0 0 6 6
use CELL  350
transform -1 0 2533 0 1 2604
box 0 0 6 6
use CELL  351
transform 1 0 2589 0 -1 2670
box 0 0 6 6
use CELL  352
transform -1 0 2647 0 1 2784
box 0 0 6 6
use CELL  353
transform -1 0 3123 0 1 2712
box 0 0 6 6
use CELL  354
transform 1 0 3236 0 1 2640
box 0 0 6 6
use CELL  355
transform -1 0 2785 0 1 2712
box 0 0 6 6
use CELL  356
transform -1 0 2822 0 1 2676
box 0 0 6 6
use CELL  357
transform -1 0 3116 0 1 2712
box 0 0 6 6
use CELL  358
transform 1 0 2775 0 1 2544
box 0 0 6 6
use CELL  359
transform -1 0 3033 0 -1 2754
box 0 0 6 6
use CELL  360
transform -1 0 3044 0 1 2592
box 0 0 6 6
use CELL  361
transform -1 0 2955 0 1 2760
box 0 0 6 6
use CELL  362
transform 1 0 2856 0 -1 2586
box 0 0 6 6
use CELL  363
transform -1 0 2704 0 1 2580
box 0 0 6 6
use CELL  364
transform 1 0 2724 0 1 2640
box 0 0 6 6
use CELL  365
transform 1 0 2986 0 1 2604
box 0 0 6 6
use CELL  366
transform 1 0 3062 0 1 2748
box 0 0 6 6
use CELL  367
transform -1 0 2702 0 1 2784
box 0 0 6 6
use CELL  368
transform 1 0 3041 0 1 2760
box 0 0 6 6
use CELL  369
transform 1 0 3064 0 1 2688
box 0 0 6 6
use CELL  370
transform -1 0 2812 0 1 2664
box 0 0 6 6
use CELL  371
transform -1 0 3134 0 1 2640
box 0 0 6 6
use CELL  372
transform 1 0 2981 0 1 2796
box 0 0 6 6
use CELL  373
transform 1 0 2669 0 -1 2850
box 0 0 6 6
use CELL  374
transform -1 0 2666 0 1 2700
box 0 0 6 6
use CELL  375
transform -1 0 2640 0 1 2784
box 0 0 6 6
use CELL  376
transform -1 0 2873 0 1 2844
box 0 0 6 6
use CELL  377
transform 1 0 2626 0 -1 2658
box 0 0 6 6
use CELL  378
transform -1 0 3197 0 1 2652
box 0 0 6 6
use CELL  379
transform -1 0 3160 0 1 2676
box 0 0 6 6
use CELL  380
transform -1 0 2612 0 1 2688
box 0 0 6 6
use CELL  381
transform 1 0 2718 0 1 2760
box 0 0 6 6
use CELL  382
transform -1 0 3043 0 1 2616
box 0 0 6 6
use CELL  383
transform -1 0 2643 0 1 2808
box 0 0 6 6
use CELL  384
transform 1 0 2748 0 -1 2622
box 0 0 6 6
use CELL  385
transform -1 0 2633 0 1 2736
box 0 0 6 6
use CELL  386
transform -1 0 2755 0 1 2640
box 0 0 6 6
use CELL  387
transform -1 0 3037 0 1 2736
box 0 0 6 6
use CELL  388
transform -1 0 2748 0 1 2604
box 0 0 6 6
use CELL  389
transform -1 0 3029 0 1 2772
box 0 0 6 6
use CELL  390
transform 1 0 2640 0 1 2544
box 0 0 6 6
use CELL  391
transform -1 0 2717 0 1 2760
box 0 0 6 6
use CELL  392
transform 1 0 2605 0 -1 2550
box 0 0 6 6
use CELL  393
transform -1 0 2619 0 1 2736
box 0 0 6 6
use CELL  394
transform 1 0 2745 0 1 2856
box 0 0 6 6
use CELL  395
transform -1 0 2740 0 1 2832
box 0 0 6 6
use CELL  396
transform -1 0 2611 0 1 2652
box 0 0 6 6
use CELL  397
transform 1 0 2950 0 -1 2778
box 0 0 6 6
use CELL  398
transform -1 0 2974 0 1 2808
box 0 0 6 6
use CELL  399
transform 1 0 2943 0 1 2820
box 0 0 6 6
use CELL  400
transform -1 0 2628 0 -1 2874
box 0 0 6 6
use CELL  401
transform 1 0 2957 0 1 2820
box 0 0 6 6
use CELL  402
transform -1 0 2598 0 1 2616
box 0 0 6 6
use CELL  403
transform -1 0 2629 0 1 2808
box 0 0 6 6
use CELL  404
transform -1 0 3106 0 1 2688
box 0 0 6 6
use CELL  405
transform -1 0 2675 0 1 2676
box 0 0 6 6
use CELL  406
transform 1 0 2705 0 -1 2550
box 0 0 6 6
use CELL  407
transform 1 0 2997 0 -1 2622
box 0 0 6 6
use CELL  408
transform 1 0 2624 0 1 2832
box 0 0 6 6
use CELL  409
transform 1 0 3017 0 1 2592
box 0 0 6 6
use CELL  410
transform -1 0 3219 0 1 2628
box 0 0 6 6
use CELL  411
transform -1 0 2623 0 1 2580
box 0 0 6 6
use CELL  412
transform -1 0 2646 0 1 2760
box 0 0 6 6
use CELL  413
transform -1 0 2644 0 1 2796
box 0 0 6 6
use CELL  414
transform -1 0 2777 0 1 2652
box 0 0 6 6
use CELL  415
transform 1 0 2794 0 -1 2694
box 0 0 6 6
use CELL  416
transform 1 0 2934 0 1 2604
box 0 0 6 6
use CELL  417
transform 1 0 2891 0 1 2580
box 0 0 6 6
use CELL  418
transform -1 0 2788 0 -1 2550
box 0 0 6 6
use CELL  419
transform -1 0 2807 0 1 2556
box 0 0 6 6
use CELL  420
transform -1 0 2896 0 -1 2574
box 0 0 6 6
use CELL  421
transform -1 0 2965 0 1 2592
box 0 0 6 6
use CELL  422
transform -1 0 2634 0 1 2700
box 0 0 6 6
use CELL  423
transform -1 0 3038 0 1 2772
box 0 0 6 6
use CELL  424
transform 1 0 2821 0 1 2712
box 0 0 6 6
use CELL  425
transform -1 0 2662 0 1 2604
box 0 0 6 6
use CELL  426
transform -1 0 3202 0 1 2664
box 0 0 6 6
use CELL  427
transform -1 0 2617 0 1 2628
box 0 0 6 6
use CELL  428
transform -1 0 2911 0 1 2580
box 0 0 6 6
use CELL  429
transform 1 0 2690 0 -1 2598
box 0 0 6 6
use CELL  430
transform 1 0 3065 0 1 2640
box 0 0 6 6
use CELL  431
transform 1 0 2683 0 -1 2598
box 0 0 6 6
use CELL  432
transform 1 0 2514 0 -1 2754
box 0 0 6 6
use CELL  433
transform 1 0 2849 0 1 2772
box 0 0 6 6
use CELL  434
transform -1 0 3003 0 1 2760
box 0 0 6 6
use CELL  435
transform -1 0 2693 0 1 2652
box 0 0 6 6
use CELL  436
transform -1 0 3084 0 1 2628
box 0 0 6 6
use CELL  437
transform -1 0 2802 0 1 2748
box 0 0 6 6
use CELL  438
transform 1 0 3022 0 1 2604
box 0 0 6 6
use CELL  439
transform 1 0 2868 0 1 2700
box 0 0 6 6
use CELL  440
transform -1 0 2669 0 1 2652
box 0 0 6 6
use CELL  441
transform 1 0 2838 0 1 2760
box 0 0 6 6
use CELL  442
transform 1 0 3004 0 -1 2766
box 0 0 6 6
use CELL  443
transform -1 0 2623 0 1 2856
box 0 0 6 6
use CELL  444
transform -1 0 2774 0 1 2628
box 0 0 6 6
use CELL  445
transform -1 0 2658 0 1 2856
box 0 0 6 6
use CELL  446
transform 1 0 2851 0 1 2844
box 0 0 6 6
use CELL  447
transform 1 0 2575 0 1 2640
box 0 0 6 6
use CELL  448
transform -1 0 3149 0 1 2640
box 0 0 6 6
use CELL  449
transform -1 0 3209 0 1 2652
box 0 0 6 6
use CELL  450
transform -1 0 2655 0 1 2880
box 0 0 6 6
use CELL  451
transform 1 0 2883 0 1 2820
box 0 0 6 6
use CELL  452
transform 1 0 2847 0 -1 2562
box 0 0 6 6
use CELL  453
transform -1 0 3193 0 -1 2694
box 0 0 6 6
use CELL  454
transform -1 0 3086 0 -1 2718
box 0 0 6 6
use CELL  455
transform 1 0 2791 0 1 2832
box 0 0 6 6
use CELL  456
transform -1 0 2713 0 1 2676
box 0 0 6 6
use CELL  457
transform -1 0 2745 0 1 2724
box 0 0 6 6
use CELL  458
transform -1 0 2725 0 -1 2538
box 0 0 6 6
use CELL  459
transform -1 0 2642 0 -1 2754
box 0 0 6 6
use CELL  460
transform -1 0 2612 0 1 2736
box 0 0 6 6
use CELL  461
transform -1 0 3002 0 1 2592
box 0 0 6 6
use CELL  462
transform -1 0 2841 0 1 2820
box 0 0 6 6
use CELL  463
transform -1 0 2702 0 1 2544
box 0 0 6 6
use CELL  464
transform 1 0 2702 0 1 2808
box 0 0 6 6
use CELL  465
transform -1 0 2938 0 1 2796
box 0 0 6 6
use CELL  466
transform 1 0 2995 0 -1 2730
box 0 0 6 6
use CELL  467
transform 1 0 3098 0 -1 2742
box 0 0 6 6
use CELL  468
transform -1 0 2687 0 1 2700
box 0 0 6 6
use CELL  469
transform 1 0 2904 0 1 2844
box 0 0 6 6
use CELL  470
transform 1 0 3167 0 1 2628
box 0 0 6 6
use CELL  471
transform -1 0 2793 0 1 2688
box 0 0 6 6
use CELL  472
transform -1 0 2694 0 1 2700
box 0 0 6 6
use CELL  473
transform 1 0 2897 0 1 2844
box 0 0 6 6
use CELL  474
transform 1 0 2654 0 1 2580
box 0 0 6 6
use CELL  475
transform 1 0 2716 0 1 2580
box 0 0 6 6
use CELL  476
transform 1 0 2888 0 -1 2646
box 0 0 6 6
use CELL  477
transform -1 0 3117 0 1 2736
box 0 0 6 6
use CELL  478
transform 1 0 2521 0 1 2556
box 0 0 6 6
use CELL  479
transform 1 0 3066 0 1 2604
box 0 0 6 6
use CELL  480
transform -1 0 2639 0 1 2760
box 0 0 6 6
use CELL  481
transform -1 0 2692 0 1 2616
box 0 0 6 6
use CELL  482
transform -1 0 2636 0 1 2724
box 0 0 6 6
use CELL  483
transform 1 0 2842 0 -1 2778
box 0 0 6 6
use CELL  484
transform -1 0 2905 0 1 2820
box 0 0 6 6
use CELL  485
transform -1 0 2624 0 1 2604
box 0 0 6 6
use CELL  486
transform -1 0 2618 0 1 2652
box 0 0 6 6
use CELL  487
transform -1 0 2672 0 1 2856
box 0 0 6 6
use CELL  488
transform -1 0 2618 0 1 2712
box 0 0 6 6
use CELL  489
transform -1 0 2738 0 1 2688
box 0 0 6 6
use CELL  490
transform 1 0 2631 0 -1 2586
box 0 0 6 6
use CELL  491
transform -1 0 2660 0 1 2724
box 0 0 6 6
use CELL  492
transform -1 0 3077 0 1 2628
box 0 0 6 6
use CELL  493
transform -1 0 2665 0 -1 2718
box 0 0 6 6
use CELL  494
transform 1 0 3184 0 -1 2658
box 0 0 6 6
use CELL  495
transform 1 0 2817 0 1 2556
box 0 0 6 6
use CELL  496
transform 1 0 2727 0 1 2568
box 0 0 6 6
use CELL  497
transform -1 0 2967 0 1 2724
box 0 0 6 6
use CELL  498
transform -1 0 3186 0 1 2688
box 0 0 6 6
use CELL  499
transform -1 0 2975 0 1 2628
box 0 0 6 6
use CELL  500
transform -1 0 3105 0 1 2664
box 0 0 6 6
use CELL  501
transform 1 0 2649 0 1 2808
box 0 0 6 6
use CELL  502
transform 1 0 2816 0 1 2544
box 0 0 6 6
use CELL  503
transform 1 0 3223 0 1 2664
box 0 0 6 6
use CELL  504
transform -1 0 3226 0 -1 2634
box 0 0 6 6
use CELL  505
transform 1 0 2915 0 1 2820
box 0 0 6 6
use CELL  506
transform -1 0 3008 0 1 2772
box 0 0 6 6
use CELL  507
transform -1 0 2661 0 1 2748
box 0 0 6 6
use CELL  508
transform -1 0 2698 0 -1 2634
box 0 0 6 6
use CELL  509
transform -1 0 3121 0 -1 2694
box 0 0 6 6
use CELL  510
transform 1 0 3146 0 1 2616
box 0 0 6 6
use CELL  511
transform -1 0 2980 0 1 2772
box 0 0 6 6
use CELL  512
transform 1 0 2625 0 1 2628
box 0 0 6 6
use CELL  513
transform 1 0 3002 0 1 2796
box 0 0 6 6
use CELL  514
transform -1 0 2626 0 1 2616
box 0 0 6 6
use CELL  515
transform -1 0 2662 0 1 2688
box 0 0 6 6
use CELL  516
transform 1 0 3227 0 -1 2634
box 0 0 6 6
use CELL  517
transform 1 0 2922 0 1 2820
box 0 0 6 6
use CELL  518
transform 1 0 3163 0 1 2664
box 0 0 6 6
use CELL  519
transform -1 0 2601 0 1 2724
box 0 0 6 6
use CELL  520
transform -1 0 2660 0 1 2796
box 0 0 6 6
use CELL  521
transform -1 0 3153 0 1 2676
box 0 0 6 6
use CELL  522
transform -1 0 3106 0 1 2616
box 0 0 6 6
use CELL  523
transform -1 0 2681 0 1 2688
box 0 0 6 6
use CELL  524
transform 1 0 2845 0 1 2748
box 0 0 6 6
use CELL  525
transform -1 0 2717 0 1 2844
box 0 0 6 6
use CELL  526
transform -1 0 2919 0 1 2760
box 0 0 6 6
use CELL  527
transform 1 0 2603 0 -1 2682
box 0 0 6 6
use CELL  528
transform 1 0 2849 0 -1 2586
box 0 0 6 6
use CELL  529
transform -1 0 3082 0 1 2616
box 0 0 6 6
use CELL  530
transform -1 0 3017 0 1 2748
box 0 0 6 6
use CELL  531
transform -1 0 2611 0 1 2820
box 0 0 6 6
use CELL  532
transform -1 0 3071 0 1 2724
box 0 0 6 6
use CELL  533
transform -1 0 3146 0 1 2676
box 0 0 6 6
use CELL  534
transform 1 0 2695 0 -1 2706
box 0 0 6 6
use CELL  535
transform -1 0 2633 0 1 2784
box 0 0 6 6
use CELL  536
transform 1 0 2936 0 1 2820
box 0 0 6 6
use CELL  537
transform -1 0 2701 0 1 2808
box 0 0 6 6
use CELL  538
transform 1 0 2557 0 1 2796
box 0 0 6 6
use CELL  539
transform -1 0 2690 0 1 2796
box 0 0 6 6
use CELL  540
transform -1 0 2602 0 1 2640
box 0 0 6 6
use CELL  541
transform 1 0 3026 0 1 2676
box 0 0 6 6
use CELL  542
transform 1 0 2643 0 1 2568
box 0 0 6 6
use CELL  543
transform -1 0 2740 0 1 2616
box 0 0 6 6
use CELL  544
transform 1 0 2650 0 1 2568
box 0 0 6 6
use CELL  545
transform 1 0 2721 0 1 2544
box 0 0 6 6
use CELL  546
transform -1 0 2625 0 -1 2718
box 0 0 6 6
use CELL  547
transform -1 0 2623 0 1 2640
box 0 0 6 6
use CELL  548
transform 1 0 2718 0 1 2628
box 0 0 6 6
use CELL  549
transform -1 0 2994 0 1 2724
box 0 0 6 6
use CELL  550
transform -1 0 2820 0 1 2784
box 0 0 6 6
use CELL  551
transform -1 0 2981 0 -1 2754
box 0 0 6 6
use CELL  552
transform -1 0 2681 0 1 2796
box 0 0 6 6
use CELL  553
transform 1 0 2604 0 -1 2610
box 0 0 6 6
use CELL  554
transform 1 0 2783 0 1 2700
box 0 0 6 6
use CELL  555
transform -1 0 2595 0 1 2676
box 0 0 6 6
use CELL  556
transform 1 0 3018 0 1 2760
box 0 0 6 6
use CELL  557
transform -1 0 2844 0 1 2748
box 0 0 6 6
use CELL  558
transform -1 0 2823 0 1 2820
box 0 0 6 6
use CELL  559
transform 1 0 2629 0 1 2556
box 0 0 6 6
use CELL  560
transform -1 0 3038 0 1 2712
box 0 0 6 6
use CELL  561
transform 1 0 3116 0 1 2652
box 0 0 6 6
use CELL  562
transform 1 0 2736 0 -1 2850
box 0 0 6 6
use CELL  563
transform -1 0 2722 0 1 2856
box 0 0 6 6
use CELL  564
transform -1 0 2865 0 1 2808
box 0 0 6 6
use CELL  565
transform -1 0 2685 0 1 2580
box 0 0 6 6
use CELL  566
transform 1 0 2533 0 1 2724
box 0 0 6 6
use CELL  567
transform -1 0 2664 0 1 2736
box 0 0 6 6
use CELL  568
transform 1 0 2726 0 1 2784
box 0 0 6 6
use CELL  569
transform -1 0 3068 0 1 2676
box 0 0 6 6
use CELL  570
transform -1 0 3038 0 1 2760
box 0 0 6 6
use CELL  571
transform -1 0 2817 0 1 2856
box 0 0 6 6
use CELL  572
transform -1 0 2733 0 1 2616
box 0 0 6 6
use CELL  573
transform -1 0 2940 0 1 2808
box 0 0 6 6
use CELL  574
transform -1 0 2858 0 1 2724
box 0 0 6 6
use CELL  575
transform 1 0 3101 0 1 2700
box 0 0 6 6
use CELL  576
transform -1 0 3117 0 1 2628
box 0 0 6 6
use CELL  577
transform -1 0 2604 0 1 2544
box 0 0 6 6
use CELL  578
transform -1 0 2641 0 1 2880
box 0 0 6 6
use CELL  579
transform 1 0 2885 0 -1 2838
box 0 0 6 6
use CELL  580
transform 1 0 2671 0 1 2520
box 0 0 6 6
use CELL  581
transform 1 0 2756 0 1 2640
box 0 0 6 6
use CELL  582
transform 1 0 3206 0 -1 2634
box 0 0 6 6
use CELL  583
transform -1 0 2699 0 1 2868
box 0 0 6 6
use CELL  584
transform -1 0 2767 0 1 2832
box 0 0 6 6
use CELL  585
transform -1 0 3130 0 1 2676
box 0 0 6 6
use CELL  586
transform -1 0 2692 0 1 2868
box 0 0 6 6
use CELL  587
transform -1 0 2663 0 1 2844
box 0 0 6 6
use CELL  588
transform 1 0 3069 0 1 2748
box 0 0 6 6
use CELL  589
transform -1 0 2752 0 1 2652
box 0 0 6 6
use CELL  590
transform 1 0 2629 0 -1 2574
box 0 0 6 6
use CELL  591
transform -1 0 3090 0 1 2676
box 0 0 6 6
use CELL  592
transform -1 0 2901 0 1 2808
box 0 0 6 6
use CELL  593
transform 1 0 3107 0 -1 2622
box 0 0 6 6
use CELL  594
transform -1 0 2737 0 -1 2862
box 0 0 6 6
use CELL  595
transform 1 0 2917 0 1 2592
box 0 0 6 6
use CELL  596
transform -1 0 2900 0 1 2652
box 0 0 6 6
use CELL  597
transform 1 0 2618 0 1 2544
box 0 0 6 6
use CELL  598
transform -1 0 2759 0 1 2724
box 0 0 6 6
use CELL  599
transform -1 0 2750 0 1 2688
box 0 0 6 6
use CELL  600
transform -1 0 2631 0 1 2604
box 0 0 6 6
use CELL  601
transform -1 0 3223 0 1 2652
box 0 0 6 6
use CELL  602
transform -1 0 2944 0 1 2580
box 0 0 6 6
use CELL  603
transform -1 0 2759 0 1 2652
box 0 0 6 6
use CELL  604
transform -1 0 2647 0 1 2664
box 0 0 6 6
use CELL  605
transform -1 0 2687 0 1 2844
box 0 0 6 6
use CELL  606
transform 1 0 3094 0 1 2712
box 0 0 6 6
use CELL  607
transform -1 0 2796 0 -1 2862
box 0 0 6 6
use CELL  608
transform -1 0 2767 0 -1 2634
box 0 0 6 6
use CELL  609
transform -1 0 2631 0 1 2688
box 0 0 6 6
use CELL  610
transform -1 0 2728 0 1 2652
box 0 0 6 6
use CELL  611
transform -1 0 2605 0 1 2748
box 0 0 6 6
use CELL  612
transform -1 0 2980 0 1 2760
box 0 0 6 6
use CELL  613
transform -1 0 2904 0 -1 2790
box 0 0 6 6
use CELL  614
transform -1 0 2725 0 1 2676
box 0 0 6 6
use CELL  615
transform -1 0 2819 0 1 2568
box 0 0 6 6
use CELL  616
transform 1 0 2929 0 1 2820
box 0 0 6 6
use CELL  617
transform -1 0 2667 0 1 2820
box 0 0 6 6
use CELL  618
transform -1 0 2679 0 1 2568
box 0 0 6 6
use CELL  619
transform -1 0 2582 0 1 2844
box 0 0 6 6
use CELL  620
transform -1 0 2634 0 1 2880
box 0 0 6 6
use CELL  621
transform -1 0 2642 0 1 2676
box 0 0 6 6
use CELL  622
transform -1 0 2718 0 1 2532
box 0 0 6 6
use CELL  623
transform -1 0 2635 0 1 2868
box 0 0 6 6
use CELL  624
transform -1 0 2662 0 -1 2886
box 0 0 6 6
use CELL  625
transform -1 0 2520 0 1 2556
box 0 0 6 6
use CELL  626
transform -1 0 2670 0 1 2532
box 0 0 6 6
use CELL  627
transform -1 0 2747 0 1 2616
box 0 0 6 6
use CELL  628
transform -1 0 2669 0 1 2580
box 0 0 6 6
use CELL  629
transform -1 0 2609 0 1 2640
box 0 0 6 6
use CELL  630
transform 1 0 2528 0 1 2748
box 0 0 6 6
use CELL  631
transform 1 0 2762 0 1 2676
box 0 0 6 6
use CELL  632
transform -1 0 2619 0 1 2688
box 0 0 6 6
use CELL  633
transform -1 0 2630 0 1 2592
box 0 0 6 6
use CELL  634
transform -1 0 2538 0 1 2628
box 0 0 6 6
use CELL  635
transform -1 0 2851 0 1 2832
box 0 0 6 6
use CELL  636
transform -1 0 2698 0 1 2568
box 0 0 6 6
use CELL  637
transform -1 0 2646 0 1 2520
box 0 0 6 6
use CELL  638
transform 1 0 2932 0 1 2592
box 0 0 6 6
use CELL  639
transform -1 0 2663 0 1 2532
box 0 0 6 6
use CELL  640
transform -1 0 2592 0 -1 2718
box 0 0 6 6
use CELL  641
transform -1 0 2605 0 1 2736
box 0 0 6 6
use CELL  642
transform 1 0 2908 0 1 2832
box 0 0 6 6
use CELL  643
transform -1 0 2931 0 1 2796
box 0 0 6 6
use CELL  644
transform 1 0 2966 0 -1 2598
box 0 0 6 6
use CELL  645
transform -1 0 2710 0 1 2568
box 0 0 6 6
use CELL  646
transform -1 0 2882 0 1 2832
box 0 0 6 6
use CELL  647
transform -1 0 2689 0 -1 2610
box 0 0 6 6
use CELL  648
transform -1 0 2619 0 1 2616
box 0 0 6 6
use CELL  649
transform -1 0 2675 0 1 2640
box 0 0 6 6
use CELL  650
transform -1 0 2722 0 1 2772
box 0 0 6 6
use CELL  651
transform -1 0 2657 0 1 2652
box 0 0 6 6
use CELL  652
transform 1 0 3122 0 -1 2706
box 0 0 6 6
use CELL  653
transform -1 0 2774 0 1 2544
box 0 0 6 6
use CELL  654
transform -1 0 3228 0 1 2640
box 0 0 6 6
use CELL  655
transform -1 0 2680 0 1 2700
box 0 0 6 6
use CELL  656
transform -1 0 2695 0 1 2688
box 0 0 6 6
use CELL  657
transform 1 0 2918 0 1 2808
box 0 0 6 6
use CELL  658
transform -1 0 2662 0 1 2832
box 0 0 6 6
use CELL  659
transform 1 0 2965 0 -1 2802
box 0 0 6 6
use CELL  660
transform 1 0 2737 0 1 2676
box 0 0 6 6
use CELL  661
transform -1 0 2624 0 1 2628
box 0 0 6 6
use CELL  662
transform 1 0 3045 0 1 2604
box 0 0 6 6
use CELL  663
transform -1 0 2996 0 1 2760
box 0 0 6 6
use CELL  664
transform -1 0 2665 0 1 2856
box 0 0 6 6
use CELL  665
transform -1 0 2723 0 1 2604
box 0 0 6 6
use CELL  666
transform -1 0 2616 0 1 2676
box 0 0 6 6
use CELL  667
transform -1 0 2695 0 1 2712
box 0 0 6 6
use CELL  668
transform 1 0 2708 0 1 2664
box 0 0 6 6
use CELL  669
transform 1 0 2638 0 -1 2586
box 0 0 6 6
use CELL  670
transform 1 0 2988 0 1 2796
box 0 0 6 6
use CELL  671
transform 1 0 2662 0 1 2592
box 0 0 6 6
use CELL  672
transform -1 0 2660 0 1 2760
box 0 0 6 6
use CELL  673
transform 1 0 2696 0 1 2844
box 0 0 6 6
use CELL  674
transform -1 0 3079 0 1 2604
box 0 0 6 6
use CELL  675
transform 1 0 2603 0 -1 2670
box 0 0 6 6
use CELL  676
transform -1 0 2703 0 1 2856
box 0 0 6 6
use CELL  677
transform -1 0 2605 0 1 2616
box 0 0 6 6
use CELL  678
transform -1 0 2818 0 1 2844
box 0 0 6 6
use CELL  679
transform -1 0 3062 0 1 2652
box 0 0 6 6
use CELL  680
transform 1 0 2636 0 -1 2562
box 0 0 6 6
use CELL  681
transform -1 0 3153 0 1 2652
box 0 0 6 6
use CELL  682
transform -1 0 2786 0 1 2688
box 0 0 6 6
use CELL  683
transform 1 0 2909 0 1 2808
box 0 0 6 6
use CELL  684
transform 1 0 2932 0 1 2748
box 0 0 6 6
use CELL  685
transform 1 0 2743 0 -1 2634
box 0 0 6 6
use CELL  686
transform -1 0 2648 0 1 2616
box 0 0 6 6
use CELL  687
transform -1 0 2853 0 1 2616
box 0 0 6 6
use CELL  688
transform -1 0 2695 0 1 2556
box 0 0 6 6
use CELL  689
transform -1 0 3019 0 1 2784
box 0 0 6 6
use CELL  690
transform -1 0 2947 0 -1 2610
box 0 0 6 6
use CELL  691
transform 1 0 2665 0 1 2664
box 0 0 6 6
use CELL  692
transform -1 0 3209 0 -1 2694
box 0 0 6 6
use CELL  693
transform 1 0 2917 0 1 2784
box 0 0 6 6
use CELL  694
transform -1 0 2688 0 1 2556
box 0 0 6 6
use CELL  695
transform 1 0 2779 0 1 2772
box 0 0 6 6
use CELL  696
transform 1 0 2882 0 1 2724
box 0 0 6 6
use CELL  697
transform 1 0 2956 0 -1 2766
box 0 0 6 6
use CELL  698
transform -1 0 2620 0 1 2700
box 0 0 6 6
use CELL  699
transform 1 0 2863 0 1 2748
box 0 0 6 6
use CELL  700
transform -1 0 3144 0 1 2700
box 0 0 6 6
use CELL  701
transform -1 0 2780 0 1 2676
box 0 0 6 6
use CELL  702
transform 1 0 2643 0 -1 2598
box 0 0 6 6
use CELL  703
transform 1 0 2592 0 -1 2790
box 0 0 6 6
use CELL  704
transform -1 0 2796 0 1 2700
box 0 0 6 6
use CELL  705
transform -1 0 2807 0 1 2640
box 0 0 6 6
use CELL  706
transform -1 0 2604 0 1 2772
box 0 0 6 6
use CELL  707
transform 1 0 3105 0 1 2676
box 0 0 6 6
use CELL  708
transform -1 0 3042 0 1 2748
box 0 0 6 6
use CELL  709
transform 1 0 3203 0 1 2640
box 0 0 6 6
use CELL  710
transform -1 0 2628 0 -1 2574
box 0 0 6 6
use CELL  711
transform 1 0 2562 0 1 2844
box 0 0 6 6
use CELL  712
transform -1 0 2617 0 1 2544
box 0 0 6 6
use CELL  713
transform -1 0 2709 0 1 2556
box 0 0 6 6
use CELL  714
transform -1 0 3003 0 1 2736
box 0 0 6 6
use CELL  715
transform -1 0 2996 0 1 2748
box 0 0 6 6
use CELL  716
transform -1 0 2788 0 1 2664
box 0 0 6 6
use CELL  717
transform -1 0 2650 0 1 2688
box 0 0 6 6
use CELL  718
transform -1 0 2742 0 -1 2802
box 0 0 6 6
use CELL  719
transform -1 0 2811 0 1 2760
box 0 0 6 6
use CELL  720
transform 1 0 2926 0 1 2580
box 0 0 6 6
use CELL  721
transform -1 0 2733 0 1 2808
box 0 0 6 6
use CELL  722
transform -1 0 3097 0 1 2724
box 0 0 6 6
use CELL  723
transform -1 0 2731 0 1 2580
box 0 0 6 6
use CELL  724
transform 1 0 3064 0 -1 2622
box 0 0 6 6
use CELL  725
transform -1 0 2619 0 1 2784
box 0 0 6 6
use CELL  726
transform -1 0 2838 0 1 2784
box 0 0 6 6
use CELL  727
transform 1 0 2647 0 1 2796
box 0 0 6 6
use CELL  728
transform 1 0 2734 0 1 2568
box 0 0 6 6
use CELL  729
transform -1 0 2836 0 1 2688
box 0 0 6 6
use CELL  730
transform 1 0 2857 0 1 2568
box 0 0 6 6
use CELL  731
transform 1 0 3065 0 -1 2742
box 0 0 6 6
use CELL  732
transform -1 0 2598 0 1 2688
box 0 0 6 6
use CELL  733
transform -1 0 2928 0 1 2832
box 0 0 6 6
use CELL  734
transform -1 0 2944 0 -1 2706
box 0 0 6 6
use CELL  735
transform -1 0 2630 0 1 2580
box 0 0 6 6
use CELL  736
transform 1 0 2606 0 1 2784
box 0 0 6 6
use CELL  737
transform -1 0 2933 0 -1 2814
box 0 0 6 6
use CELL  738
transform -1 0 2639 0 1 2832
box 0 0 6 6
use CELL  739
transform -1 0 2636 0 1 2808
box 0 0 6 6
use CELL  740
transform -1 0 2682 0 1 2676
box 0 0 6 6
use CELL  741
transform -1 0 2785 0 1 2844
box 0 0 6 6
use CELL  742
transform 1 0 2636 0 -1 2778
box 0 0 6 6
use CELL  743
transform 1 0 2962 0 1 2808
box 0 0 6 6
use CELL  744
transform -1 0 3236 0 1 2664
box 0 0 6 6
use CELL  745
transform -1 0 2632 0 1 2760
box 0 0 6 6
use CELL  746
transform -1 0 2662 0 1 2616
box 0 0 6 6
use CELL  747
transform 1 0 2562 0 1 2832
box 0 0 6 6
use CELL  748
transform 1 0 2650 0 1 2556
box 0 0 6 6
use CELL  749
transform -1 0 2813 0 1 2580
box 0 0 6 6
use CELL  750
transform -1 0 2631 0 -1 2550
box 0 0 6 6
use CELL  751
transform -1 0 2599 0 -1 2754
box 0 0 6 6
use CELL  752
transform -1 0 2803 0 1 2856
box 0 0 6 6
use CELL  753
transform 1 0 3087 0 1 2712
box 0 0 6 6
use CELL  754
transform -1 0 2754 0 1 2796
box 0 0 6 6
use CELL  755
transform -1 0 2865 0 1 2592
box 0 0 6 6
use CELL  756
transform 1 0 3052 0 1 2604
box 0 0 6 6
use CELL  757
transform 1 0 3010 0 -1 2598
box 0 0 6 6
use CELL  758
transform -1 0 2717 0 1 2628
box 0 0 6 6
use CELL  759
transform -1 0 2692 0 -1 2586
box 0 0 6 6
use CELL  760
transform -1 0 2802 0 -1 2550
box 0 0 6 6
use CELL  761
transform 1 0 2904 0 -1 2802
box 0 0 6 6
use CELL  762
transform -1 0 2987 0 1 2772
box 0 0 6 6
use CELL  763
transform -1 0 2605 0 1 2784
box 0 0 6 6
use CELL  764
transform 1 0 2889 0 1 2724
box 0 0 6 6
use CELL  765
transform -1 0 2760 0 1 2544
box 0 0 6 6
use CELL  766
transform -1 0 2837 0 1 2568
box 0 0 6 6
use CELL  767
transform -1 0 2679 0 1 2772
box 0 0 6 6
use CELL  768
transform -1 0 2684 0 1 2532
box 0 0 6 6
use CELL  769
transform -1 0 2604 0 1 2820
box 0 0 6 6
use CELL  770
transform 1 0 2618 0 1 2820
box 0 0 6 6
use CELL  771
transform 1 0 2929 0 1 2832
box 0 0 6 6
use CELL  772
transform 1 0 2707 0 -1 2874
box 0 0 6 6
use CELL  773
transform -1 0 2674 0 -1 2610
box 0 0 6 6
use CELL  774
transform -1 0 2532 0 1 2724
box 0 0 6 6
use CELL  775
transform 1 0 2958 0 -1 2802
box 0 0 6 6
use CELL  776
transform -1 0 2766 0 1 2736
box 0 0 6 6
use CELL  777
transform -1 0 2715 0 1 2640
box 0 0 6 6
use CELL  778
transform -1 0 2681 0 1 2544
box 0 0 6 6
use CELL  779
transform 1 0 2664 0 1 2520
box 0 0 6 6
use CELL  780
transform 1 0 2901 0 1 2832
box 0 0 6 6
use CELL  781
transform -1 0 3097 0 1 2736
box 0 0 6 6
use CELL  782
transform 1 0 2738 0 -1 2862
box 0 0 6 6
use CELL  783
transform -1 0 2568 0 1 2808
box 0 0 6 6
use CELL  784
transform 1 0 3019 0 -1 2730
box 0 0 6 6
use CELL  785
transform -1 0 2896 0 1 2820
box 0 0 6 6
use CELL  786
transform 1 0 2661 0 -1 2550
box 0 0 6 6
use CELL  787
transform -1 0 2721 0 1 2652
box 0 0 6 6
use CELL  788
transform -1 0 2724 0 1 2820
box 0 0 6 6
use CELL  789
transform -1 0 2715 0 1 2832
box 0 0 6 6
use CELL  790
transform -1 0 2776 0 1 2712
box 0 0 6 6
use CELL  791
transform -1 0 2714 0 1 2652
box 0 0 6 6
use CELL  792
transform 1 0 2632 0 -1 2694
box 0 0 6 6
use CELL  793
transform 1 0 3174 0 -1 2634
box 0 0 6 6
use CELL  794
transform -1 0 2656 0 1 2844
box 0 0 6 6
use CELL  795
transform 1 0 2951 0 1 2796
box 0 0 6 6
use CELL  796
transform 1 0 2587 0 -1 2766
box 0 0 6 6
use CELL  797
transform -1 0 2617 0 -1 2610
box 0 0 6 6
use CELL  798
transform 1 0 2815 0 1 2832
box 0 0 6 6
use CELL  799
transform -1 0 2996 0 1 2736
box 0 0 6 6
use CELL  800
transform -1 0 2696 0 1 2856
box 0 0 6 6
use CELL  801
transform 1 0 2970 0 1 2784
box 0 0 6 6
use CELL  802
transform 1 0 2748 0 -1 2850
box 0 0 6 6
use CELL  803
transform 1 0 2745 0 -1 2550
box 0 0 6 6
use CELL  804
transform -1 0 2612 0 1 2748
box 0 0 6 6
use CELL  805
transform -1 0 2994 0 1 2772
box 0 0 6 6
use CELL  806
transform 1 0 2648 0 -1 2754
box 0 0 6 6
use CELL  807
transform -1 0 2677 0 1 2532
box 0 0 6 6
use CELL  808
transform 1 0 3161 0 1 2688
box 0 0 6 6
use CELL  809
transform -1 0 3073 0 1 2664
box 0 0 6 6
use CELL  810
transform -1 0 2663 0 1 2568
box 0 0 6 6
use CELL  811
transform -1 0 3135 0 1 2700
box 0 0 6 6
use CELL  812
transform 1 0 2915 0 -1 2838
box 0 0 6 6
use CELL  813
transform -1 0 2637 0 1 2796
box 0 0 6 6
use CELL  814
transform -1 0 2796 0 1 2808
box 0 0 6 6
use CELL  815
transform -1 0 2772 0 1 2820
box 0 0 6 6
use CELL  816
transform -1 0 3083 0 1 2676
box 0 0 6 6
use CELL  817
transform -1 0 2775 0 1 2856
box 0 0 6 6
use CELL  818
transform 1 0 2984 0 1 2784
box 0 0 6 6
use CELL  819
transform -1 0 2635 0 1 2664
box 0 0 6 6
use CELL  820
transform 1 0 2908 0 1 2820
box 0 0 6 6
use CELL  821
transform 1 0 2755 0 1 2676
box 0 0 6 6
use CELL  822
transform -1 0 2612 0 1 2616
box 0 0 6 6
use CELL  823
transform -1 0 3038 0 1 2628
box 0 0 6 6
use CELL  824
transform -1 0 2705 0 1 2628
box 0 0 6 6
use CELL  825
transform 1 0 2883 0 1 2844
box 0 0 6 6
use CELL  826
transform -1 0 3093 0 1 2604
box 0 0 6 6
use CELL  827
transform 1 0 3046 0 1 2700
box 0 0 6 6
use CELL  828
transform -1 0 2654 0 1 2784
box 0 0 6 6
use CELL  829
transform 1 0 2599 0 -1 2694
box 0 0 6 6
use CELL  830
transform 1 0 2871 0 1 2568
box 0 0 6 6
use CELL  831
transform -1 0 3183 0 1 2652
box 0 0 6 6
use CELL  832
transform -1 0 2889 0 1 2784
box 0 0 6 6
use CELL  833
transform -1 0 2616 0 1 2592
box 0 0 6 6
use CELL  834
transform -1 0 2527 0 1 2748
box 0 0 6 6
use CELL  835
transform 1 0 3196 0 1 2688
box 0 0 6 6
use CELL  836
transform -1 0 2625 0 1 2652
box 0 0 6 6
use CELL  837
transform -1 0 2826 0 -1 2802
box 0 0 6 6
use CELL  838
transform 1 0 3155 0 1 2640
box 0 0 6 6
use CELL  839
transform 1 0 2995 0 1 2772
box 0 0 6 6
use CELL  840
transform -1 0 3111 0 1 2736
box 0 0 6 6
use CELL  841
transform -1 0 2588 0 1 2640
box 0 0 6 6
use CELL  842
transform 1 0 2748 0 -1 2538
box 0 0 6 6
use CELL  843
transform -1 0 3015 0 -1 2778
box 0 0 6 6
use CELL  844
transform 1 0 2580 0 -1 2622
box 0 0 6 6
use CELL  845
transform -1 0 3166 0 -1 2634
box 0 0 6 6
use CELL  846
transform -1 0 2942 0 1 2772
box 0 0 6 6
use CELL  847
transform 1 0 2945 0 -1 2586
box 0 0 6 6
use CELL  848
transform -1 0 2599 0 1 2700
box 0 0 6 6
use CELL  849
transform -1 0 2669 0 1 2688
box 0 0 6 6
use CELL  850
transform -1 0 2724 0 1 2796
box 0 0 6 6
use CELL  851
transform -1 0 2602 0 1 2664
box 0 0 6 6
use CELL  852
transform -1 0 3176 0 1 2664
box 0 0 6 6
use CELL  853
transform -1 0 3049 0 1 2748
box 0 0 6 6
use CELL  854
transform -1 0 2654 0 1 2640
box 0 0 6 6
use CELL  855
transform -1 0 2635 0 1 2844
box 0 0 6 6
use CELL  856
transform -1 0 2733 0 1 2724
box 0 0 6 6
use CELL  857
transform 1 0 2694 0 1 2820
box 0 0 6 6
use CELL  858
transform 1 0 2726 0 1 2868
box 0 0 6 6
use CELL  859
transform -1 0 2904 0 1 2580
box 0 0 6 6
use CELL  860
transform -1 0 2630 0 1 2856
box 0 0 6 6
use CELL  861
transform 1 0 2861 0 1 2556
box 0 0 6 6
use CELL  862
transform -1 0 2741 0 1 2604
box 0 0 6 6
use CELL  863
transform -1 0 2715 0 1 2808
box 0 0 6 6
use CELL  864
transform -1 0 2635 0 1 2772
box 0 0 6 6
use CELL  865
transform -1 0 2665 0 1 2556
box 0 0 6 6
use CELL  866
transform -1 0 2727 0 1 2712
box 0 0 6 6
use CELL  867
transform 1 0 3000 0 -1 2790
box 0 0 6 6
use CELL  868
transform 1 0 2942 0 1 2712
box 0 0 6 6
use CELL  869
transform -1 0 2645 0 1 2820
box 0 0 6 6
use CELL  870
transform -1 0 2985 0 1 2616
box 0 0 6 6
use CELL  871
transform 1 0 3050 0 1 2748
box 0 0 6 6
use CELL  872
transform -1 0 3235 0 1 2640
box 0 0 6 6
use CELL  873
transform -1 0 2606 0 1 2760
box 0 0 6 6
use CELL  874
transform -1 0 2708 0 1 2640
box 0 0 6 6
use CELL  875
transform -1 0 2795 0 -1 2550
box 0 0 6 6
use CELL  876
transform -1 0 2653 0 1 2544
box 0 0 6 6
use CELL  877
transform -1 0 2616 0 1 2772
box 0 0 6 6
use CELL  878
transform -1 0 2808 0 1 2808
box 0 0 6 6
use CELL  879
transform -1 0 2617 0 1 2820
box 0 0 6 6
use CELL  880
transform 1 0 2854 0 1 2556
box 0 0 6 6
use CELL  881
transform -1 0 2592 0 1 2748
box 0 0 6 6
use CELL  882
transform -1 0 3096 0 1 2628
box 0 0 6 6
use CELL  883
transform -1 0 2751 0 1 2820
box 0 0 6 6
use CELL  884
transform -1 0 2889 0 1 2808
box 0 0 6 6
use CELL  885
transform 1 0 2711 0 1 2568
box 0 0 6 6
use CELL  886
transform -1 0 2766 0 1 2616
box 0 0 6 6
use CELL  887
transform -1 0 2616 0 -1 2670
box 0 0 6 6
use CELL  888
transform 1 0 2709 0 -1 2778
box 0 0 6 6
use CELL  889
transform 1 0 2666 0 1 2556
box 0 0 6 6
use CELL  890
transform -1 0 2724 0 1 2568
box 0 0 6 6
use CELL  891
transform -1 0 2719 0 1 2868
box 0 0 6 6
use CELL  892
transform 1 0 2890 0 1 2844
box 0 0 6 6
use CELL  893
transform -1 0 2829 0 1 2748
box 0 0 6 6
use CELL  894
transform -1 0 2655 0 1 2604
box 0 0 6 6
use CELL  895
transform 1 0 3093 0 1 2676
box 0 0 6 6
use CELL  896
transform -1 0 2630 0 1 2676
box 0 0 6 6
use CELL  897
transform -1 0 3104 0 1 2724
box 0 0 6 6
use CELL  898
transform 1 0 2963 0 1 2784
box 0 0 6 6
use CELL  899
transform -1 0 2661 0 1 2640
box 0 0 6 6
use CELL  900
transform 1 0 3118 0 1 2736
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 2879 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 2855 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 2633 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 2640 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 2735 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 3059 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 3033 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 2818 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 2757 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 2691 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 2766 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 2708 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 2586 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 2592 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 2595 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 2586 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 2586 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 2815 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 2800 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 2802 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 2838 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 2871 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 2838 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 2921 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 2931 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 2592 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 2569 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 2943 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 2930 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 2868 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 2946 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 2861 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 2839 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 2832 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 2736 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 2740 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 2748 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 2691 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 2703 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 2706 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 2690 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 2694 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 2693 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 2745 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 2673 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 2731 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 2742 0 1 2544
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 2788 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 2797 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 2739 0 1 2544
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 2844 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 2749 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 2718 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 2736 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 2749 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 2876 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 2829 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 2883 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 2817 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 2702 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 2794 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 2785 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 2568 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 2900 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 2914 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 2820 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 2796 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 2790 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 2755 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 2755 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 2872 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 2847 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 2893 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 3122 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 3189 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 3216 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 3197 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 3183 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 3119 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 3186 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 3074 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 3095 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 3155 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 3099 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 3145 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 3171 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 3149 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 2811 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 2742 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 2788 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 2788 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 2803 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 2834 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 2791 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 2759 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 2734 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 2761 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 2801 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 2954 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 2930 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 2775 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 2821 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 2670 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 2676 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 2824 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 2826 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 3137 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 3122 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-109
transform 1 0 3114 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-110
transform 1 0 3047 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-111
transform 1 0 3130 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-112
transform 1 0 3193 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-113
transform 1 0 3144 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-114
transform 1 0 3123 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-115
transform 1 0 3081 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-116
transform 1 0 3088 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-117
transform 1 0 3059 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-118
transform 1 0 2767 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-119
transform 1 0 2773 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-120
transform 1 0 2911 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-121
transform 1 0 2959 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-122
transform 1 0 2968 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-123
transform 1 0 2996 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-124
transform 1 0 3025 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-125
transform 1 0 2953 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-126
transform 1 0 2956 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-127
transform 1 0 2992 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-128
transform 1 0 3055 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-129
transform 1 0 3105 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-130
transform 1 0 2938 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-131
transform 1 0 2851 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-132
transform 1 0 2879 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-133
transform 1 0 2632 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-134
transform 1 0 2706 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-135
transform 1 0 2702 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-136
transform 1 0 2696 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-137
transform 1 0 2711 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-138
transform 1 0 2705 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-139
transform 1 0 2708 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-140
transform 1 0 2693 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-141
transform 1 0 2885 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-142
transform 1 0 2827 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-143
transform 1 0 2705 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-144
transform 1 0 2680 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-145
transform 1 0 2860 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-146
transform 1 0 2835 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-147
transform 1 0 2927 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-148
transform 1 0 2919 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-149
transform 1 0 2938 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-150
transform 1 0 2984 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-151
transform 1 0 2631 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-152
transform 1 0 2789 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-153
transform 1 0 2786 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-154
transform 1 0 3068 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-155
transform 1 0 3018 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-156
transform 1 0 2886 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-157
transform 1 0 2856 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-158
transform 1 0 2822 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-159
transform 1 0 2770 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-160
transform 1 0 3134 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-161
transform 1 0 2653 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-162
transform 1 0 2651 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-163
transform 1 0 2871 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-164
transform 1 0 2923 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-165
transform 1 0 2956 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-166
transform 1 0 3049 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-167
transform 1 0 2875 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-168
transform 1 0 2840 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-169
transform 1 0 2863 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-170
transform 1 0 2913 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-171
transform 1 0 2894 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-172
transform 1 0 2789 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-173
transform 1 0 2813 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-174
transform 1 0 3013 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-175
transform 1 0 2957 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-176
transform 1 0 2956 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-177
transform 1 0 2936 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-178
transform 1 0 2689 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-179
transform 1 0 2724 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-180
transform 1 0 2680 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-181
transform 1 0 2677 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-182
transform 1 0 2676 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-183
transform 1 0 2682 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-184
transform 1 0 2672 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-185
transform 1 0 2668 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-186
transform 1 0 2838 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-187
transform 1 0 2807 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-188
transform 1 0 2908 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-189
transform 1 0 2835 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-190
transform 1 0 2817 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-191
transform 1 0 2764 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-192
transform 1 0 2758 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-193
transform 1 0 2727 0 1 2544
box 0 0 3 6
use FEEDTHRU  F-194
transform 1 0 2761 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-195
transform 1 0 2755 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-196
transform 1 0 2971 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-197
transform 1 0 3025 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-198
transform 1 0 2999 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-199
transform 1 0 3037 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-200
transform 1 0 2960 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-201
transform 1 0 2858 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-202
transform 1 0 2804 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-203
transform 1 0 2835 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-204
transform 1 0 2910 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-205
transform 1 0 2886 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-206
transform 1 0 2974 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-207
transform 1 0 3028 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-208
transform 1 0 3002 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-209
transform 1 0 3040 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-210
transform 1 0 2963 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-211
transform 1 0 2861 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-212
transform 1 0 2807 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-213
transform 1 0 2838 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-214
transform 1 0 2913 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-215
transform 1 0 2889 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-216
transform 1 0 2700 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-217
transform 1 0 2646 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-218
transform 1 0 2804 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-219
transform 1 0 2743 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-220
transform 1 0 2765 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-221
transform 1 0 2650 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-222
transform 1 0 2642 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-223
transform 1 0 2635 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-224
transform 1 0 2849 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-225
transform 1 0 2843 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-226
transform 1 0 2825 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-227
transform 1 0 2832 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-228
transform 1 0 2775 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-229
transform 1 0 2741 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-230
transform 1 0 2644 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-231
transform 1 0 2663 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-232
transform 1 0 2656 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-233
transform 1 0 2727 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-234
transform 1 0 2748 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-235
transform 1 0 2724 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-236
transform 1 0 2722 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-237
transform 1 0 2766 0 1 2856
box 0 0 3 6
use FEEDTHRU  F-238
transform 1 0 2809 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-239
transform 1 0 2752 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-240
transform 1 0 2787 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-241
transform 1 0 2763 0 1 2856
box 0 0 3 6
use FEEDTHRU  F-242
transform 1 0 2980 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-243
transform 1 0 2954 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-244
transform 1 0 3019 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-245
transform 1 0 3052 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-246
transform 1 0 3038 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-247
transform 1 0 3152 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-248
transform 1 0 3174 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-249
transform 1 0 2709 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-250
transform 1 0 2705 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-251
transform 1 0 2877 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-252
transform 1 0 2932 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-253
transform 1 0 2737 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-254
transform 1 0 2700 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-255
transform 1 0 2712 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-256
transform 1 0 2808 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-257
transform 1 0 2644 0 1 2868
box 0 0 3 6
use FEEDTHRU  F-258
transform 1 0 2641 0 1 2868
box 0 0 3 6
use FEEDTHRU  F-259
transform 1 0 2951 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-260
transform 1 0 2977 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-261
transform 1 0 2994 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-262
transform 1 0 3056 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-263
transform 1 0 3098 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-264
transform 1 0 3089 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-265
transform 1 0 3058 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-266
transform 1 0 3044 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-267
transform 1 0 3097 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-268
transform 1 0 3062 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-269
transform 1 0 3029 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-270
transform 1 0 2907 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-271
transform 1 0 2934 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-272
transform 1 0 2963 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-273
transform 1 0 3047 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-274
transform 1 0 3050 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-275
transform 1 0 3055 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-276
transform 1 0 3014 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-277
transform 1 0 3049 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-278
transform 1 0 3010 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-279
transform 1 0 2960 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-280
transform 1 0 2914 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-281
transform 1 0 2908 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-282
transform 1 0 2934 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-283
transform 1 0 2887 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-284
transform 1 0 2890 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-285
transform 1 0 2865 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-286
transform 1 0 2839 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-287
transform 1 0 2799 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-288
transform 1 0 2814 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-289
transform 1 0 2769 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-290
transform 1 0 2751 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-291
transform 1 0 2992 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-292
transform 1 0 2972 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-293
transform 1 0 3016 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-294
transform 1 0 3047 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-295
transform 1 0 2969 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-296
transform 1 0 2974 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-297
transform 1 0 2962 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-298
transform 1 0 2895 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-299
transform 1 0 2866 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-300
transform 1 0 2849 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-301
transform 1 0 2706 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-302
transform 1 0 2715 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-303
transform 1 0 2742 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-304
transform 1 0 2811 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-305
transform 1 0 2856 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-306
transform 1 0 2778 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-307
transform 1 0 2754 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-308
transform 1 0 2685 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-309
transform 1 0 2675 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-310
transform 1 0 2678 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-311
transform 1 0 2687 0 1 2856
box 0 0 3 6
use FEEDTHRU  F-312
transform 1 0 2667 0 1 2868
box 0 0 3 6
use FEEDTHRU  F-313
transform 1 0 2786 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-314
transform 1 0 2815 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-315
transform 1 0 2841 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-316
transform 1 0 2800 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-317
transform 1 0 2786 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-318
transform 1 0 2788 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-319
transform 1 0 2783 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-320
transform 1 0 2762 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-321
transform 1 0 2749 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-322
transform 1 0 2675 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-323
transform 1 0 2684 0 1 2856
box 0 0 3 6
use FEEDTHRU  F-324
transform 1 0 2993 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-325
transform 1 0 2653 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-326
transform 1 0 2715 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-327
transform 1 0 2736 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-328
transform 1 0 2766 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-329
transform 1 0 2654 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-330
transform 1 0 2788 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-331
transform 1 0 2669 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-332
transform 1 0 3025 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-333
transform 1 0 3037 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-334
transform 1 0 3008 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-335
transform 1 0 2677 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-336
transform 1 0 2701 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-337
transform 1 0 2708 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-338
transform 1 0 2689 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-339
transform 1 0 2671 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-340
transform 1 0 2669 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-341
transform 1 0 2675 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-342
transform 1 0 2674 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-343
transform 1 0 2662 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-344
transform 1 0 2683 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-345
transform 1 0 2707 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-346
transform 1 0 2714 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-347
transform 1 0 2695 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-348
transform 1 0 2677 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-349
transform 1 0 2675 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-350
transform 1 0 2681 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-351
transform 1 0 2680 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-352
transform 1 0 2668 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-353
transform 1 0 2643 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-354
transform 1 0 2938 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-355
transform 1 0 2889 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-356
transform 1 0 2865 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-357
transform 1 0 2806 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-358
transform 1 0 2681 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-359
transform 1 0 2683 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-360
transform 1 0 2998 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-361
transform 1 0 2708 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-362
transform 1 0 2988 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-363
transform 1 0 2912 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-364
transform 1 0 2975 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-365
transform 1 0 2724 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-366
transform 1 0 2720 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-367
transform 1 0 2727 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-368
transform 1 0 2730 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-369
transform 1 0 2672 0 1 2856
box 0 0 3 6
use FEEDTHRU  F-370
transform 1 0 3062 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-371
transform 1 0 3062 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-372
transform 1 0 3107 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-373
transform 1 0 3135 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-374
transform 1 0 3167 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-375
transform 1 0 3111 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-376
transform 1 0 3157 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-377
transform 1 0 3168 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-378
transform 1 0 3200 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-379
transform 1 0 3157 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-380
transform 1 0 3097 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-381
transform 1 0 3019 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-382
transform 1 0 2981 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-383
transform 1 0 2932 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-384
transform 1 0 2884 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-385
transform 1 0 2787 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-386
transform 1 0 2749 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-387
transform 1 0 2793 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-388
transform 1 0 2760 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-389
transform 1 0 2767 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-390
transform 1 0 2760 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-391
transform 1 0 2811 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-392
transform 1 0 2778 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-393
transform 1 0 2702 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-394
transform 1 0 2711 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-395
transform 1 0 2679 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-396
transform 1 0 2681 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-397
transform 1 0 2697 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-398
transform 1 0 2667 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-399
transform 1 0 2699 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-400
transform 1 0 2684 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-401
transform 1 0 2693 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-402
transform 1 0 2696 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-403
transform 1 0 2854 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-404
transform 1 0 2883 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-405
transform 1 0 2968 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-406
transform 1 0 2930 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-407
transform 1 0 2734 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-408
transform 1 0 2734 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-409
transform 1 0 2990 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-410
transform 1 0 2752 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-411
transform 1 0 2777 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-412
transform 1 0 2774 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-413
transform 1 0 2749 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-414
transform 1 0 2740 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-415
transform 1 0 2740 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-416
transform 1 0 2743 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-417
transform 1 0 2731 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-418
transform 1 0 2721 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-419
transform 1 0 2702 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-420
transform 1 0 2739 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-421
transform 1 0 2769 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-422
transform 1 0 2751 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-423
transform 1 0 2761 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-424
transform 1 0 2663 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-425
transform 1 0 2681 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-426
transform 1 0 2643 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-427
transform 1 0 2652 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-428
transform 1 0 2630 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-429
transform 1 0 2803 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-430
transform 1 0 2840 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-431
transform 1 0 2681 0 1 2856
box 0 0 3 6
use FEEDTHRU  F-432
transform 1 0 2743 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-433
transform 1 0 2798 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-434
transform 1 0 2792 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-435
transform 1 0 2774 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-436
transform 1 0 2871 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-437
transform 1 0 2892 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-438
transform 1 0 2781 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-439
transform 1 0 2831 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-440
transform 1 0 2882 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-441
transform 1 0 2896 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-442
transform 1 0 2915 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-443
transform 1 0 2999 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-444
transform 1 0 3022 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-445
transform 1 0 3010 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-446
transform 1 0 3077 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-447
transform 1 0 2760 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-448
transform 1 0 2781 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-449
transform 1 0 3071 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-450
transform 1 0 3002 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-451
transform 1 0 2991 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-452
transform 1 0 2947 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-453
transform 1 0 2911 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-454
transform 1 0 2862 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-455
transform 1 0 2819 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-456
transform 1 0 2807 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-457
transform 1 0 2774 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-458
transform 1 0 2758 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-459
transform 1 0 2731 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-460
transform 1 0 2702 0 1 2544
box 0 0 3 6
use FEEDTHRU  F-461
transform 1 0 3027 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-462
transform 1 0 2670 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-463
transform 1 0 2667 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-464
transform 1 0 2690 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-465
transform 1 0 2672 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-466
transform 1 0 2667 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-467
transform 1 0 2672 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-468
transform 1 0 2694 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-469
transform 1 0 2751 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-470
transform 1 0 2798 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-471
transform 1 0 2812 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-472
transform 1 0 2835 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-473
transform 1 0 2863 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-474
transform 1 0 2825 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-475
transform 1 0 2815 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-476
transform 1 0 2705 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-477
transform 1 0 2715 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-478
transform 1 0 2705 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-479
transform 1 0 2790 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-480
transform 1 0 2674 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-481
transform 1 0 2674 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-482
transform 1 0 2660 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-483
transform 1 0 2679 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-484
transform 1 0 2727 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-485
transform 1 0 2731 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-486
transform 1 0 2739 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-487
transform 1 0 2742 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-488
transform 1 0 2760 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-489
transform 1 0 2724 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-490
transform 1 0 2700 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-491
transform 1 0 2687 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-492
transform 1 0 2733 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-493
transform 1 0 2737 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-494
transform 1 0 2745 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-495
transform 1 0 2702 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-496
transform 1 0 2697 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-497
transform 1 0 2708 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-498
transform 1 0 2703 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-499
transform 1 0 2699 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-500
transform 1 0 3092 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-501
transform 1 0 3050 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-502
transform 1 0 2931 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-503
transform 1 0 2923 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-504
transform 1 0 2876 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-505
transform 1 0 2914 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-506
transform 1 0 2777 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-507
transform 1 0 3092 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-508
transform 1 0 3130 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-509
transform 1 0 3071 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-510
transform 1 0 3111 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-511
transform 1 0 3092 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-512
transform 1 0 3107 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-513
transform 1 0 3044 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-514
transform 1 0 3041 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-515
transform 1 0 3094 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-516
transform 1 0 3059 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-517
transform 1 0 3026 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-518
transform 1 0 3074 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-519
transform 1 0 3095 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-520
transform 1 0 2820 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-521
transform 1 0 2865 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-522
transform 1 0 2984 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-523
transform 1 0 2853 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-524
transform 1 0 2709 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-525
transform 1 0 2746 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-526
transform 1 0 2715 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-527
transform 1 0 2809 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-528
transform 1 0 2796 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-529
transform 1 0 3046 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-530
transform 1 0 2684 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-531
transform 1 0 2644 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-532
transform 1 0 3002 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-533
transform 1 0 2962 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-534
transform 1 0 2956 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-535
transform 1 0 2930 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-536
transform 1 0 2971 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-537
transform 1 0 2924 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-538
transform 1 0 2905 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-539
transform 1 0 2891 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-540
transform 1 0 2873 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-541
transform 1 0 2824 0 1 2856
box 0 0 3 6
use FEEDTHRU  F-542
transform 1 0 3023 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-543
transform 1 0 2979 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-544
transform 1 0 2646 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-545
transform 1 0 2672 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-546
transform 1 0 2675 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-547
transform 1 0 2670 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-548
transform 1 0 2666 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-549
transform 1 0 2667 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-550
transform 1 0 2655 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-551
transform 1 0 2667 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-552
transform 1 0 2877 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-553
transform 1 0 2863 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-554
transform 1 0 2848 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-555
transform 1 0 2883 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-556
transform 1 0 2875 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-557
transform 1 0 2855 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-558
transform 1 0 2873 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-559
transform 1 0 2849 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-560
transform 1 0 2736 0 1 2544
box 0 0 3 6
use FEEDTHRU  F-561
transform 1 0 2774 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-562
transform 1 0 2733 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-563
transform 1 0 2715 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-564
transform 1 0 2727 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-565
transform 1 0 3146 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-566
transform 1 0 3090 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-567
transform 1 0 3126 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-568
transform 1 0 3137 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-569
transform 1 0 2758 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-570
transform 1 0 2768 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-571
transform 1 0 2765 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-572
transform 1 0 2752 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-573
transform 1 0 2852 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-574
transform 1 0 2725 0 1 2856
box 0 0 3 6
use FEEDTHRU  F-575
transform 1 0 2705 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-576
transform 1 0 2728 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-577
transform 1 0 2754 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-578
transform 1 0 2763 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-579
transform 1 0 2793 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-580
transform 1 0 2778 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-581
transform 1 0 2752 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-582
transform 1 0 2754 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-583
transform 1 0 2742 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-584
transform 1 0 2721 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-585
transform 1 0 2740 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-586
transform 1 0 2762 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-587
transform 1 0 2768 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-588
transform 1 0 3173 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-589
transform 1 0 3136 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-590
transform 1 0 3179 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-591
transform 1 0 3142 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-592
transform 1 0 3088 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-593
transform 1 0 3016 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-594
transform 1 0 2978 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-595
transform 1 0 2857 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-596
transform 1 0 2752 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-597
transform 1 0 2752 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-598
transform 1 0 2787 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-599
transform 1 0 2793 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-600
transform 1 0 2889 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-601
transform 1 0 2924 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-602
transform 1 0 2966 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-603
transform 1 0 2942 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-604
transform 1 0 2926 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-605
transform 1 0 2891 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-606
transform 1 0 2911 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-607
transform 1 0 2898 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-608
transform 1 0 2902 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-609
transform 1 0 2825 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-610
transform 1 0 2875 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-611
transform 1 0 2802 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-612
transform 1 0 2784 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-613
transform 1 0 2803 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-614
transform 1 0 2790 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-615
transform 1 0 2808 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-616
transform 1 0 2775 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-617
transform 1 0 2763 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-618
transform 1 0 2740 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-619
transform 1 0 2724 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-620
transform 1 0 2728 0 1 2856
box 0 0 3 6
use FEEDTHRU  F-621
transform 1 0 2683 0 1 2868
box 0 0 3 6
use FEEDTHRU  F-622
transform 1 0 2722 0 1 2856
box 0 0 3 6
use FEEDTHRU  F-623
transform 1 0 3086 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-624
transform 1 0 3053 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-625
transform 1 0 2768 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-626
transform 1 0 2775 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-627
transform 1 0 2772 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-628
transform 1 0 2739 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-629
transform 1 0 2764 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-630
transform 1 0 2766 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-631
transform 1 0 2754 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-632
transform 1 0 2739 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-633
transform 1 0 2811 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-634
transform 1 0 2806 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-635
transform 1 0 2918 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-636
transform 1 0 2932 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-637
transform 1 0 2912 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-638
transform 1 0 2927 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-639
transform 1 0 2802 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-640
transform 1 0 2840 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-641
transform 1 0 2830 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-642
transform 1 0 2864 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-643
transform 1 0 2866 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-644
transform 1 0 2873 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-645
transform 1 0 2905 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-646
transform 1 0 2874 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-647
transform 1 0 2848 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-648
transform 1 0 2804 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-649
transform 1 0 2810 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-650
transform 1 0 2789 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-651
transform 1 0 2820 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-652
transform 1 0 2928 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-653
transform 1 0 2751 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-654
transform 1 0 2775 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-655
transform 1 0 2775 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-656
transform 1 0 2815 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-657
transform 1 0 2781 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-658
transform 1 0 2813 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-659
transform 1 0 2791 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-660
transform 1 0 2817 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-661
transform 1 0 2818 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-662
transform 1 0 3065 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-663
transform 1 0 2704 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-664
transform 1 0 2744 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-665
transform 1 0 2769 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-666
transform 1 0 2775 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-667
transform 1 0 2758 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-668
transform 1 0 2838 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-669
transform 1 0 2920 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-670
transform 1 0 3007 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-671
transform 1 0 3062 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-672
transform 1 0 3089 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-673
transform 1 0 3127 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-674
transform 1 0 3068 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-675
transform 1 0 3108 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-676
transform 1 0 2911 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-677
transform 1 0 2845 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-678
transform 1 0 2928 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-679
transform 1 0 2973 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-680
transform 1 0 3014 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-681
transform 1 0 3077 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-682
transform 1 0 3062 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-683
transform 1 0 3061 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-684
transform 1 0 3032 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-685
transform 1 0 3085 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-686
transform 1 0 3037 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-687
transform 1 0 3017 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-688
transform 1 0 2976 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-689
transform 1 0 2954 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-690
transform 1 0 2917 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-691
transform 1 0 2934 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-692
transform 1 0 2924 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-693
transform 1 0 3219 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-694
transform 1 0 3124 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-695
transform 1 0 3070 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-696
transform 1 0 2842 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-697
transform 1 0 2830 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-698
transform 1 0 2874 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-699
transform 1 0 2916 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-700
transform 1 0 2871 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-701
transform 1 0 2933 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-702
transform 1 0 2895 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-703
transform 1 0 2766 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-704
transform 1 0 2778 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-705
transform 1 0 2790 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-706
transform 1 0 2810 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-707
transform 1 0 2836 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-708
transform 1 0 2844 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-709
transform 1 0 2993 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-710
transform 1 0 2699 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-711
transform 1 0 2714 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-712
transform 1 0 2766 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-713
transform 1 0 2780 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-714
transform 1 0 2798 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-715
transform 1 0 2818 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-716
transform 1 0 2799 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-717
transform 1 0 2805 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-718
transform 1 0 2945 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-719
transform 1 0 3023 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-720
transform 1 0 2990 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-721
transform 1 0 3025 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-722
transform 1 0 2981 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-723
transform 1 0 3013 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-724
transform 1 0 2950 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-725
transform 1 0 2948 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-726
transform 1 0 2838 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-727
transform 1 0 2811 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-728
transform 1 0 2771 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-729
transform 1 0 2808 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-730
transform 1 0 2835 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-731
transform 1 0 2898 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-732
transform 1 0 2943 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-733
transform 1 0 2960 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-734
transform 1 0 2908 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-735
transform 1 0 3094 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-736
transform 1 0 3148 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-737
transform 1 0 3185 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-738
transform 1 0 3028 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-739
transform 1 0 2990 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-740
transform 1 0 2922 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-741
transform 1 0 2903 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-742
transform 1 0 2719 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-743
transform 1 0 2743 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-744
transform 1 0 2751 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-745
transform 1 0 2755 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-746
transform 1 0 2745 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-747
transform 1 0 2763 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-748
transform 1 0 2772 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-749
transform 1 0 3165 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-750
transform 1 0 3197 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-751
transform 1 0 3154 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-752
transform 1 0 2890 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-753
transform 1 0 2867 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-754
transform 1 0 2872 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-755
transform 1 0 2869 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-756
transform 1 0 2751 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-757
transform 1 0 2736 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-758
transform 1 0 2777 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-759
transform 1 0 2797 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-760
transform 1 0 2808 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-761
transform 1 0 2743 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-762
transform 1 0 2746 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-763
transform 1 0 2921 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-764
transform 1 0 2935 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-765
transform 1 0 2945 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-766
transform 1 0 2987 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-767
transform 1 0 2933 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-768
transform 1 0 2965 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-769
transform 1 0 2927 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-770
transform 1 0 2953 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-771
transform 1 0 2954 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-772
transform 1 0 2857 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-773
transform 1 0 3003 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-774
transform 1 0 3009 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-775
transform 1 0 3059 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-776
transform 1 0 3015 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-777
transform 1 0 3065 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-778
transform 1 0 2931 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-779
transform 1 0 2881 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-780
transform 1 0 2856 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-781
transform 1 0 2861 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-782
transform 1 0 2820 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-783
transform 1 0 2880 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-784
transform 1 0 2814 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-785
transform 1 0 2887 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-786
transform 1 0 2862 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-787
transform 1 0 2873 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-788
transform 1 0 2826 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-789
transform 1 0 2796 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-790
transform 1 0 2977 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-791
transform 1 0 3043 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-792
transform 1 0 3011 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-793
transform 1 0 3043 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-794
transform 1 0 3082 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-795
transform 1 0 3034 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-796
transform 1 0 3053 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-797
transform 1 0 3050 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-798
transform 1 0 3056 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-799
transform 1 0 3017 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-800
transform 1 0 2980 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-801
transform 1 0 2971 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-802
transform 1 0 2946 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-803
transform 1 0 2823 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-804
transform 1 0 2828 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-805
transform 1 0 2914 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-806
transform 1 0 2966 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-807
transform 1 0 2973 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-808
transform 1 0 3020 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-809
transform 1 0 3028 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-810
transform 1 0 2841 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-811
transform 1 0 2889 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-812
transform 1 0 2781 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-813
transform 1 0 2797 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-814
transform 1 0 2781 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-815
transform 1 0 3160 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-816
transform 1 0 3159 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-817
transform 1 0 3191 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-818
transform 1 0 3108 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-819
transform 1 0 3134 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-820
transform 1 0 3125 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-821
transform 1 0 2736 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-822
transform 1 0 3047 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-823
transform 1 0 3089 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-824
transform 1 0 2822 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-825
transform 1 0 2833 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-826
transform 1 0 2850 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-827
transform 1 0 2902 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-828
transform 1 0 2870 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-829
transform 1 0 2878 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-830
transform 1 0 2888 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-831
transform 1 0 2882 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-832
transform 1 0 2858 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-833
transform 1 0 3044 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-834
transform 1 0 2969 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-835
transform 1 0 2716 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-836
transform 1 0 2724 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-837
transform 1 0 2722 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-838
transform 1 0 2772 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-839
transform 1 0 2799 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-840
transform 1 0 2880 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-841
transform 1 0 2882 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-842
transform 1 0 2924 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-843
transform 1 0 2909 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-844
transform 1 0 2929 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-845
transform 1 0 2915 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-846
transform 1 0 2959 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-847
transform 1 0 2892 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-848
transform 1 0 2863 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-849
transform 1 0 2846 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-850
transform 1 0 2818 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-851
transform 1 0 2829 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-852
transform 1 0 2836 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-853
transform 1 0 2858 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-854
transform 1 0 2896 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-855
transform 1 0 2901 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-856
transform 1 0 2971 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-857
transform 1 0 2806 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-858
transform 1 0 2797 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-859
transform 1 0 2799 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-860
transform 1 0 2835 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-861
transform 1 0 2812 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-862
transform 1 0 2822 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-863
transform 1 0 2860 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-864
transform 1 0 2832 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-865
transform 1 0 2809 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-866
transform 1 0 2795 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-867
transform 1 0 2748 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-868
transform 1 0 2877 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-869
transform 1 0 2910 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-870
transform 1 0 2868 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-871
transform 1 0 2823 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-872
transform 1 0 2821 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-873
transform 1 0 2818 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-874
transform 1 0 3015 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-875
transform 1 0 2990 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-876
transform 1 0 3029 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-877
transform 1 0 3038 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-878
transform 1 0 3056 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-879
transform 1 0 3085 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-880
transform 1 0 3078 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-881
transform 1 0 2947 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-882
transform 1 0 2880 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-883
transform 1 0 2851 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-884
transform 1 0 2840 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-885
transform 1 0 2812 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-886
transform 1 0 2817 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-887
transform 1 0 2796 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-888
transform 1 0 2812 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-889
transform 1 0 2738 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-890
transform 1 0 2760 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-891
transform 1 0 2829 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-892
transform 1 0 2822 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-893
transform 1 0 2840 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-894
transform 1 0 2846 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-895
transform 1 0 2860 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-896
transform 1 0 2837 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-897
transform 1 0 2872 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-898
transform 1 0 2726 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-899
transform 1 0 2754 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-900
transform 1 0 2811 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-901
transform 1 0 2720 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-902
transform 1 0 2748 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-903
transform 1 0 2800 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-904
transform 1 0 2781 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-905
transform 1 0 2799 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-906
transform 1 0 2748 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-907
transform 1 0 2739 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-908
transform 1 0 3046 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-909
transform 1 0 3029 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-910
transform 1 0 2981 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-911
transform 1 0 2969 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-912
transform 1 0 3013 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-913
transform 1 0 3008 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-914
transform 1 0 3041 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-915
transform 1 0 2993 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-916
transform 1 0 2946 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-917
transform 1 0 2917 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-918
transform 1 0 2944 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-919
transform 1 0 3001 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-920
transform 1 0 3061 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-921
transform 1 0 3102 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-922
transform 1 0 3140 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-923
transform 1 0 3113 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-924
transform 1 0 3105 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-925
transform 1 0 3074 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-926
transform 1 0 3121 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-927
transform 1 0 3083 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-928
transform 1 0 3056 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-929
transform 1 0 3016 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-930
transform 1 0 3028 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-931
transform 1 0 2929 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-932
transform 1 0 2977 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-933
transform 1 0 3043 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-934
transform 1 0 3084 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-935
transform 1 0 3122 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-936
transform 1 0 3200 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-937
transform 1 0 3186 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-938
transform 1 0 3059 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-939
transform 1 0 3106 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-940
transform 1 0 3065 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-941
transform 1 0 3038 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-942
transform 1 0 3028 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-943
transform 1 0 3040 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-944
transform 1 0 2743 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-945
transform 1 0 2740 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-946
transform 1 0 2728 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-947
transform 1 0 2790 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-948
transform 1 0 2859 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-949
transform 1 0 2894 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-950
transform 1 0 2930 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-951
transform 1 0 2915 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-952
transform 1 0 2920 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-953
transform 1 0 2909 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-954
transform 1 0 2974 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-955
transform 1 0 2904 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-956
transform 1 0 2899 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-957
transform 1 0 2918 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-958
transform 1 0 2895 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-959
transform 1 0 2941 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-960
transform 1 0 2892 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-961
transform 1 0 2868 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-962
transform 1 0 2851 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-963
transform 1 0 2972 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-964
transform 1 0 2972 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-965
transform 1 0 2967 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-966
transform 1 0 2993 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-967
transform 1 0 3016 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-968
transform 1 0 3058 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-969
transform 1 0 3050 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-970
transform 1 0 2893 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-971
transform 1 0 2879 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-972
transform 1 0 2985 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-973
transform 1 0 2901 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-974
transform 1 0 2877 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-975
transform 1 0 2837 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-976
transform 1 0 2866 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-977
transform 1 0 2864 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-978
transform 1 0 2951 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-979
transform 1 0 2869 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-980
transform 1 0 2900 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-981
transform 1 0 2885 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-982
transform 1 0 3044 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-983
transform 1 0 2978 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-984
transform 1 0 2977 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-985
transform 1 0 2939 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-986
transform 1 0 2989 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-987
transform 1 0 2935 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-988
transform 1 0 2905 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-989
transform 1 0 2895 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-990
transform 1 0 2884 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-991
transform 1 0 2869 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-992
transform 1 0 2844 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-993
transform 1 0 2871 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-994
transform 1 0 2892 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-995
transform 1 0 2880 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-996
transform 1 0 2897 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-997
transform 1 0 3068 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-998
transform 1 0 3041 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-999
transform 1 0 2923 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1000
transform 1 0 2939 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1001
transform 1 0 2963 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1002
transform 1 0 2921 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1003
transform 1 0 2886 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1004
transform 1 0 2751 0 1 2544
box 0 0 3 6
use FEEDTHRU  F-1005
transform 1 0 2791 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-1006
transform 1 0 2800 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-1007
transform 1 0 2787 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1008
transform 1 0 2789 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-1009
transform 1 0 2803 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-1010
transform 1 0 2823 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1011
transform 1 0 2848 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1012
transform 1 0 2785 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-1013
transform 1 0 2785 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-1014
transform 1 0 2760 0 1 2856
box 0 0 3 6
use FEEDTHRU  F-1015
transform 1 0 2808 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-1016
transform 1 0 2853 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-1017
transform 1 0 2749 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-1018
transform 1 0 2987 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1019
transform 1 0 2941 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-1020
transform 1 0 2922 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-1021
transform 1 0 2981 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-1022
transform 1 0 2929 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1023
transform 1 0 2980 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1024
transform 1 0 2887 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-1025
transform 1 0 2876 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-1026
transform 1 0 2860 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1027
transform 1 0 2910 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1028
transform 1 0 2890 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-1029
transform 1 0 2879 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-1030
transform 1 0 2863 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1031
transform 1 0 2857 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-1032
transform 1 0 2832 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-1033
transform 1 0 2987 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1034
transform 1 0 2961 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1035
transform 1 0 2883 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-1036
transform 1 0 2853 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-1037
transform 1 0 2819 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-1038
transform 1 0 2782 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-1039
transform 1 0 2767 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-1040
transform 1 0 2766 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1041
transform 1 0 2866 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-1042
transform 1 0 2824 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1043
transform 1 0 2829 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1044
transform 1 0 2854 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1045
transform 1 0 2828 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1046
transform 1 0 2827 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1047
transform 1 0 2897 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1048
transform 1 0 2899 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1049
transform 1 0 2933 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1050
transform 1 0 2949 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1051
transform 1 0 2877 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-1052
transform 1 0 2847 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-1053
transform 1 0 2813 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-1054
transform 1 0 2776 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-1055
transform 1 0 2761 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-1056
transform 1 0 2804 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-1057
transform 1 0 2838 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-1058
transform 1 0 2931 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-1059
transform 1 0 2976 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1060
transform 1 0 3017 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1061
transform 1 0 3080 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1062
transform 1 0 3065 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1063
transform 1 0 3064 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1064
transform 1 0 2878 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1065
transform 1 0 2896 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-1066
transform 1 0 2877 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-1067
transform 1 0 2998 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1068
transform 1 0 2975 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-1069
transform 1 0 2955 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-1070
transform 1 0 3001 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1071
transform 1 0 2978 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-1072
transform 1 0 2958 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-1073
transform 1 0 2935 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1074
transform 1 0 3005 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-1075
transform 1 0 2965 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-1076
transform 1 0 2999 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1077
transform 1 0 2928 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1078
transform 1 0 2847 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-1079
transform 1 0 2820 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-1080
transform 1 0 2789 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-1081
transform 1 0 2916 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1082
transform 1 0 2850 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-1083
transform 1 0 2823 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-1084
transform 1 0 2792 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-1085
transform 1 0 2815 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1086
transform 1 0 2843 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-1087
transform 1 0 2842 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-1088
transform 1 0 2862 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1089
transform 1 0 2896 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1090
transform 1 0 2874 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-1091
transform 1 0 2898 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-1092
transform 1 0 2853 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-1093
transform 1 0 2880 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-1094
transform 1 0 2827 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-1095
transform 1 0 2821 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-1096
transform 1 0 2823 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1097
transform 1 0 2849 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1098
transform 1 0 2848 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1099
transform 1 0 2876 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1100
transform 1 0 2876 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1101
transform 1 0 2852 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1102
transform 1 0 2843 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1103
transform 1 0 2842 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1104
transform 1 0 3124 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1105
transform 1 0 3086 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1106
transform 1 0 3059 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-1107
transform 1 0 3041 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1108
transform 1 0 3059 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1109
transform 1 0 3038 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1110
transform 1 0 3148 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1111
transform 1 0 3102 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1112
transform 1 0 3020 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1113
transform 1 0 3053 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1114
transform 1 0 3032 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1115
transform 1 0 2995 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1116
transform 1 0 2987 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1117
transform 1 0 3158 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1118
transform 1 0 3098 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1119
transform 1 0 2975 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1120
transform 1 0 2970 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-1121
transform 1 0 2996 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-1122
transform 1 0 2938 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1123
transform 1 0 3055 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1124
transform 1 0 2989 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1125
transform 1 0 2966 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-1126
transform 1 0 3016 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1127
transform 1 0 2984 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1128
transform 1 0 3028 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1129
transform 1 0 2927 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1130
transform 1 0 3026 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1131
transform 1 0 2763 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-1132
transform 1 0 2733 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-1133
transform 1 0 2712 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-1134
transform 1 0 2785 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-1135
transform 1 0 2801 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-1136
transform 1 0 2832 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-1137
transform 1 0 2787 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1138
transform 1 0 2953 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1139
transform 1 0 2912 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1140
transform 1 0 2917 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1141
transform 1 0 2951 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1142
transform 1 0 2981 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1143
transform 1 0 2957 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1144
transform 1 0 2812 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1145
transform 1 0 2773 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-1146
transform 1 0 2767 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-1147
transform 1 0 2776 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-1148
transform 1 0 2770 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-1149
transform 1 0 2751 0 1 2856
box 0 0 3 6
use FEEDTHRU  F-1150
transform 1 0 3019 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1151
transform 1 0 3061 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1152
transform 1 0 2945 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1153
transform 1 0 3117 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1154
transform 1 0 2984 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1155
transform 1 0 2827 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-1156
transform 1 0 2833 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-1157
transform 1 0 2847 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-1158
transform 1 0 2865 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-1159
transform 1 0 2901 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-1160
transform 1 0 2914 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-1161
transform 1 0 2962 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-1162
transform 1 0 2971 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-1163
transform 1 0 2926 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-1164
transform 1 0 2902 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1165
transform 1 0 2916 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-1166
transform 1 0 2936 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-1167
transform 1 0 2953 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1168
transform 1 0 2995 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1169
transform 1 0 2957 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1170
transform 1 0 2959 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1171
transform 1 0 2996 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1172
transform 1 0 3035 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1173
transform 1 0 3008 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1174
transform 1 0 2955 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1175
transform 1 0 2959 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-1176
transform 1 0 2926 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-1177
transform 1 0 2874 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-1178
transform 1 0 2927 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1179
transform 1 0 2951 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1180
transform 1 0 2814 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-1181
transform 1 0 2830 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1182
transform 1 0 2851 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-1183
transform 1 0 2826 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-1184
transform 1 0 2833 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-1185
transform 1 0 2850 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-1186
transform 1 0 2778 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-1187
transform 1 0 2773 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-1188
transform 1 0 3129 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1189
transform 1 0 3014 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1190
transform 1 0 2939 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1191
transform 1 0 2948 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1192
transform 1 0 2933 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1193
transform 1 0 2903 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1194
transform 1 0 2901 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1195
transform 1 0 2707 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-1196
transform 1 0 2732 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-1197
transform 1 0 2874 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-1198
transform 1 0 2865 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-1199
transform 1 0 2879 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-1200
transform 1 0 2868 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-1201
transform 1 0 2893 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-1202
transform 1 0 2872 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1203
transform 1 0 2826 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1204
transform 1 0 2861 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1205
transform 1 0 2885 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1206
transform 1 0 2891 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1207
transform 1 0 2797 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-1208
transform 1 0 2803 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-1209
transform 1 0 2811 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-1210
transform 1 0 2856 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-1211
transform 1 0 2912 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1212
transform 1 0 2867 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-1213
transform 1 0 2853 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-1214
transform 1 0 2859 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-1215
transform 1 0 2823 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-1216
transform 1 0 2757 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-1217
transform 1 0 2737 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-1218
transform 1 0 2766 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-1219
transform 1 0 2925 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-1220
transform 1 0 2793 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-1221
transform 1 0 2816 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1222
transform 1 0 2800 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1223
transform 1 0 2804 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1224
transform 1 0 2796 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-1225
transform 1 0 2820 0 1 2808
box 0 0 3 6
use FEEDTHRU  F-1226
transform 1 0 2877 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-1227
transform 1 0 2746 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-1228
transform 1 0 2775 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-1229
transform 1 0 2808 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-1230
transform 1 0 2868 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1231
transform 1 0 2897 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1232
transform 1 0 2640 0 1 2532
box 0 0 3 6
use FEEDTHRU  F-1233
transform 1 0 2870 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1234
transform 1 0 2846 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1235
transform 1 0 2782 0 1 2556
box 0 0 3 6
use FEEDTHRU  F-1236
transform 1 0 2834 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1237
transform 1 0 2834 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1238
transform 1 0 2828 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1239
transform 1 0 2836 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1240
transform 1 0 2856 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1241
transform 1 0 2878 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1242
transform 1 0 2855 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1243
transform 1 0 2854 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1244
transform 1 0 2870 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1245
transform 1 0 2864 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1246
transform 1 0 2882 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1247
transform 1 0 2810 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1248
transform 1 0 2957 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1249
transform 1 0 2951 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1250
transform 1 0 3058 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1251
transform 1 0 2995 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-1252
transform 1 0 2826 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-1253
transform 1 0 2801 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-1254
transform 1 0 2711 0 1 2544
box 0 0 3 6
use FEEDTHRU  F-1255
transform 1 0 3170 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1256
transform 1 0 3114 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1257
transform 1 0 2983 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1258
transform 1 0 3002 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1259
transform 1 0 3005 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1260
transform 1 0 2996 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1261
transform 1 0 2967 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1262
transform 1 0 2904 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-1263
transform 1 0 2871 0 1 2592
box 0 0 3 6
use FEEDTHRU  F-1264
transform 1 0 2935 0 1 2580
box 0 0 3 6
use FEEDTHRU  F-1265
transform 1 0 2887 0 1 2568
box 0 0 3 6
use FEEDTHRU  F-1266
transform 1 0 2956 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1267
transform 1 0 2766 0 1 2604
box 0 0 3 6
use FEEDTHRU  F-1268
transform 1 0 2817 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1269
transform 1 0 2840 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1270
transform 1 0 2846 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1271
transform 1 0 2852 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1272
transform 1 0 2836 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1273
transform 1 0 2871 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-1274
transform 1 0 2900 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1275
transform 1 0 3032 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1276
transform 1 0 2888 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1277
transform 1 0 2862 0 1 2616
box 0 0 3 6
use FEEDTHRU  F-1278
transform 1 0 2796 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1279
transform 1 0 2776 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-1280
transform 1 0 2765 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-1281
transform 1 0 2721 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1282
transform 1 0 2784 0 1 2796
box 0 0 3 6
use FEEDTHRU  F-1283
transform 1 0 2803 0 1 2844
box 0 0 3 6
use FEEDTHRU  F-1284
transform 1 0 2854 0 1 2832
box 0 0 3 6
use FEEDTHRU  F-1285
transform 1 0 2805 0 1 2820
box 0 0 3 6
use FEEDTHRU  F-1286
transform 1 0 2758 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-1287
transform 1 0 2748 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-1288
transform 1 0 2766 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-1289
transform 1 0 2730 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1290
transform 1 0 2774 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-1291
transform 1 0 2800 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-1292
transform 1 0 2805 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1293
transform 1 0 2824 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1294
transform 1 0 2807 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1295
transform 1 0 2803 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1296
transform 1 0 2819 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1297
transform 1 0 2807 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1298
transform 1 0 2801 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1299
transform 1 0 2769 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1300
transform 1 0 2909 0 1 2628
box 0 0 3 6
use FEEDTHRU  F-1301
transform 1 0 2978 0 1 2640
box 0 0 3 6
use FEEDTHRU  F-1302
transform 1 0 2918 0 1 2652
box 0 0 3 6
use FEEDTHRU  F-1303
transform 1 0 3022 0 1 2664
box 0 0 3 6
use FEEDTHRU  F-1304
transform 1 0 2903 0 1 2676
box 0 0 3 6
use FEEDTHRU  F-1305
transform 1 0 2935 0 1 2688
box 0 0 3 6
use FEEDTHRU  F-1306
transform 1 0 2907 0 1 2700
box 0 0 3 6
use FEEDTHRU  F-1307
transform 1 0 2893 0 1 2712
box 0 0 3 6
use FEEDTHRU  F-1308
transform 1 0 2873 0 1 2724
box 0 0 3 6
use FEEDTHRU  F-1309
transform 1 0 2881 0 1 2736
box 0 0 3 6
use FEEDTHRU  F-1310
transform 1 0 2899 0 1 2748
box 0 0 3 6
use FEEDTHRU  F-1311
transform 1 0 2880 0 1 2760
box 0 0 3 6
use FEEDTHRU  F-1312
transform 1 0 2855 0 1 2772
box 0 0 3 6
use FEEDTHRU  F-1313
transform 1 0 2847 0 1 2784
box 0 0 3 6
use FEEDTHRU  F-1314
transform 1 0 2847 0 1 2796
box 0 0 3 6
<< end >>
