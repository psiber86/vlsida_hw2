magic
tech scmos
timestamp 1395743131
<< m1p >>
use CELL  1
transform -1 0 1946 0 1 1024
box 0 0 6 6
use CELL  2
transform 1 0 1790 0 1 1757
box 0 0 6 6
use CELL  3
transform 1 0 1896 0 1 1393
box 0 0 6 6
use CELL  4
transform 1 0 1730 0 1 971
box 0 0 6 6
use CELL  5
transform 1 0 1945 0 1 1476
box 0 0 6 6
use CELL  6
transform 1 0 1734 0 1 1267
box 0 0 6 6
use CELL  7
transform -1 0 1842 0 -1 1482
box 0 0 6 6
use CELL  8
transform 1 0 1922 0 1 878
box 0 0 6 6
use CELL  9
transform 1 0 1941 0 1 899
box 0 0 6 6
use CELL  10
transform 1 0 1829 0 1 1775
box 0 0 6 6
use CELL  11
transform 1 0 2010 0 1 1476
box 0 0 6 6
use CELL  12
transform 1 0 1887 0 1 1766
box 0 0 6 6
use CELL  13
transform -1 0 1846 0 1 1168
box 0 0 6 6
use CELL  14
transform 1 0 1917 0 1 1537
box 0 0 6 6
use CELL  15
transform 1 0 1737 0 -1 1340
box 0 0 6 6
use CELL  16
transform 1 0 1853 0 -1 1725
box 0 0 6 6
use CELL  17
transform 1 0 1810 0 1 869
box 0 0 6 6
use CELL  18
transform 1 0 1957 0 1 1537
box 0 0 6 6
use CELL  19
transform 1 0 1794 0 1 869
box 0 0 6 6
use CELL  20
transform -1 0 1900 0 -1 1750
box 0 0 6 6
use CELL  21
transform 1 0 1873 0 1 1766
box 0 0 6 6
use CELL  22
transform -1 0 1755 0 1 836
box 0 0 6 6
use CELL  23
transform 1 0 2027 0 1 1267
box 0 0 6 6
use CELL  24
transform -1 0 1756 0 -1 1543
box 0 0 6 6
use CELL  25
transform 1 0 1845 0 1 1775
box 0 0 6 6
use CELL  26
transform 1 0 1804 0 1 1775
box 0 0 6 6
use CELL  27
transform -1 0 1953 0 -1 1030
box 0 0 6 6
use CELL  28
transform 1 0 1934 0 1 899
box 0 0 6 6
use CELL  29
transform 1 0 1913 0 1 971
box 0 0 6 6
use CELL  30
transform 1 0 1762 0 1 1766
box 0 0 6 6
use CELL  31
transform -1 0 1923 0 1 1655
box 0 0 6 6
use CELL  32
transform 1 0 1780 0 1 1537
box 0 0 6 6
use CELL  33
transform 1 0 1790 0 1 1766
box 0 0 6 6
use CELL  34
transform 1 0 1820 0 1 1766
box 0 0 6 6
use CELL  35
transform 1 0 1838 0 1 1766
box 0 0 6 6
use CELL  36
transform -1 0 1734 0 1 1087
box 0 0 6 6
use CELL  37
transform 1 0 1798 0 -1 1482
box 0 0 6 6
use CELL  38
transform -1 0 1711 0 1 1610
box 0 0 6 6
use CELL  39
transform -1 0 1780 0 1 1655
box 0 0 6 6
use CELL  40
transform -1 0 2030 0 -1 1482
box 0 0 6 6
use CELL  41
transform 1 0 1908 0 1 1766
box 0 0 6 6
use CELL  42
transform 1 0 1908 0 1 1744
box 0 0 6 6
use CELL  43
transform 1 0 1844 0 1 878
box 0 0 6 6
use CELL  44
transform -1 0 1952 0 1 1393
box 0 0 6 6
use CELL  45
transform 1 0 1794 0 1 851
box 0 0 6 6
use CELL  46
transform 1 0 1896 0 -1 1704
box 0 0 6 6
use CELL  47
transform 1 0 1741 0 1 1698
box 0 0 6 6
use CELL  48
transform 1 0 1764 0 1 878
box 0 0 6 6
use CELL  49
transform 1 0 1910 0 1 1087
box 0 0 6 6
use CELL  50
transform -1 0 2036 0 1 1393
box 0 0 6 6
use CELL  51
transform -1 0 1830 0 1 836
box 0 0 6 6
use CELL  52
transform -1 0 1856 0 1 928
box 0 0 6 6
use CELL  53
transform -1 0 1926 0 1 971
box 0 0 6 6
use CELL  54
transform 1 0 1794 0 1 878
box 0 0 6 6
use CELL  55
transform -1 0 1743 0 1 1610
box 0 0 6 6
use CELL  56
transform -1 0 1916 0 1 1610
box 0 0 6 6
use CELL  57
transform 1 0 1858 0 1 878
box 0 0 6 6
use CELL  58
transform 1 0 1769 0 1 1766
box 0 0 6 6
use CELL  59
transform -1 0 1800 0 -1 1543
box 0 0 6 6
use CELL  60
transform 1 0 1852 0 1 1757
box 0 0 6 6
use CELL  61
transform -1 0 1909 0 -1 1093
box 0 0 6 6
use CELL  62
transform -1 0 1872 0 1 1393
box 0 0 6 6
use CELL  63
transform 1 0 1710 0 -1 905
box 0 0 6 6
use CELL  64
transform -1 0 1735 0 1 1476
box 0 0 6 6
use CELL  65
transform 1 0 1776 0 1 1766
box 0 0 6 6
use CELL  66
transform 1 0 1808 0 1 1024
box 0 0 6 6
use CELL  67
transform -1 0 1825 0 1 1168
box 0 0 6 6
use CELL  68
transform 1 0 1901 0 1 1757
box 0 0 6 6
use CELL  69
transform 1 0 1901 0 1 1744
box 0 0 6 6
use CELL  70
transform 1 0 1913 0 1 1719
box 0 0 6 6
use CELL  71
transform 1 0 1741 0 1 1719
box 0 0 6 6
use CELL  72
transform 1 0 2010 0 1 1537
box 0 0 6 6
use CELL  73
transform 1 0 1779 0 1 1087
box 0 0 6 6
use CELL  74
transform -1 0 1741 0 -1 1093
box 0 0 6 6
use CELL  75
transform 1 0 1858 0 1 851
box 0 0 6 6
use CELL  76
transform 1 0 1893 0 1 851
box 0 0 6 6
use CELL  77
transform 1 0 1801 0 1 851
box 0 0 6 6
use CELL  78
transform 1 0 1717 0 1 971
box 0 0 6 6
use CELL  79
transform -1 0 1948 0 1 1334
box 0 0 6 6
use CELL  80
transform 1 0 1886 0 1 851
box 0 0 6 6
use CELL  81
transform 1 0 1776 0 1 1757
box 0 0 6 6
use CELL  82
transform 1 0 1785 0 1 851
box 0 0 6 6
use CELL  83
transform 1 0 1965 0 1 1334
box 0 0 6 6
use CELL  84
transform 1 0 1873 0 1 1087
box 0 0 6 6
use CELL  85
transform 1 0 1815 0 1 836
box 0 0 6 6
use CELL  86
transform 1 0 2003 0 1 1537
box 0 0 6 6
use CELL  87
transform -1 0 1775 0 1 1744
box 0 0 6 6
use CELL  88
transform -1 0 1839 0 1 1393
box 0 0 6 6
use CELL  89
transform -1 0 1748 0 1 1024
box 0 0 6 6
use CELL  90
transform 1 0 1680 0 -1 1750
box 0 0 6 6
use CELL  91
transform 1 0 1755 0 1 1744
box 0 0 6 6
use CELL  92
transform 1 0 1847 0 1 1334
box 0 0 6 6
use CELL  93
transform 1 0 1739 0 1 971
box 0 0 6 6
use CELL  94
transform -1 0 1975 0 1 971
box 0 0 6 6
use CELL  95
transform 1 0 1923 0 1 928
box 0 0 6 6
use CELL  96
transform 1 0 1741 0 1 878
box 0 0 6 6
use CELL  97
transform 1 0 1893 0 1 860
box 0 0 6 6
use CELL  98
transform 1 0 1941 0 1 1087
box 0 0 6 6
use CELL  99
transform -1 0 1693 0 -1 1750
box 0 0 6 6
use CELL  100
transform -1 0 1971 0 1 1655
box 0 0 6 6
use CELL  101
transform 1 0 2037 0 -1 1399
box 0 0 6 6
use CELL  102
transform 1 0 1825 0 1 928
box 0 0 6 6
use CELL  103
transform -1 0 1754 0 1 928
box 0 0 6 6
use CELL  104
transform -1 0 1981 0 1 1610
box 0 0 6 6
use CELL  105
transform 1 0 1986 0 -1 1093
box 0 0 6 6
use CELL  106
transform 1 0 1798 0 1 1168
box 0 0 6 6
use CELL  107
transform -1 0 1716 0 -1 977
box 0 0 6 6
use CELL  108
transform 1 0 1819 0 1 860
box 0 0 6 6
use CELL  109
transform 1 0 1887 0 1 1757
box 0 0 6 6
use CELL  110
transform 1 0 1954 0 1 1610
box 0 0 6 6
use CELL  111
transform 1 0 1829 0 1 1757
box 0 0 6 6
use CELL  112
transform -1 0 1869 0 1 1537
box 0 0 6 6
use CELL  113
transform 1 0 1819 0 1 971
box 0 0 6 6
use CELL  114
transform 1 0 1736 0 -1 1543
box 0 0 6 6
use CELL  115
transform -1 0 1812 0 -1 1750
box 0 0 6 6
use CELL  116
transform 1 0 1771 0 1 869
box 0 0 6 6
use CELL  117
transform 1 0 1959 0 -1 1482
box 0 0 6 6
use CELL  118
transform 1 0 1813 0 1 1757
box 0 0 6 6
use CELL  119
transform 1 0 1819 0 1 869
box 0 0 6 6
use CELL  120
transform 1 0 1977 0 1 1393
box 0 0 6 6
use CELL  121
transform 1 0 1968 0 1 1024
box 0 0 6 6
use CELL  122
transform 1 0 1885 0 1 1744
box 0 0 6 6
use CELL  123
transform 1 0 1843 0 1 1744
box 0 0 6 6
use CELL  124
transform 1 0 2028 0 -1 1093
box 0 0 6 6
use CELL  125
transform -1 0 1797 0 -1 1174
box 0 0 6 6
use CELL  126
transform -1 0 1761 0 1 1698
box 0 0 6 6
use CELL  127
transform 1 0 1806 0 1 1719
box 0 0 6 6
use CELL  128
transform 1 0 1760 0 1 928
box 0 0 6 6
use CELL  129
transform -1 0 1909 0 -1 1616
box 0 0 6 6
use CELL  130
transform 1 0 1759 0 1 899
box 0 0 6 6
use CELL  131
transform -1 0 1922 0 -1 934
box 0 0 6 6
use CELL  132
transform -1 0 1797 0 1 836
box 0 0 6 6
use CELL  133
transform 1 0 1851 0 1 878
box 0 0 6 6
use CELL  134
transform 1 0 1827 0 1 1698
box 0 0 6 6
use CELL  135
transform 1 0 1850 0 1 1698
box 0 0 6 6
use CELL  136
transform 1 0 1815 0 1 899
box 0 0 6 6
use CELL  137
transform 1 0 1721 0 1 1610
box 0 0 6 6
use CELL  138
transform 1 0 1787 0 1 899
box 0 0 6 6
use CELL  139
transform -1 0 1779 0 -1 1543
box 0 0 6 6
use CELL  140
transform -1 0 1791 0 -1 842
box 0 0 6 6
use CELL  141
transform 1 0 2022 0 1 1168
box 0 0 6 6
use CELL  142
transform -1 0 1916 0 1 1393
box 0 0 6 6
use CELL  143
transform 1 0 1975 0 1 1024
box 0 0 6 6
use CELL  144
transform -1 0 1917 0 1 1334
box 0 0 6 6
use CELL  145
transform 1 0 1831 0 1 899
box 0 0 6 6
use CELL  146
transform 1 0 1787 0 -1 1273
box 0 0 6 6
use CELL  147
transform -1 0 1800 0 1 1794
box 0 0 6 6
use CELL  148
transform 1 0 1958 0 1 1334
box 0 0 6 6
use CELL  149
transform 1 0 1760 0 1 1334
box 0 0 6 6
use CELL  150
transform 1 0 1770 0 -1 1800
box 0 0 6 6
use CELL  151
transform 1 0 1771 0 1 1267
box 0 0 6 6
use CELL  152
transform -1 0 2056 0 1 1168
box 0 0 6 6
use CELL  153
transform 1 0 1748 0 1 860
box 0 0 6 6
use CELL  154
transform -1 0 1730 0 1 971
box 0 0 6 6
use CELL  155
transform -1 0 1978 0 1 1655
box 0 0 6 6
use CELL  156
transform 1 0 1778 0 1 860
box 0 0 6 6
use CELL  157
transform 1 0 1809 0 1 1087
box 0 0 6 6
use CELL  158
transform 1 0 1769 0 1 1775
box 0 0 6 6
use CELL  159
transform 1 0 1770 0 1 1024
box 0 0 6 6
use CELL  160
transform 1 0 1755 0 1 1775
box 0 0 6 6
use CELL  161
transform -1 0 1822 0 1 1087
box 0 0 6 6
use CELL  162
transform 1 0 1762 0 1 1775
box 0 0 6 6
use CELL  163
transform -1 0 1903 0 -1 934
box 0 0 6 6
use CELL  164
transform 1 0 1866 0 1 928
box 0 0 6 6
use CELL  165
transform 1 0 2031 0 -1 1482
box 0 0 6 6
use CELL  166
transform -1 0 1882 0 -1 1616
box 0 0 6 6
use CELL  167
transform -1 0 1732 0 1 899
box 0 0 6 6
use CELL  168
transform 1 0 1797 0 1 1744
box 0 0 6 6
use CELL  169
transform 1 0 1893 0 1 1334
box 0 0 6 6
use CELL  170
transform -1 0 2000 0 -1 1174
box 0 0 6 6
use CELL  171
transform -1 0 1778 0 1 1087
box 0 0 6 6
use CELL  172
transform -1 0 1750 0 1 1334
box 0 0 6 6
use CELL  173
transform 1 0 1950 0 1 1537
box 0 0 6 6
use CELL  174
transform 1 0 1777 0 1 1024
box 0 0 6 6
use CELL  175
transform 1 0 1820 0 1 1698
box 0 0 6 6
use CELL  176
transform 1 0 1806 0 1 1698
box 0 0 6 6
use CELL  177
transform -1 0 2043 0 -1 1482
box 0 0 6 6
use CELL  178
transform 1 0 1776 0 1 1698
box 0 0 6 6
use CELL  179
transform 1 0 1762 0 1 836
box 0 0 6 6
use CELL  180
transform 1 0 1698 0 1 1610
box 0 0 6 6
use CELL  181
transform -1 0 1934 0 1 1267
box 0 0 6 6
use CELL  182
transform 1 0 1755 0 1 1719
box 0 0 6 6
use CELL  183
transform 1 0 1853 0 1 1655
box 0 0 6 6
use CELL  184
transform 1 0 1820 0 1 1719
box 0 0 6 6
use CELL  185
transform 1 0 1790 0 1 1719
box 0 0 6 6
use CELL  186
transform 1 0 1783 0 1 1719
box 0 0 6 6
use CELL  187
transform -1 0 1742 0 1 1476
box 0 0 6 6
use CELL  188
transform -1 0 1793 0 1 1537
box 0 0 6 6
use CELL  189
transform 1 0 1767 0 1 1655
box 0 0 6 6
use CELL  190
transform 1 0 1894 0 1 1087
box 0 0 6 6
use CELL  191
transform 1 0 1881 0 1 1537
box 0 0 6 6
use CELL  192
transform 1 0 1807 0 1 928
box 0 0 6 6
use CELL  193
transform 1 0 1774 0 1 928
box 0 0 6 6
use CELL  194
transform 1 0 1728 0 -1 1399
box 0 0 6 6
use CELL  195
transform 1 0 1813 0 1 1698
box 0 0 6 6
use CELL  196
transform 1 0 1728 0 1 1024
box 0 0 6 6
use CELL  197
transform 1 0 1869 0 1 1655
box 0 0 6 6
use CELL  198
transform -1 0 1799 0 1 1087
box 0 0 6 6
use CELL  199
transform 1 0 2031 0 -1 1543
box 0 0 6 6
use CELL  200
transform 1 0 1824 0 1 1024
box 0 0 6 6
use CELL  201
transform 1 0 1984 0 1 1393
box 0 0 6 6
use CELL  202
transform 1 0 1862 0 1 1655
box 0 0 6 6
use CELL  203
transform -1 0 1824 0 1 1537
box 0 0 6 6
use CELL  204
transform 1 0 1982 0 1 1024
box 0 0 6 6
use CELL  205
transform 1 0 1776 0 1 1334
box 0 0 6 6
use CELL  206
transform -1 0 1796 0 -1 1340
box 0 0 6 6
use CELL  207
transform 1 0 1762 0 1 971
box 0 0 6 6
use CELL  208
transform 1 0 1834 0 1 928
box 0 0 6 6
use CELL  209
transform -1 0 1830 0 -1 1482
box 0 0 6 6
use CELL  210
transform -1 0 1749 0 1 1476
box 0 0 6 6
use CELL  211
transform -1 0 1770 0 -1 1482
box 0 0 6 6
use CELL  212
transform 1 0 1781 0 1 928
box 0 0 6 6
use CELL  213
transform 1 0 1924 0 -1 1616
box 0 0 6 6
use CELL  214
transform -1 0 1782 0 1 1744
box 0 0 6 6
use CELL  215
transform 1 0 1888 0 1 878
box 0 0 6 6
use CELL  216
transform 1 0 2023 0 -1 1399
box 0 0 6 6
use CELL  217
transform 1 0 1766 0 1 1537
box 0 0 6 6
use CELL  218
transform 1 0 1834 0 1 1698
box 0 0 6 6
use CELL  219
transform -1 0 1824 0 -1 1661
box 0 0 6 6
use CELL  220
transform 1 0 1762 0 1 1719
box 0 0 6 6
use CELL  221
transform 1 0 1769 0 1 1719
box 0 0 6 6
use CELL  222
transform 1 0 1908 0 -1 884
box 0 0 6 6
use CELL  223
transform 1 0 1871 0 -1 1340
box 0 0 6 6
use CELL  224
transform 1 0 1797 0 1 1719
box 0 0 6 6
use CELL  225
transform 1 0 1815 0 -1 1030
box 0 0 6 6
use CELL  226
transform -1 0 1789 0 1 1334
box 0 0 6 6
use CELL  227
transform -1 0 1827 0 1 1794
box 0 0 6 6
use CELL  228
transform 1 0 1936 0 1 1610
box 0 0 6 6
use CELL  229
transform 1 0 1843 0 1 928
box 0 0 6 6
use CELL  230
transform 1 0 1832 0 -1 1661
box 0 0 6 6
use CELL  231
transform 1 0 1762 0 1 1744
box 0 0 6 6
use CELL  232
transform 1 0 1806 0 1 1393
box 0 0 6 6
use CELL  233
transform -1 0 1816 0 -1 1482
box 0 0 6 6
use CELL  234
transform -1 0 1816 0 1 971
box 0 0 6 6
use CELL  235
transform 1 0 1783 0 1 1698
box 0 0 6 6
use CELL  236
transform 1 0 1763 0 -1 1030
box 0 0 6 6
use CELL  237
transform 1 0 1790 0 1 1698
box 0 0 6 6
use CELL  238
transform -1 0 2021 0 -1 1174
box 0 0 6 6
use CELL  239
transform -1 0 1770 0 1 1267
box 0 0 6 6
use CELL  240
transform -1 0 1784 0 1 1267
box 0 0 6 6
use CELL  241
transform 1 0 1843 0 1 1698
box 0 0 6 6
use CELL  242
transform 1 0 1755 0 1 971
box 0 0 6 6
use CELL  243
transform -1 0 1750 0 1 1610
box 0 0 6 6
use CELL  244
transform 1 0 1846 0 1 1655
box 0 0 6 6
use CELL  245
transform 1 0 1839 0 1 1655
box 0 0 6 6
use CELL  246
transform 1 0 1860 0 -1 1482
box 0 0 6 6
use CELL  247
transform 1 0 1722 0 -1 1543
box 0 0 6 6
use CELL  248
transform 1 0 1802 0 1 1655
box 0 0 6 6
use CELL  249
transform 1 0 1838 0 -1 1340
box 0 0 6 6
use CELL  250
transform 1 0 1787 0 1 971
box 0 0 6 6
use CELL  251
transform 1 0 1881 0 1 878
box 0 0 6 6
use CELL  252
transform 1 0 1771 0 1 1476
box 0 0 6 6
use CELL  253
transform -1 0 1735 0 1 1537
box 0 0 6 6
use CELL  254
transform 1 0 1889 0 1 1698
box 0 0 6 6
use CELL  255
transform -1 0 1958 0 1 1168
box 0 0 6 6
use CELL  256
transform 1 0 1878 0 1 899
box 0 0 6 6
use CELL  257
transform 1 0 1885 0 1 899
box 0 0 6 6
use CELL  258
transform 1 0 2036 0 -1 1174
box 0 0 6 6
use CELL  259
transform 1 0 1767 0 1 928
box 0 0 6 6
use CELL  260
transform 1 0 1904 0 1 928
box 0 0 6 6
use CELL  261
transform 1 0 1954 0 1 1024
box 0 0 6 6
use CELL  262
transform 1 0 1999 0 1 1267
box 0 0 6 6
use CELL  263
transform 1 0 1852 0 1 971
box 0 0 6 6
use CELL  264
transform 1 0 1927 0 1 971
box 0 0 6 6
use CELL  265
transform 1 0 1924 0 -1 1174
box 0 0 6 6
use CELL  266
transform -1 0 1923 0 -1 1616
box 0 0 6 6
use CELL  267
transform 1 0 1968 0 1 1610
box 0 0 6 6
use CELL  268
transform 1 0 1800 0 -1 1093
box 0 0 6 6
use CELL  269
transform 1 0 1734 0 1 860
box 0 0 6 6
use CELL  270
transform 1 0 1792 0 1 1393
box 0 0 6 6
use CELL  271
transform -1 0 2063 0 1 1168
box 0 0 6 6
use CELL  272
transform 1 0 1764 0 1 860
box 0 0 6 6
use CELL  273
transform 1 0 1753 0 -1 1661
box 0 0 6 6
use CELL  274
transform 1 0 1784 0 -1 1616
box 0 0 6 6
use CELL  275
transform 1 0 1794 0 1 860
box 0 0 6 6
use CELL  276
transform 1 0 1810 0 1 860
box 0 0 6 6
use CELL  277
transform -1 0 1740 0 1 928
box 0 0 6 6
use CELL  278
transform 1 0 1826 0 1 860
box 0 0 6 6
use CELL  279
transform 1 0 1844 0 1 860
box 0 0 6 6
use CELL  280
transform 1 0 1858 0 1 860
box 0 0 6 6
use CELL  281
transform 1 0 1872 0 1 860
box 0 0 6 6
use CELL  282
transform 1 0 1886 0 1 860
box 0 0 6 6
use CELL  283
transform 1 0 1900 0 1 860
box 0 0 6 6
use CELL  284
transform -1 0 2070 0 1 1168
box 0 0 6 6
use CELL  285
transform -1 0 1805 0 1 899
box 0 0 6 6
use CELL  286
transform 1 0 1754 0 -1 1399
box 0 0 6 6
use CELL  287
transform 1 0 1883 0 1 1719
box 0 0 6 6
use CELL  288
transform 1 0 1890 0 1 1719
box 0 0 6 6
use CELL  289
transform 1 0 1940 0 -1 1273
box 0 0 6 6
use CELL  290
transform 1 0 1843 0 1 1087
box 0 0 6 6
use CELL  291
transform -1 0 1999 0 1 1087
box 0 0 6 6
use CELL  292
transform 1 0 1819 0 1 878
box 0 0 6 6
use CELL  293
transform 1 0 1813 0 1 1744
box 0 0 6 6
use CELL  294
transform 1 0 1757 0 1 878
box 0 0 6 6
use CELL  295
transform 1 0 1771 0 1 878
box 0 0 6 6
use CELL  296
transform 1 0 1785 0 1 878
box 0 0 6 6
use CELL  297
transform 1 0 2034 0 1 1267
box 0 0 6 6
use CELL  298
transform 1 0 1836 0 1 1744
box 0 0 6 6
use CELL  299
transform -1 0 1716 0 1 1794
box 0 0 6 6
use CELL  300
transform 1 0 1797 0 1 1698
box 0 0 6 6
use CELL  301
transform 1 0 1866 0 1 899
box 0 0 6 6
use CELL  302
transform 1 0 1878 0 -1 934
box 0 0 6 6
use CELL  303
transform 1 0 1824 0 1 899
box 0 0 6 6
use CELL  304
transform -1 0 1768 0 1 1698
box 0 0 6 6
use CELL  305
transform 1 0 1813 0 1 1719
box 0 0 6 6
use CELL  306
transform 1 0 1776 0 -1 1725
box 0 0 6 6
use CELL  307
transform 1 0 1773 0 1 899
box 0 0 6 6
use CELL  308
transform 1 0 1780 0 1 899
box 0 0 6 6
use CELL  309
transform 1 0 1803 0 -1 977
box 0 0 6 6
use CELL  310
transform 1 0 1806 0 1 899
box 0 0 6 6
use CELL  311
transform -1 0 1884 0 1 1476
box 0 0 6 6
use CELL  312
transform 1 0 1931 0 1 1655
box 0 0 6 6
use CELL  313
transform 1 0 1854 0 1 899
box 0 0 6 6
use CELL  314
transform 1 0 1933 0 1 1698
box 0 0 6 6
use CELL  315
transform -1 0 1782 0 -1 1399
box 0 0 6 6
use CELL  316
transform -1 0 1757 0 1 1334
box 0 0 6 6
use CELL  317
transform 1 0 1839 0 -1 1725
box 0 0 6 6
use CELL  318
transform 1 0 1867 0 1 878
box 0 0 6 6
use CELL  319
transform -1 0 1772 0 -1 905
box 0 0 6 6
use CELL  320
transform 1 0 1897 0 1 899
box 0 0 6 6
use CELL  321
transform -1 0 1799 0 -1 1030
box 0 0 6 6
use CELL  322
transform 1 0 1945 0 1 1168
box 0 0 6 6
use CELL  323
transform 1 0 1961 0 1 1024
box 0 0 6 6
use CELL  324
transform 1 0 1949 0 -1 1340
box 0 0 6 6
use CELL  325
transform 1 0 1748 0 1 1267
box 0 0 6 6
use CELL  326
transform 1 0 1980 0 1 1476
box 0 0 6 6
use CELL  327
transform 1 0 1801 0 1 878
box 0 0 6 6
use CELL  328
transform 1 0 1979 0 1 1537
box 0 0 6 6
use CELL  329
transform -1 0 1876 0 1 1024
box 0 0 6 6
use CELL  330
transform 1 0 1865 0 1 860
box 0 0 6 6
use CELL  331
transform 1 0 1780 0 1 1476
box 0 0 6 6
use CELL  332
transform 1 0 1820 0 1 1744
box 0 0 6 6
use CELL  333
transform 1 0 1794 0 -1 977
box 0 0 6 6
use CELL  334
transform 1 0 1850 0 1 1744
box 0 0 6 6
use CELL  335
transform 1 0 1871 0 1 1744
box 0 0 6 6
use CELL  336
transform 1 0 1878 0 1 1744
box 0 0 6 6
use CELL  337
transform 1 0 1722 0 -1 1482
box 0 0 6 6
use CELL  338
transform 1 0 1879 0 1 869
box 0 0 6 6
use CELL  339
transform 1 0 1835 0 1 860
box 0 0 6 6
use CELL  340
transform 1 0 1851 0 1 860
box 0 0 6 6
use CELL  341
transform -1 0 1891 0 -1 1482
box 0 0 6 6
use CELL  342
transform 1 0 1806 0 -1 1543
box 0 0 6 6
use CELL  343
transform 1 0 1962 0 1 971
box 0 0 6 6
use CELL  344
transform -1 0 1805 0 -1 1399
box 0 0 6 6
use CELL  345
transform -1 0 1776 0 -1 1174
box 0 0 6 6
use CELL  346
transform 1 0 1757 0 1 869
box 0 0 6 6
use CELL  347
transform -1 0 1860 0 1 1024
box 0 0 6 6
use CELL  348
transform 1 0 1785 0 1 869
box 0 0 6 6
use CELL  349
transform 1 0 1801 0 1 869
box 0 0 6 6
use CELL  350
transform 1 0 1749 0 -1 1174
box 0 0 6 6
use CELL  351
transform 1 0 1835 0 1 869
box 0 0 6 6
use CELL  352
transform 1 0 1851 0 1 869
box 0 0 6 6
use CELL  353
transform 1 0 1865 0 1 869
box 0 0 6 6
use CELL  354
transform 1 0 1835 0 1 878
box 0 0 6 6
use CELL  355
transform -1 0 1909 0 -1 1399
box 0 0 6 6
use CELL  356
transform 1 0 1747 0 1 899
box 0 0 6 6
use CELL  357
transform 1 0 1904 0 1 899
box 0 0 6 6
use CELL  358
transform 1 0 1746 0 1 971
box 0 0 6 6
use CELL  359
transform 1 0 1934 0 1 971
box 0 0 6 6
use CELL  360
transform 1 0 1934 0 1 1087
box 0 0 6 6
use CELL  361
transform 1 0 1842 0 -1 1030
box 0 0 6 6
use CELL  362
transform 1 0 2029 0 1 1168
box 0 0 6 6
use CELL  363
transform 1 0 1748 0 1 1698
box 0 0 6 6
use CELL  364
transform 1 0 1998 0 1 1476
box 0 0 6 6
use CELL  365
transform 1 0 1757 0 1 1537
box 0 0 6 6
use CELL  366
transform -1 0 1750 0 1 1087
box 0 0 6 6
use CELL  367
transform 1 0 2014 0 1 1087
box 0 0 6 6
use CELL  368
transform 1 0 1783 0 1 1757
box 0 0 6 6
use CELL  369
transform 1 0 1797 0 1 1757
box 0 0 6 6
use CELL  370
transform 1 0 1840 0 1 971
box 0 0 6 6
use CELL  371
transform 1 0 1845 0 1 1757
box 0 0 6 6
use CELL  372
transform 1 0 1868 0 1 1267
box 0 0 6 6
use CELL  373
transform -1 0 1753 0 1 1393
box 0 0 6 6
use CELL  374
transform 1 0 1781 0 1 1655
box 0 0 6 6
use CELL  375
transform 1 0 1972 0 1 1334
box 0 0 6 6
use CELL  376
transform -1 0 1749 0 1 1537
box 0 0 6 6
use CELL  377
transform 1 0 1813 0 1 1766
box 0 0 6 6
use CELL  378
transform 1 0 1984 0 1 1267
box 0 0 6 6
use CELL  379
transform 1 0 1757 0 1 860
box 0 0 6 6
use CELL  380
transform -1 0 1778 0 1 1610
box 0 0 6 6
use CELL  381
transform 1 0 1771 0 1 860
box 0 0 6 6
use CELL  382
transform 1 0 1785 0 1 860
box 0 0 6 6
use CELL  383
transform 1 0 1741 0 1 928
box 0 0 6 6
use CELL  384
transform -1 0 1817 0 -1 1661
box 0 0 6 6
use CELL  385
transform 1 0 1895 0 1 878
box 0 0 6 6
use CELL  386
transform 1 0 1733 0 -1 905
box 0 0 6 6
use CELL  387
transform -1 0 1832 0 1 1267
box 0 0 6 6
use CELL  388
transform 1 0 2043 0 1 1168
box 0 0 6 6
use CELL  389
transform 1 0 1901 0 1 971
box 0 0 6 6
use CELL  390
transform 1 0 1783 0 1 1393
box 0 0 6 6
use CELL  391
transform 1 0 1897 0 1 1719
box 0 0 6 6
use CELL  392
transform -1 0 1904 0 1 1267
box 0 0 6 6
use CELL  393
transform 1 0 1769 0 1 971
box 0 0 6 6
use CELL  394
transform 1 0 1751 0 1 1024
box 0 0 6 6
use CELL  395
transform 1 0 1921 0 -1 1482
box 0 0 6 6
use CELL  396
transform 1 0 1741 0 1 860
box 0 0 6 6
use CELL  397
transform 1 0 1879 0 1 860
box 0 0 6 6
use CELL  398
transform -1 0 1757 0 1 1087
box 0 0 6 6
use CELL  399
transform 1 0 1741 0 1 869
box 0 0 6 6
use CELL  400
transform 1 0 1893 0 1 869
box 0 0 6 6
use CELL  401
transform 1 0 1692 0 1 1537
box 0 0 6 6
use CELL  402
transform 1 0 1801 0 1 860
box 0 0 6 6
use CELL  403
transform 1 0 2002 0 1 1393
box 0 0 6 6
use CELL  404
transform -1 0 1930 0 1 1655
box 0 0 6 6
use CELL  405
transform -1 0 1831 0 1 1655
box 0 0 6 6
use CELL  406
transform 1 0 1927 0 1 899
box 0 0 6 6
use CELL  407
transform 1 0 1941 0 1 971
box 0 0 6 6
use CELL  408
transform 1 0 1769 0 1 1757
box 0 0 6 6
use CELL  409
transform 1 0 1741 0 1 1267
box 0 0 6 6
use CELL  410
transform 1 0 1874 0 -1 884
box 0 0 6 6
use CELL  411
transform 1 0 2020 0 1 1267
box 0 0 6 6
use CELL  412
transform -1 0 1935 0 -1 1543
box 0 0 6 6
use CELL  413
transform -1 0 2006 0 1 1087
box 0 0 6 6
use CELL  414
transform -1 0 1789 0 1 1744
box 0 0 6 6
use CELL  415
transform 1 0 1740 0 1 899
box 0 0 6 6
use CELL  416
transform 1 0 1873 0 1 1757
box 0 0 6 6
use CELL  417
transform 1 0 1741 0 1 1655
box 0 0 6 6
use CELL  418
transform 1 0 1906 0 1 1719
box 0 0 6 6
use CELL  419
transform -1 0 1833 0 -1 1725
box 0 0 6 6
use CELL  420
transform -1 0 1961 0 1 971
box 0 0 6 6
use CELL  421
transform 1 0 1769 0 1 1393
box 0 0 6 6
use CELL  422
transform -1 0 1958 0 -1 1482
box 0 0 6 6
use CELL  423
transform 1 0 1748 0 1 1744
box 0 0 6 6
use CELL  424
transform 1 0 1755 0 1 1757
box 0 0 6 6
use CELL  425
transform 1 0 1812 0 1 1794
box 0 0 6 6
use CELL  426
transform -1 0 1844 0 1 899
box 0 0 6 6
use CELL  427
transform -1 0 1865 0 -1 977
box 0 0 6 6
use CELL  428
transform 1 0 1762 0 1 1757
box 0 0 6 6
use CELL  429
transform 1 0 1748 0 1 1757
box 0 0 6 6
use CELL  430
transform 1 0 1872 0 1 851
box 0 0 6 6
use CELL  431
transform 1 0 1879 0 1 851
box 0 0 6 6
use CELL  432
transform -1 0 1869 0 1 1024
box 0 0 6 6
use CELL  433
transform -1 0 1748 0 1 1168
box 0 0 6 6
use CELL  434
transform 1 0 1865 0 1 851
box 0 0 6 6
use CELL  435
transform 1 0 1778 0 1 851
box 0 0 6 6
use CELL  436
transform 1 0 1900 0 1 851
box 0 0 6 6
use CELL  437
transform -1 0 1766 0 1 1655
box 0 0 6 6
use CELL  438
transform 1 0 1947 0 -1 1661
box 0 0 6 6
use CELL  439
transform -1 0 1896 0 1 928
box 0 0 6 6
use CELL  440
transform 1 0 1851 0 1 851
box 0 0 6 6
use CELL  441
transform 1 0 1844 0 1 851
box 0 0 6 6
use CELL  442
transform 1 0 1826 0 1 851
box 0 0 6 6
use CELL  443
transform 1 0 1835 0 1 851
box 0 0 6 6
use CELL  444
transform 1 0 1800 0 1 1610
box 0 0 6 6
use CELL  445
transform 1 0 1948 0 1 971
box 0 0 6 6
use CELL  446
transform 1 0 1710 0 1 1719
box 0 0 6 6
use CELL  447
transform 1 0 1771 0 1 851
box 0 0 6 6
use CELL  448
transform 1 0 1845 0 1 1766
box 0 0 6 6
use CELL  449
transform 1 0 1961 0 1 1610
box 0 0 6 6
use CELL  450
transform 1 0 1919 0 1 1698
box 0 0 6 6
use CELL  451
transform -1 0 1723 0 1 899
box 0 0 6 6
use CELL  452
transform -1 0 1892 0 1 1334
box 0 0 6 6
use CELL  453
transform 1 0 1741 0 1 1744
box 0 0 6 6
use CELL  454
transform 1 0 1818 0 1 1610
box 0 0 6 6
use CELL  455
transform 1 0 1741 0 1 1757
box 0 0 6 6
use CELL  456
transform -1 0 1794 0 1 928
box 0 0 6 6
use CELL  457
transform 1 0 1799 0 1 1334
box 0 0 6 6
use CELL  458
transform 1 0 1757 0 1 1476
box 0 0 6 6
use CELL  459
transform -1 0 2012 0 -1 1273
box 0 0 6 6
use CELL  460
transform 1 0 1804 0 1 1757
box 0 0 6 6
use CELL  461
transform 1 0 2021 0 -1 1093
box 0 0 6 6
use CELL  462
transform 1 0 1783 0 1 1766
box 0 0 6 6
use CELL  463
transform 1 0 1797 0 1 1766
box 0 0 6 6
use CELL  464
transform 1 0 1829 0 1 1766
box 0 0 6 6
use CELL  465
transform 1 0 1894 0 1 1757
box 0 0 6 6
use CELL  466
transform -1 0 1763 0 1 1267
box 0 0 6 6
use CELL  467
transform 1 0 1827 0 1 1537
box 0 0 6 6
use CELL  468
transform -1 0 1811 0 -1 1174
box 0 0 6 6
use CELL  469
transform 1 0 1880 0 1 1757
box 0 0 6 6
use CELL  470
transform 1 0 1716 0 -1 1340
box 0 0 6 6
use CELL  471
transform 1 0 1838 0 1 1757
box 0 0 6 6
use CELL  472
transform 1 0 1981 0 1 1334
box 0 0 6 6
use CELL  473
transform 1 0 1820 0 1 1757
box 0 0 6 6
use CELL  474
transform 1 0 1911 0 -1 905
box 0 0 6 6
use CELL  475
transform 1 0 1826 0 1 878
box 0 0 6 6
use CELL  476
transform -1 0 1909 0 1 1698
box 0 0 6 6
use CELL  477
transform 1 0 1769 0 1 1334
box 0 0 6 6
use CELL  478
transform 1 0 1786 0 1 1024
box 0 0 6 6
use CELL  479
transform 1 0 1756 0 1 836
box 0 0 6 6
use CELL  480
transform 1 0 1748 0 1 1719
box 0 0 6 6
use CELL  481
transform 1 0 1831 0 1 971
box 0 0 6 6
use CELL  482
transform -1 0 1983 0 1 1267
box 0 0 6 6
use CELL  483
transform -1 0 1918 0 -1 1704
box 0 0 6 6
use CELL  484
transform 1 0 1765 0 1 1610
box 0 0 6 6
use CELL  485
transform 1 0 1748 0 1 878
box 0 0 6 6
use CELL  486
transform 1 0 1810 0 1 878
box 0 0 6 6
use CELL  487
transform -1 0 1833 0 1 1744
box 0 0 6 6
use CELL  488
transform 1 0 1730 0 1 1610
box 0 0 6 6
use CELL  489
transform -1 0 1723 0 1 1794
box 0 0 6 6
use CELL  490
transform 1 0 1757 0 1 851
box 0 0 6 6
use CELL  491
transform 1 0 1712 0 1 1610
box 0 0 6 6
use CELL  492
transform 1 0 1764 0 1 851
box 0 0 6 6
use CELL  493
transform 1 0 1970 0 -1 1399
box 0 0 6 6
use CELL  494
transform -1 0 1865 0 -1 934
box 0 0 6 6
use CELL  495
transform 1 0 1735 0 1 1168
box 0 0 6 6
use CELL  496
transform 1 0 1741 0 1 1775
box 0 0 6 6
use CELL  497
transform 1 0 1748 0 1 1775
box 0 0 6 6
use CELL  498
transform -1 0 2030 0 -1 1543
box 0 0 6 6
use CELL  499
transform 1 0 1776 0 1 1775
box 0 0 6 6
use CELL  500
transform -1 0 1921 0 1 878
box 0 0 6 6
use CELL  501
transform -1 0 1729 0 1 1334
box 0 0 6 6
use CELL  502
transform 1 0 1894 0 1 1766
box 0 0 6 6
use CELL  503
transform 1 0 1880 0 1 1766
box 0 0 6 6
use CELL  504
transform 1 0 1852 0 1 1766
box 0 0 6 6
use CELL  505
transform -1 0 2023 0 1 1537
box 0 0 6 6
use CELL  506
transform -1 0 1946 0 1 1655
box 0 0 6 6
use CELL  507
transform 1 0 1989 0 1 1024
box 0 0 6 6
use CELL  508
transform 1 0 1803 0 1 1794
box 0 0 6 6
use CELL  509
transform 1 0 1967 0 -1 1174
box 0 0 6 6
use CELL  510
transform 1 0 1741 0 1 1766
box 0 0 6 6
use CELL  511
transform -1 0 1849 0 1 1610
box 0 0 6 6
use CELL  512
transform -1 0 1734 0 -1 1174
box 0 0 6 6
use CELL  513
transform 1 0 1844 0 1 1267
box 0 0 6 6
use CELL  514
transform -1 0 1953 0 1 1267
box 0 0 6 6
use CELL  515
transform 1 0 1847 0 -1 905
box 0 0 6 6
use CELL  516
transform 1 0 1748 0 1 1766
box 0 0 6 6
use CELL  517
transform 1 0 1734 0 1 1766
box 0 0 6 6
use CELL  518
transform 1 0 1988 0 1 1334
box 0 0 6 6
use CELL  519
transform 1 0 1798 0 1 836
box 0 0 6 6
use CELL  520
transform 1 0 1742 0 1 836
box 0 0 6 6
use CELL  521
transform 1 0 1735 0 1 836
box 0 0 6 6
use CELL  522
transform 1 0 1728 0 1 836
box 0 0 6 6
use CELL  523
transform -1 0 1943 0 1 928
box 0 0 6 6
use CELL  524
transform 1 0 1804 0 1 1766
box 0 0 6 6
use CELL  525
transform 1 0 1783 0 1 1775
box 0 0 6 6
use CELL  526
transform 1 0 1790 0 1 1775
box 0 0 6 6
use CELL  527
transform 1 0 1797 0 1 1775
box 0 0 6 6
use CELL  528
transform 1 0 1877 0 -1 1030
box 0 0 6 6
use CELL  529
transform 1 0 1735 0 -1 1399
box 0 0 6 6
use CELL  530
transform 1 0 1888 0 1 1610
box 0 0 6 6
use CELL  531
transform 1 0 1734 0 1 869
box 0 0 6 6
use CELL  532
transform 1 0 1900 0 1 869
box 0 0 6 6
use CELL  533
transform -1 0 1818 0 -1 1174
box 0 0 6 6
use CELL  534
transform 1 0 1735 0 1 1024
box 0 0 6 6
use CELL  535
transform 1 0 1857 0 1 1393
box 0 0 6 6
use CELL  536
transform 1 0 1734 0 1 1775
box 0 0 6 6
use CELL  537
transform -1 0 1852 0 1 1719
box 0 0 6 6
use CELL  538
transform 1 0 2017 0 1 1476
box 0 0 6 6
use CELL  539
transform 1 0 1756 0 1 1168
box 0 0 6 6
use CELL  540
transform 1 0 1734 0 1 1655
box 0 0 6 6
use CELL  541
transform 1 0 1926 0 1 1698
box 0 0 6 6
use CELL  542
transform 1 0 1793 0 1 1610
box 0 0 6 6
use CELL  543
transform 1 0 1734 0 1 1719
box 0 0 6 6
use CELL  544
transform 1 0 1920 0 1 1719
box 0 0 6 6
use CELL  545
transform 1 0 1734 0 1 1744
box 0 0 6 6
use CELL  546
transform 1 0 1734 0 1 1757
box 0 0 6 6
use CELL  547
transform 1 0 1908 0 1 1757
box 0 0 6 6
use CELL  548
transform 1 0 1769 0 1 1698
box 0 0 6 6
use CELL  549
transform -1 0 2013 0 -1 1093
box 0 0 6 6
use CELL  550
transform 1 0 1748 0 1 869
box 0 0 6 6
use CELL  551
transform 1 0 1764 0 1 869
box 0 0 6 6
use CELL  552
transform 1 0 1778 0 1 869
box 0 0 6 6
use CELL  553
transform -1 0 1829 0 -1 1340
box 0 0 6 6
use CELL  554
transform 1 0 1786 0 -1 1093
box 0 0 6 6
use CELL  555
transform -1 0 1769 0 1 1168
box 0 0 6 6
use CELL  556
transform 1 0 1750 0 -1 1482
box 0 0 6 6
use CELL  557
transform -1 0 1764 0 -1 1800
box 0 0 6 6
use CELL  558
transform 1 0 1826 0 1 869
box 0 0 6 6
use CELL  559
transform 1 0 1844 0 1 869
box 0 0 6 6
use CELL  560
transform -1 0 1722 0 1 878
box 0 0 6 6
use CELL  561
transform 1 0 1858 0 1 869
box 0 0 6 6
use CELL  562
transform 1 0 1872 0 1 869
box 0 0 6 6
use CELL  563
transform 1 0 1805 0 1 1267
box 0 0 6 6
use CELL  564
transform -1 0 1964 0 1 1393
box 0 0 6 6
use CELL  565
transform 1 0 1901 0 1 1766
box 0 0 6 6
use CELL  566
transform 1 0 1819 0 1 851
box 0 0 6 6
use CELL  567
transform 1 0 1813 0 1 1775
box 0 0 6 6
use CELL  568
transform 1 0 1734 0 1 851
box 0 0 6 6
use CELL  569
transform 1 0 1741 0 1 851
box 0 0 6 6
use CELL  570
transform 1 0 1748 0 1 851
box 0 0 6 6
use CELL  571
transform 1 0 1778 0 1 878
box 0 0 6 6
use CELL  572
transform 1 0 1755 0 1 1766
box 0 0 6 6
use CELL  573
transform 1 0 1817 0 1 1476
box 0 0 6 6
use CELL  574
transform 1 0 1886 0 1 869
box 0 0 6 6
use CELL  575
transform 1 0 1778 0 1 971
box 0 0 6 6
use CELL  576
transform 1 0 1838 0 1 1775
box 0 0 6 6
use CELL  577
transform 1 0 1918 0 1 899
box 0 0 6 6
use CELL  578
transform -1 0 1842 0 1 1610
box 0 0 6 6
use CELL  579
transform -1 0 1757 0 1 1610
box 0 0 6 6
use CELL  580
transform 1 0 1852 0 1 1775
box 0 0 6 6
use CELL  581
transform 1 0 1873 0 1 1775
box 0 0 6 6
use CELL  582
transform 1 0 1880 0 1 1775
box 0 0 6 6
use CELL  583
transform 1 0 1887 0 1 1775
box 0 0 6 6
use CELL  584
transform 1 0 1894 0 1 1775
box 0 0 6 6
use CELL  585
transform 1 0 1901 0 1 1775
box 0 0 6 6
use CELL  586
transform 1 0 1908 0 1 1775
box 0 0 6 6
use CELL  587
transform 1 0 1810 0 1 851
box 0 0 6 6
use CELL  588
transform 1 0 1820 0 1 1775
box 0 0 6 6
use CELL  589
transform 1 0 1730 0 1 1334
box 0 0 6 6
use CELL  590
transform 1 0 1734 0 1 1698
box 0 0 6 6
use CELL  591
transform -1 0 2019 0 -1 1273
box 0 0 6 6
use CELL  592
transform 1 0 1959 0 1 1655
box 0 0 6 6
use CELL  593
transform -1 0 1970 0 -1 1543
box 0 0 6 6
use CELL  594
transform -1 0 1764 0 1 1610
box 0 0 6 6
use CELL  595
transform 1 0 1790 0 -1 1750
box 0 0 6 6
use CELL  596
transform 1 0 1930 0 1 928
box 0 0 6 6
use CELL  597
transform -1 0 1941 0 1 1334
box 0 0 6 6
use CELL  598
transform 1 0 1902 0 1 878
box 0 0 6 6
use CELL  599
transform 1 0 1734 0 1 878
box 0 0 6 6
use CELL  600
transform 1 0 1800 0 -1 934
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 1889 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 1871 0 1 971
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 1933 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 1857 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 1857 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 1824 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 1943 0 1 928
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 1900 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 1888 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 1897 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 1763 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 1891 0 1 1744
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 1903 0 1 1719
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 1909 0 1 1698
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 1937 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 1933 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 1985 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 1971 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 1996 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 1754 0 1 851
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 1754 0 1 860
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 1754 0 1 869
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 1754 0 1 878
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 1756 0 1 899
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 1757 0 1 928
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 1752 0 1 971
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 1760 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 1757 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 1788 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 1754 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 1757 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 1766 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 1889 0 1 971
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 1884 0 1 928
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 1872 0 1 899
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 1864 0 1 878
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 1924 0 1 899
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 1916 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 1971 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 2000 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 1883 0 1 1698
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 1871 0 1 1719
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 1862 0 1 1744
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 1864 0 1 1757
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 1864 0 1 1766
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 1864 0 1 1775
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 1836 0 1 1794
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 1741 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 1800 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 1790 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 1808 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 1718 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 1799 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 1796 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 2004 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 1877 0 1 1719
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 1868 0 1 1744
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 1870 0 1 1757
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 1870 0 1 1766
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 1870 0 1 1775
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 1839 0 1 1794
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 2017 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 2020 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 1978 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 1821 0 1 836
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 1841 0 1 851
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 1841 0 1 860
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 1841 0 1 869
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 1841 0 1 878
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 1844 0 1 899
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 1895 0 1 971
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 1922 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 1977 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 2009 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 1993 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 1894 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 1812 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 1930 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 1910 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 1880 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 1854 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 1860 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 1723 0 1 899
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 1870 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 1971 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 2003 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 1974 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 1919 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 1892 0 1 971
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 1812 0 1 836
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 1832 0 1 851
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 1832 0 1 860
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 1832 0 1 869
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 1832 0 1 878
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 1988 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 1974 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 1999 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 1955 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 1990 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 2006 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 1983 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 1928 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 1769 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 1849 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 1757 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 1766 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 1782 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 2008 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-109
transform 1 0 2007 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-110
transform 1 0 1997 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-111
transform 1 0 1948 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-112
transform 1 0 1986 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-113
transform 1 0 2000 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-114
transform 1 0 1951 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-115
transform 1 0 1953 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-116
transform 1 0 1953 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-117
transform 1 0 1973 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-118
transform 1 0 1974 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-119
transform 1 0 1923 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-120
transform 1 0 1964 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-121
transform 1 0 1936 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-122
transform 1 0 1938 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-123
transform 1 0 1897 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-124
transform 1 0 1899 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-125
transform 1 0 1886 0 1 1698
box 0 0 3 6
use FEEDTHRU  F-126
transform 1 0 1874 0 1 1719
box 0 0 3 6
use FEEDTHRU  F-127
transform 1 0 1865 0 1 1744
box 0 0 3 6
use FEEDTHRU  F-128
transform 1 0 1867 0 1 1757
box 0 0 3 6
use FEEDTHRU  F-129
transform 1 0 1867 0 1 1766
box 0 0 3 6
use FEEDTHRU  F-130
transform 1 0 1867 0 1 1775
box 0 0 3 6
use FEEDTHRU  F-131
transform 1 0 1879 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-132
transform 1 0 1827 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-133
transform 1 0 1810 0 1 1757
box 0 0 3 6
use FEEDTHRU  F-134
transform 1 0 1810 0 1 1766
box 0 0 3 6
use FEEDTHRU  F-135
transform 1 0 1810 0 1 1775
box 0 0 3 6
use FEEDTHRU  F-136
transform 1 0 1800 0 1 1794
box 0 0 3 6
use FEEDTHRU  F-137
transform 1 0 1944 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-138
transform 1 0 1828 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-139
transform 1 0 1870 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-140
transform 1 0 1911 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-141
transform 1 0 1897 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-142
transform 1 0 1934 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-143
transform 1 0 1816 0 1 851
box 0 0 3 6
use FEEDTHRU  F-144
transform 1 0 1816 0 1 860
box 0 0 3 6
use FEEDTHRU  F-145
transform 1 0 1816 0 1 869
box 0 0 3 6
use FEEDTHRU  F-146
transform 1 0 1816 0 1 878
box 0 0 3 6
use FEEDTHRU  F-147
transform 1 0 1821 0 1 899
box 0 0 3 6
use FEEDTHRU  F-148
transform 1 0 1831 0 1 928
box 0 0 3 6
use FEEDTHRU  F-149
transform 1 0 1750 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-150
transform 1 0 1722 0 1 1698
box 0 0 3 6
use FEEDTHRU  F-151
transform 1 0 1719 0 1 1719
box 0 0 3 6
use FEEDTHRU  F-152
transform 1 0 1781 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-153
transform 1 0 1782 0 1 836
box 0 0 3 6
use FEEDTHRU  F-154
transform 1 0 1807 0 1 851
box 0 0 3 6
use FEEDTHRU  F-155
transform 1 0 1807 0 1 860
box 0 0 3 6
use FEEDTHRU  F-156
transform 1 0 1807 0 1 869
box 0 0 3 6
use FEEDTHRU  F-157
transform 1 0 1807 0 1 878
box 0 0 3 6
use FEEDTHRU  F-158
transform 1 0 1812 0 1 899
box 0 0 3 6
use FEEDTHRU  F-159
transform 1 0 1822 0 1 928
box 0 0 3 6
use FEEDTHRU  F-160
transform 1 0 1934 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-161
transform 1 0 1910 0 1 971
box 0 0 3 6
use FEEDTHRU  F-162
transform 1 0 1910 0 1 928
box 0 0 3 6
use FEEDTHRU  F-163
transform 1 0 1891 0 1 899
box 0 0 3 6
use FEEDTHRU  F-164
transform 1 0 1937 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-165
transform 1 0 1900 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-166
transform 1 0 1914 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-167
transform 1 0 1873 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-168
transform 1 0 1841 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-169
transform 1 0 1858 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-170
transform 1 0 1885 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-171
transform 1 0 1873 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-172
transform 1 0 1859 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-173
transform 1 0 1835 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-174
transform 1 0 1854 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-175
transform 1 0 1842 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-176
transform 1 0 1824 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-177
transform 1 0 1898 0 1 971
box 0 0 3 6
use FEEDTHRU  F-178
transform 1 0 1925 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-179
transform 1 0 1980 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-180
transform 1 0 2012 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-181
transform 1 0 1996 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-182
transform 1 0 1929 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-183
transform 1 0 1952 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-184
transform 1 0 1927 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-185
transform 1 0 1947 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-186
transform 1 0 1882 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-187
transform 1 0 1911 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-188
transform 1 0 1754 0 1 928
box 0 0 3 6
use FEEDTHRU  F-189
transform 1 0 1736 0 1 971
box 0 0 3 6
use FEEDTHRU  F-190
transform 1 0 1748 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-191
transform 1 0 1753 0 1 899
box 0 0 3 6
use FEEDTHRU  F-192
transform 1 0 1803 0 1 1744
box 0 0 3 6
use FEEDTHRU  F-193
transform 1 0 1825 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-194
transform 1 0 1977 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-195
transform 1 0 1976 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-196
transform 1 0 1930 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-197
transform 1 0 1956 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-198
transform 1 0 1791 0 1 851
box 0 0 3 6
use FEEDTHRU  F-199
transform 1 0 1791 0 1 860
box 0 0 3 6
use FEEDTHRU  F-200
transform 1 0 1791 0 1 869
box 0 0 3 6
use FEEDTHRU  F-201
transform 1 0 1791 0 1 878
box 0 0 3 6
use FEEDTHRU  F-202
transform 1 0 1796 0 1 899
box 0 0 3 6
use FEEDTHRU  F-203
transform 1 0 1794 0 1 928
box 0 0 3 6
use FEEDTHRU  F-204
transform 1 0 1775 0 1 971
box 0 0 3 6
use FEEDTHRU  F-205
transform 1 0 1783 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-206
transform 1 0 1806 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-207
transform 1 0 1837 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-208
transform 1 0 1913 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-209
transform 1 0 1760 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-210
transform 1 0 1830 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-211
transform 1 0 1851 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-212
transform 1 0 1832 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-213
transform 1 0 1811 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-214
transform 1 0 1861 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-215
transform 1 0 1852 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-216
transform 1 0 1802 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-217
transform 1 0 1915 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-218
transform 1 0 1892 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-219
transform 1 0 1799 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-220
transform 1 0 1839 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-221
transform 1 0 1867 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-222
transform 1 0 1894 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-223
transform 1 0 1865 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-224
transform 1 0 1844 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-225
transform 1 0 1863 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-226
transform 1 0 1851 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-227
transform 1 0 1845 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-228
transform 1 0 1812 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-229
transform 1 0 1848 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-230
transform 1 0 1815 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-231
transform 1 0 1931 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-232
transform 1 0 1907 0 1 971
box 0 0 3 6
use FEEDTHRU  F-233
transform 1 0 1913 0 1 928
box 0 0 3 6
use FEEDTHRU  F-234
transform 1 0 1894 0 1 899
box 0 0 3 6
use FEEDTHRU  F-235
transform 1 0 1829 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-236
transform 1 0 1842 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-237
transform 1 0 1807 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-238
transform 1 0 1792 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-239
transform 1 0 1830 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-240
transform 1 0 1814 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-241
transform 1 0 1803 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-242
transform 1 0 1778 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-243
transform 1 0 1793 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-244
transform 1 0 1914 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-245
transform 1 0 1877 0 1 1698
box 0 0 3 6
use FEEDTHRU  F-246
transform 1 0 1942 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-247
transform 1 0 1935 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-248
transform 1 0 1803 0 1 1698
box 0 0 3 6
use FEEDTHRU  F-249
transform 1 0 1803 0 1 1719
box 0 0 3 6
use FEEDTHRU  F-250
transform 1 0 1818 0 1 1794
box 0 0 3 6
use FEEDTHRU  F-251
transform 1 0 1835 0 1 1775
box 0 0 3 6
use FEEDTHRU  F-252
transform 1 0 1835 0 1 1766
box 0 0 3 6
use FEEDTHRU  F-253
transform 1 0 1835 0 1 1757
box 0 0 3 6
use FEEDTHRU  F-254
transform 1 0 1833 0 1 1744
box 0 0 3 6
use FEEDTHRU  F-255
transform 1 0 1934 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-256
transform 1 0 1926 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-257
transform 1 0 1967 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-258
transform 1 0 1939 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-259
transform 1 0 1941 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-260
transform 1 0 1900 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-261
transform 1 0 1902 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-262
transform 1 0 1856 0 1 1698
box 0 0 3 6
use FEEDTHRU  F-263
transform 1 0 1961 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-264
transform 1 0 1947 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-265
transform 1 0 1898 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-266
transform 1 0 1820 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-267
transform 1 0 1823 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-268
transform 1 0 1878 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-269
transform 1 0 1859 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-270
transform 1 0 1895 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-271
transform 1 0 1918 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-272
transform 1 0 1888 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-273
transform 1 0 1848 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-274
transform 1 0 1825 0 1 971
box 0 0 3 6
use FEEDTHRU  F-275
transform 1 0 1840 0 1 928
box 0 0 3 6
use FEEDTHRU  F-276
transform 1 0 1862 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-277
transform 1 0 1921 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-278
transform 1 0 1900 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-279
transform 1 0 1880 0 1 971
box 0 0 3 6
use FEEDTHRU  F-280
transform 1 0 1893 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-281
transform 1 0 1903 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-282
transform 1 0 1922 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-283
transform 1 0 1899 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-284
transform 1 0 1916 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-285
transform 1 0 1933 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-286
transform 1 0 1916 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-287
transform 1 0 1883 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-288
transform 1 0 1865 0 1 971
box 0 0 3 6
use FEEDTHRU  F-289
transform 1 0 1887 0 1 928
box 0 0 3 6
use FEEDTHRU  F-290
transform 1 0 1875 0 1 899
box 0 0 3 6
use FEEDTHRU  F-291
transform 1 0 1837 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-292
transform 1 0 1839 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-293
transform 1 0 1833 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-294
transform 1 0 1815 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-295
transform 1 0 1959 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-296
transform 1 0 1962 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-297
transform 1 0 1985 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-298
transform 1 0 1819 0 1 928
box 0 0 3 6
use FEEDTHRU  F-299
transform 1 0 1800 0 1 971
box 0 0 3 6
use FEEDTHRU  F-300
transform 1 0 1821 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-301
transform 1 0 1855 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-302
transform 1 0 1882 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-303
transform 1 0 1836 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-304
transform 1 0 1816 0 1 971
box 0 0 3 6
use FEEDTHRU  F-305
transform 1 0 1922 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-306
transform 1 0 1939 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-307
transform 1 0 1922 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-308
transform 1 0 1932 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-309
transform 1 0 1955 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-310
transform 1 0 1930 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-311
transform 1 0 1899 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-312
transform 1 0 1885 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-313
transform 1 0 1887 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-314
transform 1 0 1880 0 1 1698
box 0 0 3 6
use FEEDTHRU  F-315
transform 1 0 1880 0 1 1719
box 0 0 3 6
use FEEDTHRU  F-316
transform 1 0 1866 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-317
transform 1 0 1884 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-318
transform 1 0 1883 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-319
transform 1 0 1886 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-320
transform 1 0 1893 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-321
transform 1 0 1833 0 1 1719
box 0 0 3 6
use FEEDTHRU  F-322
transform 1 0 1793 0 1 899
box 0 0 3 6
use FEEDTHRU  F-323
transform 1 0 1797 0 1 928
box 0 0 3 6
use FEEDTHRU  F-324
transform 1 0 1784 0 1 971
box 0 0 3 6
use FEEDTHRU  F-325
transform 1 0 1805 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-326
transform 1 0 1828 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-327
transform 1 0 1858 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-328
transform 1 0 1817 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-329
transform 1 0 1811 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-330
transform 1 0 1827 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-331
transform 1 0 1849 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-332
transform 1 0 1876 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-333
transform 1 0 1838 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-334
transform 1 0 1860 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-335
transform 1 0 1869 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-336
transform 1 0 1848 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-337
transform 1 0 1891 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-338
transform 1 0 1903 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-339
transform 1 0 1874 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-340
transform 1 0 1862 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-341
transform 1 0 1881 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-342
transform 1 0 1828 0 1 971
box 0 0 3 6
use FEEDTHRU  F-343
transform 1 0 1851 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-344
transform 1 0 1885 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-345
transform 1 0 1804 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-346
transform 1 0 1818 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-347
transform 1 0 1796 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-348
transform 1 0 1856 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-349
transform 1 0 1928 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-350
transform 1 0 1937 0 1 1024
box 0 0 3 6
use FEEDTHRU  F-351
transform 1 0 1875 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-352
transform 1 0 1830 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-353
transform 1 0 1859 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-354
transform 1 0 1840 0 1 1698
box 0 0 3 6
use FEEDTHRU  F-355
transform 1 0 1836 0 1 1719
box 0 0 3 6
use FEEDTHRU  F-356
transform 1 0 1869 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-357
transform 1 0 1872 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-358
transform 1 0 1887 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-359
transform 1 0 1809 0 1 1794
box 0 0 3 6
use FEEDTHRU  F-360
transform 1 0 1826 0 1 1775
box 0 0 3 6
use FEEDTHRU  F-361
transform 1 0 1826 0 1 1766
box 0 0 3 6
use FEEDTHRU  F-362
transform 1 0 1826 0 1 1757
box 0 0 3 6
use FEEDTHRU  F-363
transform 1 0 1837 0 1 971
box 0 0 3 6
use FEEDTHRU  F-364
transform 1 0 1856 0 1 928
box 0 0 3 6
use FEEDTHRU  F-365
transform 1 0 1846 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-366
transform 1 0 1846 0 1 971
box 0 0 3 6
use FEEDTHRU  F-367
transform 1 0 1716 0 1 1719
box 0 0 3 6
use FEEDTHRU  F-368
transform 1 0 1710 0 1 1698
box 0 0 3 6
use FEEDTHRU  F-369
transform 1 0 1747 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-370
transform 1 0 1727 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-371
transform 1 0 1763 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-372
transform 1 0 1777 0 1 1476
box 0 0 3 6
use FEEDTHRU  F-373
transform 1 0 1789 0 1 1393
box 0 0 3 6
use FEEDTHRU  F-374
transform 1 0 1766 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-375
transform 1 0 1784 0 1 1267
box 0 0 3 6
use FEEDTHRU  F-376
transform 1 0 1833 0 1 1537
box 0 0 3 6
use FEEDTHRU  F-377
transform 1 0 1931 0 1 1087
box 0 0 3 6
use FEEDTHRU  F-378
transform 1 0 1958 0 1 1168
box 0 0 3 6
use FEEDTHRU  F-379
transform 1 0 1862 0 1 1698
box 0 0 3 6
use FEEDTHRU  F-380
transform 1 0 1896 0 1 1655
box 0 0 3 6
use FEEDTHRU  F-381
transform 1 0 1855 0 1 1610
box 0 0 3 6
use FEEDTHRU  F-382
transform 1 0 1877 0 1 1334
box 0 0 3 6
use FEEDTHRU  F-383
transform 1 0 1893 0 1 1393
box 0 0 3 6
<< metal1 >>
rect 1783 833 1787 834
rect 1813 833 1820 834
rect 1822 833 1829 834
rect 1753 843 1756 844
rect 1783 843 1809 844
rect 1792 845 1818 846
rect 1766 847 1793 848
rect 1813 847 1834 848
rect 1822 849 1843 850
rect 1717 876 1866 877
rect 1919 876 1927 877
rect 1720 885 1893 886
rect 1721 887 1725 888
rect 1755 887 1758 888
rect 1727 889 1755 890
rect 1770 889 1795 890
rect 1792 891 1798 892
rect 1808 891 1814 892
rect 1817 891 1823 892
rect 1842 891 1846 892
rect 1833 893 1843 894
rect 1865 893 1874 894
rect 1876 893 1916 894
rect 1878 895 1896 896
rect 1912 895 1926 896
rect 1922 897 1932 898
rect 1711 906 1725 907
rect 1735 906 1842 907
rect 1745 908 1753 909
rect 1803 908 1821 909
rect 1792 910 1805 911
rect 1822 910 1833 911
rect 1813 912 1824 913
rect 1845 912 1852 913
rect 1873 912 1886 913
rect 1876 914 1889 915
rect 1895 914 1915 915
rect 1912 916 1921 917
rect 1892 918 1912 919
rect 1857 920 1892 921
rect 1925 920 1939 921
rect 1737 922 1939 923
rect 1738 924 1755 925
rect 1727 926 1756 927
rect 1721 935 1726 936
rect 1737 935 1756 936
rect 1753 937 1759 938
rect 1776 937 1796 938
rect 1785 939 1799 940
rect 1795 941 1824 942
rect 1801 943 1821 944
rect 1811 945 1833 946
rect 1817 947 1861 948
rect 1826 949 1842 950
rect 1829 951 1842 952
rect 1838 953 1858 954
rect 1847 955 1895 956
rect 1854 957 1873 958
rect 1866 959 1889 960
rect 1882 961 1945 962
rect 1881 963 1960 964
rect 1885 965 1891 966
rect 1893 965 1939 966
rect 1896 967 1922 968
rect 1908 969 1915 970
rect 1966 969 1974 970
rect 1714 978 1719 979
rect 1729 978 1772 979
rect 1737 980 1750 981
rect 1746 982 1759 983
rect 1753 984 1762 985
rect 1764 984 1804 985
rect 1801 986 1823 987
rect 1826 986 1850 987
rect 1829 988 1853 989
rect 1828 990 1841 991
rect 1838 992 1861 993
rect 1817 994 1838 995
rect 1809 996 1817 997
rect 1861 996 1875 997
rect 1866 998 1885 999
rect 1872 1000 1942 1001
rect 1881 1002 1929 1003
rect 1807 1004 1930 1005
rect 1785 1006 1807 1007
rect 1776 1008 1785 1009
rect 1847 1008 1882 1009
rect 1800 1010 1847 1011
rect 1890 1010 1949 1011
rect 1856 1012 1891 1013
rect 1893 1012 1921 1013
rect 1896 1014 1924 1015
rect 1899 1016 1927 1017
rect 1899 1018 1903 1019
rect 1908 1018 1933 1019
rect 1911 1020 1936 1021
rect 1914 1022 1918 1023
rect 1938 1022 1994 1023
rect 1743 1031 1771 1032
rect 1732 1033 1743 1034
rect 1749 1033 1765 1034
rect 1748 1035 1753 1036
rect 1758 1035 1768 1036
rect 1758 1037 1762 1038
rect 1790 1037 2033 1038
rect 1819 1039 1829 1040
rect 1806 1041 1830 1042
rect 1784 1043 1808 1044
rect 1822 1043 1857 1044
rect 1837 1045 1848 1046
rect 1852 1045 1887 1046
rect 1803 1047 1854 1048
rect 1804 1049 1839 1050
rect 1858 1049 1893 1050
rect 1810 1051 1860 1052
rect 1861 1051 1868 1052
rect 1840 1053 1869 1054
rect 1864 1055 1902 1056
rect 1871 1057 1879 1058
rect 1890 1057 1945 1058
rect 1849 1059 1890 1060
rect 1797 1061 1851 1062
rect 1797 1063 1801 1064
rect 1899 1063 1949 1064
rect 1917 1065 1973 1066
rect 1884 1067 1918 1068
rect 1920 1067 1976 1068
rect 1926 1069 1982 1070
rect 1929 1071 1985 1072
rect 1929 1073 1939 1074
rect 1932 1075 1987 1076
rect 1932 1077 2026 1078
rect 1935 1079 1980 1080
rect 1923 1081 1979 1082
rect 1923 1083 1995 1084
rect 1954 1085 1991 1086
rect 2004 1085 2009 1086
rect 1729 1094 1740 1095
rect 1729 1096 1848 1097
rect 1742 1098 1746 1099
rect 1743 1100 1751 1101
rect 1758 1100 1790 1101
rect 1767 1102 1784 1103
rect 1767 1104 1839 1105
rect 1773 1106 1781 1107
rect 1776 1108 1827 1109
rect 1802 1110 1881 1111
rect 1807 1112 1839 1113
rect 1820 1114 1875 1115
rect 1823 1116 1872 1117
rect 1853 1118 1863 1119
rect 1856 1120 1884 1121
rect 1868 1122 1896 1123
rect 1886 1124 1969 1125
rect 1859 1126 1887 1127
rect 1829 1128 1860 1129
rect 1792 1130 1830 1131
rect 1889 1130 1920 1131
rect 1889 1132 1926 1133
rect 1917 1134 1935 1135
rect 1898 1136 1917 1137
rect 1844 1138 1899 1139
rect 1923 1138 1941 1139
rect 1901 1140 1923 1141
rect 1877 1142 1902 1143
rect 1850 1144 1878 1145
rect 1770 1146 1851 1147
rect 1929 1146 2048 1147
rect 1932 1148 1960 1149
rect 1904 1150 1932 1151
rect 1892 1152 1905 1153
rect 1948 1152 1963 1153
rect 1975 1152 2005 1153
rect 1954 1154 1975 1155
rect 1978 1154 2011 1155
rect 1981 1156 2014 1157
rect 1984 1158 2008 1159
rect 1986 1160 2069 1161
rect 1994 1162 2002 1163
rect 1972 1164 2002 1165
rect 2040 1164 2055 1165
rect 2051 1166 2066 1167
rect 1743 1175 1848 1176
rect 1746 1177 1827 1178
rect 1755 1179 1790 1180
rect 1757 1181 1786 1182
rect 1761 1183 1769 1184
rect 1764 1185 1851 1186
rect 1765 1187 1784 1188
rect 1771 1189 1822 1190
rect 1775 1191 1783 1192
rect 1779 1193 1881 1194
rect 1788 1195 1828 1196
rect 1806 1197 1825 1198
rect 1806 1199 1830 1200
rect 1812 1201 1863 1202
rect 1816 1203 1884 1204
rect 1818 1205 1860 1206
rect 1830 1207 1858 1208
rect 1838 1209 2062 1210
rect 1839 1211 1878 1212
rect 1841 1213 1890 1214
rect 1842 1215 1945 1216
rect 1844 1217 1902 1218
rect 1845 1219 1887 1220
rect 1860 1221 1875 1222
rect 1866 1223 1896 1224
rect 1875 1225 1905 1226
rect 1887 1227 1982 1228
rect 1893 1229 1917 1230
rect 1896 1231 1920 1232
rect 1911 1233 1932 1234
rect 1914 1235 1947 1236
rect 1917 1237 1935 1238
rect 1922 1239 1954 1240
rect 1923 1241 1941 1242
rect 1928 1243 1933 1244
rect 1935 1243 2020 1244
rect 1959 1245 1979 1246
rect 1960 1247 2059 1248
rect 1962 1249 2017 1250
rect 1863 1251 2018 1252
rect 1963 1253 2069 1254
rect 1972 1255 2005 1256
rect 1986 1257 2045 1258
rect 1991 1259 2008 1260
rect 1995 1261 2002 1262
rect 1994 1263 2011 1264
rect 1997 1265 2014 1266
rect 1717 1274 1725 1275
rect 1748 1274 1753 1275
rect 1755 1274 1759 1275
rect 1761 1274 1798 1275
rect 1768 1276 1822 1277
rect 1767 1278 1786 1279
rect 1782 1280 1825 1281
rect 1788 1282 1843 1283
rect 1791 1284 1831 1285
rect 1812 1286 1834 1287
rect 1812 1288 1819 1289
rect 1815 1290 1982 1291
rect 1836 1292 1861 1293
rect 1839 1294 1873 1295
rect 1842 1296 1864 1297
rect 1845 1298 1867 1299
rect 1857 1300 1949 1301
rect 1860 1302 1897 1303
rect 1863 1304 1876 1305
rect 1878 1304 1979 1305
rect 1881 1306 1912 1307
rect 1884 1308 1888 1309
rect 1893 1308 2011 1309
rect 1900 1310 1918 1311
rect 1914 1312 1930 1313
rect 1923 1314 1934 1315
rect 1924 1316 1976 1317
rect 1927 1318 1936 1319
rect 1930 1320 1998 1321
rect 1946 1322 1973 1323
rect 1951 1324 1964 1325
rect 1950 1326 1980 1327
rect 1956 1328 1992 1329
rect 1960 1330 2036 1331
rect 1982 1332 1995 1333
rect 1741 1341 1765 1342
rect 1748 1343 1762 1344
rect 1752 1345 1785 1346
rect 1767 1347 1791 1348
rect 1758 1349 1768 1350
rect 1773 1349 1998 1350
rect 1793 1351 1841 1352
rect 1797 1353 1820 1354
rect 1812 1355 1829 1356
rect 1824 1357 1882 1358
rect 1830 1359 1844 1360
rect 1815 1361 1832 1362
rect 1833 1361 1853 1362
rect 1836 1363 1856 1364
rect 1849 1365 1888 1366
rect 1863 1367 1883 1368
rect 1845 1369 1865 1370
rect 1875 1369 1936 1370
rect 1878 1371 1895 1372
rect 1860 1373 1880 1374
rect 1888 1373 1940 1374
rect 1915 1375 1939 1376
rect 1914 1377 1951 1378
rect 1924 1379 1966 1380
rect 1900 1381 1924 1382
rect 1927 1381 1969 1382
rect 1930 1383 1954 1384
rect 1943 1385 2019 1386
rect 1956 1387 2001 1388
rect 1933 1389 1957 1390
rect 1979 1389 2022 1390
rect 2009 1391 2042 1392
rect 1729 1400 1737 1401
rect 1740 1400 1762 1401
rect 1744 1402 1794 1403
rect 1751 1404 1844 1405
rect 1755 1406 1809 1407
rect 1761 1408 1829 1409
rect 1764 1410 1781 1411
rect 1767 1412 1838 1413
rect 1768 1414 1832 1415
rect 1778 1416 1791 1417
rect 1800 1416 1850 1417
rect 1805 1418 1820 1419
rect 1831 1418 1853 1419
rect 1834 1420 1841 1421
rect 1840 1422 1859 1423
rect 1843 1424 1856 1425
rect 1852 1426 1865 1427
rect 1855 1428 1868 1429
rect 1861 1430 1880 1431
rect 1867 1432 1886 1433
rect 1870 1434 1887 1435
rect 1873 1436 1889 1437
rect 1882 1438 1963 1439
rect 1821 1440 1883 1441
rect 1894 1440 1972 1441
rect 1898 1442 1936 1443
rect 1901 1444 1939 1445
rect 1904 1446 1924 1447
rect 1907 1448 1948 1449
rect 1928 1450 1954 1451
rect 1931 1452 1957 1453
rect 1934 1454 1950 1455
rect 1937 1456 1966 1457
rect 1940 1458 1969 1459
rect 1943 1460 2025 1461
rect 1972 1462 1998 1463
rect 1975 1464 2001 1465
rect 1978 1466 2042 1467
rect 1987 1468 2039 1469
rect 2018 1470 2035 1471
rect 2005 1472 2036 1473
rect 2021 1474 2032 1475
rect 1696 1483 1871 1484
rect 1723 1485 1734 1486
rect 1730 1487 1738 1488
rect 1723 1489 1731 1490
rect 1744 1489 1809 1490
rect 1744 1491 1794 1492
rect 1747 1493 1806 1494
rect 1751 1495 1789 1496
rect 1765 1497 1805 1498
rect 1764 1499 1779 1500
rect 1791 1499 1832 1500
rect 1799 1501 1802 1502
rect 1811 1501 1954 1502
rect 1813 1503 1826 1504
rect 1816 1505 1835 1506
rect 1819 1507 1850 1508
rect 1825 1509 1844 1510
rect 1831 1511 1835 1512
rect 1846 1511 1853 1512
rect 1855 1511 1862 1512
rect 1867 1511 1883 1512
rect 1870 1513 1874 1514
rect 1876 1513 1923 1514
rect 1894 1515 1905 1516
rect 1898 1517 1913 1518
rect 1901 1519 1916 1520
rect 1900 1521 1932 1522
rect 1928 1523 1949 1524
rect 1934 1525 1962 1526
rect 1945 1527 1964 1528
rect 1975 1527 1990 1528
rect 1987 1529 2002 1530
rect 1972 1531 1987 1532
rect 1998 1531 2009 1532
rect 2005 1533 2029 1534
rect 2021 1535 2026 1536
rect 2028 1535 2033 1536
rect 1693 1544 1862 1545
rect 1706 1546 1720 1547
rect 1728 1546 1765 1547
rect 1730 1548 1738 1549
rect 1738 1550 1749 1551
rect 1745 1552 1760 1553
rect 1779 1552 1805 1553
rect 1791 1554 1802 1555
rect 1795 1556 1814 1557
rect 1810 1558 1826 1559
rect 1813 1560 1823 1561
rect 1816 1562 1838 1563
rect 1816 1564 1850 1565
rect 1822 1566 1835 1567
rect 1825 1568 1859 1569
rect 1828 1570 1865 1571
rect 1831 1572 1877 1573
rect 1844 1574 1946 1575
rect 1846 1576 1973 1577
rect 1856 1578 1966 1579
rect 1870 1580 1934 1581
rect 1871 1582 1913 1583
rect 1874 1584 1916 1585
rect 1883 1586 1949 1587
rect 1886 1588 1901 1589
rect 1894 1590 1922 1591
rect 1895 1592 1980 1593
rect 1898 1594 1940 1595
rect 1901 1596 1943 1597
rect 1931 1598 1978 1599
rect 1934 1600 1987 1601
rect 1936 1602 2019 1603
rect 1949 1604 1999 1605
rect 1952 1606 2002 1607
rect 1989 1608 2008 1609
rect 1699 1617 1707 1618
rect 1713 1617 1720 1618
rect 1725 1617 1739 1618
rect 1728 1619 1749 1620
rect 1752 1619 1783 1620
rect 1722 1621 1752 1622
rect 1755 1621 1765 1622
rect 1762 1623 1770 1624
rect 1779 1623 1795 1624
rect 1785 1625 1829 1626
rect 1791 1627 1810 1628
rect 1801 1629 1817 1630
rect 1776 1631 1801 1632
rect 1775 1633 1798 1634
rect 1813 1633 1820 1634
rect 1825 1633 1912 1634
rect 1831 1635 1861 1636
rect 1871 1635 1908 1636
rect 1874 1637 1881 1638
rect 1883 1637 1913 1638
rect 1886 1639 1889 1640
rect 1895 1639 1915 1640
rect 1894 1641 1945 1642
rect 1901 1643 1904 1644
rect 1898 1645 1901 1646
rect 1856 1647 1898 1648
rect 1915 1647 1929 1648
rect 1928 1649 1950 1650
rect 1931 1651 1958 1652
rect 1934 1653 1939 1654
rect 1952 1653 1955 1654
rect 1711 1662 1749 1663
rect 1723 1664 1752 1665
rect 1757 1664 1765 1665
rect 1759 1666 1762 1667
rect 1763 1666 1798 1667
rect 1766 1668 1810 1669
rect 1778 1670 1801 1671
rect 1794 1672 1816 1673
rect 1801 1674 1958 1675
rect 1804 1676 1823 1677
rect 1826 1676 1834 1677
rect 1841 1676 1861 1677
rect 1857 1678 1904 1679
rect 1863 1680 1898 1681
rect 1878 1682 1916 1683
rect 1881 1684 1889 1685
rect 1884 1686 1919 1687
rect 1887 1688 1901 1689
rect 1894 1690 1936 1691
rect 1910 1692 1939 1693
rect 1912 1694 1949 1695
rect 1941 1696 1955 1697
rect 1969 1696 1977 1697
rect 1711 1705 1718 1706
rect 1720 1705 1724 1706
rect 1759 1705 1764 1706
rect 1834 1705 1848 1706
rect 1837 1707 1842 1708
rect 1857 1707 1914 1708
rect 1863 1709 1905 1710
rect 1872 1711 1885 1712
rect 1875 1713 1888 1714
rect 1878 1715 1908 1716
rect 1878 1717 1901 1718
rect 1904 1717 1911 1718
rect 1916 1717 1938 1718
rect 1711 1726 1718 1727
rect 1720 1726 1750 1727
rect 1770 1726 1785 1727
rect 1804 1726 1832 1727
rect 1780 1728 1805 1729
rect 1780 1730 1792 1731
rect 1831 1730 1882 1731
rect 1834 1732 1844 1733
rect 1834 1734 1841 1735
rect 1837 1736 1908 1737
rect 1847 1738 1858 1739
rect 1863 1738 1873 1739
rect 1866 1740 1876 1741
rect 1869 1742 1879 1743
rect 1892 1742 1905 1743
rect 1681 1751 1689 1752
rect 1780 1751 1785 1752
rect 1801 1751 1805 1752
rect 1827 1751 1832 1752
rect 1834 1751 1837 1752
rect 1869 1751 1872 1752
rect 1866 1753 1869 1754
rect 1863 1755 1866 1756
rect 1892 1755 1899 1756
rect 1714 1782 1869 1783
rect 1801 1784 1812 1785
rect 1810 1786 1828 1787
rect 1819 1788 1837 1789
rect 1837 1790 1866 1791
rect 1840 1792 1872 1793
rect 1714 1801 1719 1802
rect 1762 1801 1841 1802
rect 1774 1803 1802 1804
rect 1795 1805 1838 1806
rect 1810 1807 1814 1808
rect 1819 1807 1823 1808
<< metal2 >>
rect 1783 833 1784 837
rect 1786 833 1787 837
rect 1813 833 1814 837
rect 1819 833 1820 837
rect 1822 833 1823 837
rect 1828 833 1829 837
rect 1753 841 1754 844
rect 1755 843 1756 852
rect 1783 841 1784 844
rect 1808 843 1809 852
rect 1792 841 1793 846
rect 1817 845 1818 852
rect 1766 841 1767 848
rect 1792 847 1793 852
rect 1813 841 1814 848
rect 1833 847 1834 852
rect 1822 841 1823 850
rect 1842 849 1843 852
rect 1755 858 1756 861
rect 1755 856 1756 859
rect 1792 858 1793 861
rect 1792 856 1793 859
rect 1808 858 1809 861
rect 1808 856 1809 859
rect 1817 858 1818 861
rect 1817 856 1818 859
rect 1833 858 1834 861
rect 1833 856 1834 859
rect 1842 858 1843 861
rect 1842 856 1843 859
rect 1755 867 1756 870
rect 1755 865 1756 868
rect 1792 867 1793 870
rect 1792 865 1793 868
rect 1808 867 1809 870
rect 1808 865 1809 868
rect 1817 867 1818 870
rect 1817 865 1818 868
rect 1833 867 1834 870
rect 1833 865 1834 868
rect 1842 867 1843 870
rect 1842 865 1843 868
rect 1717 876 1718 879
rect 1865 876 1866 879
rect 1755 876 1756 879
rect 1755 874 1756 877
rect 1792 876 1793 879
rect 1792 874 1793 877
rect 1808 876 1809 879
rect 1808 874 1809 877
rect 1817 876 1818 879
rect 1817 874 1818 877
rect 1833 876 1834 879
rect 1833 874 1834 877
rect 1842 876 1843 879
rect 1842 874 1843 877
rect 1919 876 1920 879
rect 1926 876 1927 879
rect 1720 883 1721 886
rect 1892 885 1893 900
rect 1721 887 1722 900
rect 1724 887 1725 900
rect 1755 883 1756 888
rect 1757 887 1758 900
rect 1727 889 1728 900
rect 1754 889 1755 900
rect 1770 889 1771 900
rect 1794 889 1795 900
rect 1792 883 1793 892
rect 1797 891 1798 900
rect 1808 883 1809 892
rect 1813 891 1814 900
rect 1817 883 1818 892
rect 1822 891 1823 900
rect 1842 883 1843 892
rect 1845 891 1846 900
rect 1833 883 1834 894
rect 1842 893 1843 900
rect 1865 883 1866 894
rect 1873 893 1874 900
rect 1876 893 1877 900
rect 1915 893 1916 900
rect 1878 883 1879 896
rect 1895 895 1896 900
rect 1912 883 1913 896
rect 1925 895 1926 900
rect 1922 897 1923 900
rect 1931 897 1932 900
rect 1711 904 1712 907
rect 1724 904 1725 907
rect 1735 906 1736 929
rect 1841 906 1842 929
rect 1745 908 1746 929
rect 1752 908 1753 929
rect 1757 904 1758 909
rect 1758 908 1759 929
rect 1803 904 1804 909
rect 1820 908 1821 929
rect 1792 910 1793 929
rect 1804 910 1805 929
rect 1822 904 1823 911
rect 1832 910 1833 929
rect 1813 904 1814 913
rect 1823 912 1824 929
rect 1845 904 1846 913
rect 1851 904 1852 913
rect 1873 904 1874 913
rect 1885 912 1886 929
rect 1876 904 1877 915
rect 1888 914 1889 929
rect 1895 904 1896 915
rect 1914 914 1915 929
rect 1912 904 1913 917
rect 1920 916 1921 929
rect 1892 904 1893 919
rect 1911 918 1912 929
rect 1857 920 1858 929
rect 1891 920 1892 929
rect 1925 904 1926 921
rect 1938 904 1939 921
rect 1737 904 1738 923
rect 1938 922 1939 929
rect 1738 924 1739 929
rect 1754 904 1755 925
rect 1727 904 1728 927
rect 1755 926 1756 929
rect 1944 926 1945 929
rect 1945 904 1946 927
rect 1721 935 1722 972
rect 1725 935 1726 972
rect 1737 935 1738 972
rect 1755 933 1756 936
rect 1753 937 1754 972
rect 1758 933 1759 938
rect 1776 937 1777 972
rect 1795 933 1796 938
rect 1785 939 1786 972
rect 1798 933 1799 940
rect 1795 941 1796 972
rect 1823 933 1824 942
rect 1801 943 1802 972
rect 1820 933 1821 944
rect 1811 945 1812 972
rect 1832 933 1833 946
rect 1817 947 1818 972
rect 1860 933 1861 948
rect 1826 949 1827 972
rect 1841 933 1842 950
rect 1829 951 1830 972
rect 1841 951 1842 972
rect 1838 953 1839 972
rect 1857 933 1858 954
rect 1847 955 1848 972
rect 1894 933 1895 956
rect 1854 933 1855 958
rect 1872 957 1873 972
rect 1866 959 1867 972
rect 1888 933 1889 960
rect 1882 933 1883 962
rect 1944 933 1945 962
rect 1881 963 1882 972
rect 1959 963 1960 972
rect 1885 933 1886 966
rect 1890 965 1891 972
rect 1893 965 1894 972
rect 1938 933 1939 966
rect 1896 967 1897 972
rect 1921 967 1922 972
rect 1898 933 1899 970
rect 1899 969 1900 972
rect 1908 969 1909 972
rect 1914 933 1915 970
rect 1911 969 1912 972
rect 1911 933 1912 970
rect 1966 969 1967 972
rect 1973 969 1974 972
rect 1714 976 1715 979
rect 1718 976 1719 979
rect 1729 978 1730 1025
rect 1771 978 1772 1025
rect 1737 976 1738 981
rect 1749 980 1750 1025
rect 1746 982 1747 1025
rect 1758 982 1759 1025
rect 1753 976 1754 985
rect 1761 984 1762 1025
rect 1764 984 1765 1025
rect 1803 984 1804 1025
rect 1801 976 1802 987
rect 1822 986 1823 1025
rect 1826 976 1827 987
rect 1849 986 1850 1025
rect 1829 976 1830 989
rect 1852 988 1853 1025
rect 1828 990 1829 1025
rect 1840 990 1841 1025
rect 1838 976 1839 993
rect 1860 976 1861 993
rect 1817 976 1818 995
rect 1837 994 1838 1025
rect 1809 996 1810 1025
rect 1816 996 1817 1025
rect 1861 996 1862 1025
rect 1874 996 1875 1025
rect 1866 976 1867 999
rect 1884 998 1885 1025
rect 1872 976 1873 1001
rect 1941 1000 1942 1025
rect 1881 976 1882 1003
rect 1928 976 1929 1003
rect 1807 976 1808 1005
rect 1929 1004 1930 1025
rect 1785 976 1786 1007
rect 1806 1006 1807 1025
rect 1776 976 1777 1009
rect 1784 1008 1785 1025
rect 1847 976 1848 1009
rect 1881 1008 1882 1025
rect 1800 1010 1801 1025
rect 1846 1010 1847 1025
rect 1890 976 1891 1011
rect 1948 1010 1949 1025
rect 1856 976 1857 1013
rect 1890 1012 1891 1025
rect 1893 976 1894 1013
rect 1920 1012 1921 1025
rect 1896 976 1897 1015
rect 1923 1014 1924 1025
rect 1899 976 1900 1017
rect 1926 1016 1927 1025
rect 1899 1018 1900 1025
rect 1902 976 1903 1019
rect 1908 976 1909 1019
rect 1932 1018 1933 1025
rect 1911 976 1912 1021
rect 1935 1020 1936 1025
rect 1914 976 1915 1023
rect 1917 1022 1918 1025
rect 1938 1022 1939 1025
rect 1993 1022 1994 1025
rect 1743 1029 1744 1032
rect 1770 1031 1771 1088
rect 1732 1033 1733 1088
rect 1742 1033 1743 1088
rect 1749 1029 1750 1034
rect 1764 1029 1765 1034
rect 1748 1035 1749 1088
rect 1752 1035 1753 1088
rect 1758 1029 1759 1036
rect 1767 1035 1768 1088
rect 1758 1037 1759 1088
rect 1761 1029 1762 1038
rect 1790 1037 1791 1088
rect 2032 1037 2033 1088
rect 1819 1029 1820 1040
rect 1828 1029 1829 1040
rect 1806 1029 1807 1042
rect 1829 1041 1830 1088
rect 1784 1029 1785 1044
rect 1807 1043 1808 1088
rect 1822 1029 1823 1044
rect 1856 1043 1857 1088
rect 1837 1029 1838 1046
rect 1847 1045 1848 1088
rect 1852 1029 1853 1046
rect 1886 1045 1887 1088
rect 1803 1029 1804 1048
rect 1853 1047 1854 1088
rect 1804 1049 1805 1088
rect 1838 1049 1839 1088
rect 1858 1029 1859 1050
rect 1892 1049 1893 1088
rect 1810 1051 1811 1088
rect 1859 1051 1860 1088
rect 1861 1029 1862 1052
rect 1867 1029 1868 1052
rect 1840 1029 1841 1054
rect 1868 1053 1869 1088
rect 1864 1029 1865 1056
rect 1901 1055 1902 1088
rect 1871 1057 1872 1088
rect 1878 1029 1879 1058
rect 1890 1029 1891 1058
rect 1944 1029 1945 1058
rect 1849 1029 1850 1060
rect 1889 1059 1890 1088
rect 1797 1029 1798 1062
rect 1850 1061 1851 1088
rect 1797 1063 1798 1088
rect 1800 1029 1801 1064
rect 1899 1029 1900 1064
rect 1948 1063 1949 1088
rect 1917 1029 1918 1066
rect 1972 1065 1973 1088
rect 1884 1029 1885 1068
rect 1917 1067 1918 1088
rect 1920 1029 1921 1068
rect 1975 1067 1976 1088
rect 1926 1029 1927 1070
rect 1981 1069 1982 1088
rect 1929 1029 1930 1072
rect 1984 1071 1985 1088
rect 1929 1073 1930 1088
rect 1938 1029 1939 1074
rect 1932 1029 1933 1076
rect 1986 1029 1987 1076
rect 1932 1077 1933 1088
rect 2025 1077 2026 1088
rect 1935 1029 1936 1080
rect 1979 1029 1980 1080
rect 1923 1029 1924 1082
rect 1978 1081 1979 1088
rect 1923 1083 1924 1088
rect 1994 1083 1995 1088
rect 1954 1085 1955 1088
rect 1990 1085 1991 1088
rect 2004 1085 2005 1088
rect 2008 1085 2009 1088
rect 1729 1092 1730 1095
rect 1739 1092 1740 1095
rect 1729 1096 1730 1169
rect 1847 1096 1848 1169
rect 1742 1092 1743 1099
rect 1745 1092 1746 1099
rect 1743 1100 1744 1169
rect 1750 1100 1751 1169
rect 1758 1092 1759 1101
rect 1789 1100 1790 1169
rect 1767 1092 1768 1103
rect 1783 1102 1784 1169
rect 1767 1104 1768 1169
rect 1838 1092 1839 1105
rect 1773 1092 1774 1107
rect 1780 1092 1781 1107
rect 1776 1092 1777 1109
rect 1826 1108 1827 1169
rect 1802 1110 1803 1169
rect 1880 1110 1881 1169
rect 1807 1092 1808 1113
rect 1838 1112 1839 1169
rect 1820 1092 1821 1115
rect 1874 1114 1875 1169
rect 1823 1116 1824 1169
rect 1871 1092 1872 1117
rect 1853 1092 1854 1119
rect 1862 1118 1863 1169
rect 1856 1092 1857 1121
rect 1883 1120 1884 1169
rect 1868 1092 1869 1123
rect 1895 1122 1896 1169
rect 1886 1092 1887 1125
rect 1968 1124 1969 1169
rect 1859 1092 1860 1127
rect 1886 1126 1887 1169
rect 1829 1092 1830 1129
rect 1859 1128 1860 1169
rect 1792 1130 1793 1169
rect 1829 1130 1830 1169
rect 1889 1092 1890 1131
rect 1919 1130 1920 1169
rect 1889 1132 1890 1169
rect 1925 1132 1926 1169
rect 1917 1092 1918 1135
rect 1934 1134 1935 1169
rect 1898 1092 1899 1137
rect 1916 1136 1917 1169
rect 1844 1138 1845 1169
rect 1898 1138 1899 1169
rect 1923 1092 1924 1139
rect 1940 1138 1941 1169
rect 1901 1092 1902 1141
rect 1922 1140 1923 1169
rect 1877 1092 1878 1143
rect 1901 1142 1902 1169
rect 1850 1092 1851 1145
rect 1877 1144 1878 1169
rect 1770 1092 1771 1147
rect 1850 1146 1851 1169
rect 1929 1092 1930 1147
rect 2047 1146 2048 1169
rect 1932 1092 1933 1149
rect 1959 1148 1960 1169
rect 1904 1092 1905 1151
rect 1931 1150 1932 1169
rect 1892 1092 1893 1153
rect 1904 1152 1905 1169
rect 1948 1092 1949 1153
rect 1962 1152 1963 1169
rect 1975 1092 1976 1153
rect 2004 1152 2005 1169
rect 1954 1092 1955 1155
rect 1974 1154 1975 1169
rect 1978 1092 1979 1155
rect 2010 1154 2011 1169
rect 1981 1092 1982 1157
rect 2013 1156 2014 1169
rect 1984 1092 1985 1159
rect 2007 1158 2008 1169
rect 1986 1160 1987 1169
rect 2068 1160 2069 1169
rect 1994 1092 1995 1163
rect 2001 1092 2002 1163
rect 1972 1092 1973 1165
rect 2001 1164 2002 1169
rect 2040 1164 2041 1169
rect 2054 1164 2055 1169
rect 2051 1166 2052 1169
rect 2065 1166 2066 1169
rect 1743 1173 1744 1176
rect 1847 1173 1848 1176
rect 1746 1173 1747 1178
rect 1826 1173 1827 1178
rect 1755 1179 1756 1268
rect 1789 1173 1790 1180
rect 1757 1173 1758 1182
rect 1785 1181 1786 1268
rect 1761 1183 1762 1268
rect 1768 1183 1769 1268
rect 1764 1173 1765 1186
rect 1850 1173 1851 1186
rect 1765 1187 1766 1268
rect 1783 1173 1784 1188
rect 1771 1173 1772 1190
rect 1821 1189 1822 1268
rect 1775 1191 1776 1268
rect 1782 1191 1783 1268
rect 1779 1193 1780 1268
rect 1880 1173 1881 1194
rect 1788 1195 1789 1268
rect 1827 1195 1828 1268
rect 1806 1173 1807 1198
rect 1824 1197 1825 1268
rect 1806 1199 1807 1268
rect 1829 1173 1830 1200
rect 1812 1201 1813 1268
rect 1862 1173 1863 1202
rect 1816 1173 1817 1204
rect 1883 1173 1884 1204
rect 1818 1205 1819 1268
rect 1859 1173 1860 1206
rect 1830 1207 1831 1268
rect 1857 1207 1858 1268
rect 1838 1173 1839 1210
rect 2061 1173 2062 1210
rect 1839 1211 1840 1268
rect 1877 1173 1878 1212
rect 1841 1173 1842 1214
rect 1889 1173 1890 1214
rect 1842 1215 1843 1268
rect 1944 1215 1945 1268
rect 1844 1173 1845 1218
rect 1901 1173 1902 1218
rect 1845 1219 1846 1268
rect 1886 1173 1887 1220
rect 1860 1221 1861 1268
rect 1874 1173 1875 1222
rect 1866 1223 1867 1268
rect 1895 1173 1896 1224
rect 1875 1225 1876 1268
rect 1904 1173 1905 1226
rect 1887 1227 1888 1268
rect 1981 1227 1982 1268
rect 1893 1229 1894 1268
rect 1916 1173 1917 1230
rect 1896 1231 1897 1268
rect 1919 1173 1920 1232
rect 1898 1173 1899 1234
rect 1899 1233 1900 1268
rect 1911 1233 1912 1268
rect 1931 1173 1932 1234
rect 1914 1235 1915 1268
rect 1946 1173 1947 1236
rect 1917 1237 1918 1268
rect 1934 1173 1935 1238
rect 1922 1173 1923 1240
rect 1953 1173 1954 1240
rect 1923 1241 1924 1268
rect 1940 1173 1941 1242
rect 1928 1173 1929 1244
rect 1932 1243 1933 1268
rect 1935 1243 1936 1268
rect 2019 1173 2020 1244
rect 1959 1173 1960 1246
rect 1978 1245 1979 1268
rect 1960 1247 1961 1268
rect 2058 1173 2059 1248
rect 1962 1173 1963 1250
rect 2016 1173 2017 1250
rect 1863 1251 1864 1268
rect 2017 1251 2018 1268
rect 1963 1253 1964 1268
rect 2068 1173 2069 1254
rect 1972 1255 1973 1268
rect 2004 1173 2005 1256
rect 1974 1173 1975 1258
rect 1975 1257 1976 1268
rect 1986 1173 1987 1258
rect 2044 1173 2045 1258
rect 1991 1259 1992 1268
rect 2007 1173 2008 1260
rect 1995 1173 1996 1262
rect 2001 1173 2002 1262
rect 1994 1263 1995 1268
rect 2010 1173 2011 1264
rect 1997 1265 1998 1268
rect 2013 1173 2014 1266
rect 1717 1274 1718 1335
rect 1724 1274 1725 1335
rect 1748 1274 1749 1335
rect 1752 1272 1753 1275
rect 1755 1272 1756 1275
rect 1758 1274 1759 1335
rect 1761 1272 1762 1275
rect 1797 1274 1798 1335
rect 1768 1272 1769 1277
rect 1821 1272 1822 1277
rect 1767 1278 1768 1335
rect 1785 1272 1786 1279
rect 1782 1272 1783 1281
rect 1824 1272 1825 1281
rect 1788 1272 1789 1283
rect 1842 1272 1843 1283
rect 1791 1284 1792 1335
rect 1830 1284 1831 1335
rect 1812 1272 1813 1287
rect 1833 1286 1834 1335
rect 1812 1288 1813 1335
rect 1818 1272 1819 1289
rect 1815 1290 1816 1335
rect 1981 1272 1982 1291
rect 1836 1292 1837 1335
rect 1860 1272 1861 1293
rect 1839 1272 1840 1295
rect 1872 1272 1873 1295
rect 1842 1296 1843 1335
rect 1863 1272 1864 1297
rect 1845 1298 1846 1335
rect 1866 1272 1867 1299
rect 1857 1272 1858 1301
rect 1948 1272 1949 1301
rect 1860 1302 1861 1335
rect 1896 1272 1897 1303
rect 1863 1304 1864 1335
rect 1875 1272 1876 1305
rect 1878 1304 1879 1335
rect 1978 1272 1979 1305
rect 1881 1306 1882 1335
rect 1911 1272 1912 1307
rect 1884 1308 1885 1335
rect 1887 1272 1888 1309
rect 1893 1272 1894 1309
rect 2010 1272 2011 1309
rect 1900 1310 1901 1335
rect 1917 1272 1918 1311
rect 1914 1272 1915 1313
rect 1929 1272 1930 1313
rect 1923 1272 1924 1315
rect 1933 1314 1934 1335
rect 1924 1316 1925 1335
rect 1975 1272 1976 1317
rect 1927 1318 1928 1335
rect 1935 1272 1936 1319
rect 1930 1320 1931 1335
rect 1997 1272 1998 1321
rect 1946 1322 1947 1335
rect 1972 1272 1973 1323
rect 1951 1272 1952 1325
rect 1963 1272 1964 1325
rect 1950 1326 1951 1335
rect 1979 1326 1980 1335
rect 1956 1328 1957 1335
rect 1991 1272 1992 1329
rect 1960 1272 1961 1331
rect 2035 1272 2036 1331
rect 1982 1332 1983 1335
rect 1994 1272 1995 1333
rect 1741 1339 1742 1342
rect 1764 1341 1765 1394
rect 1748 1343 1749 1394
rect 1761 1343 1762 1394
rect 1752 1339 1753 1346
rect 1784 1339 1785 1346
rect 1767 1339 1768 1348
rect 1790 1347 1791 1394
rect 1758 1339 1759 1350
rect 1767 1349 1768 1394
rect 1773 1339 1774 1350
rect 1997 1349 1998 1394
rect 1793 1351 1794 1394
rect 1840 1351 1841 1394
rect 1797 1339 1798 1354
rect 1819 1353 1820 1394
rect 1812 1339 1813 1356
rect 1828 1355 1829 1394
rect 1824 1339 1825 1358
rect 1881 1339 1882 1358
rect 1830 1339 1831 1360
rect 1843 1359 1844 1394
rect 1815 1339 1816 1362
rect 1831 1361 1832 1394
rect 1833 1339 1834 1362
rect 1852 1361 1853 1394
rect 1836 1339 1837 1364
rect 1855 1363 1856 1394
rect 1849 1365 1850 1394
rect 1887 1339 1888 1366
rect 1863 1339 1864 1368
rect 1882 1367 1883 1394
rect 1845 1339 1846 1370
rect 1864 1369 1865 1394
rect 1875 1339 1876 1370
rect 1935 1369 1936 1394
rect 1878 1339 1879 1372
rect 1894 1371 1895 1394
rect 1860 1339 1861 1374
rect 1879 1373 1880 1394
rect 1884 1339 1885 1374
rect 1885 1373 1886 1394
rect 1888 1373 1889 1394
rect 1939 1339 1940 1374
rect 1915 1339 1916 1376
rect 1938 1375 1939 1394
rect 1914 1377 1915 1394
rect 1950 1377 1951 1394
rect 1924 1339 1925 1380
rect 1965 1379 1966 1394
rect 1900 1339 1901 1382
rect 1923 1381 1924 1394
rect 1927 1339 1928 1382
rect 1968 1381 1969 1394
rect 1930 1339 1931 1384
rect 1953 1383 1954 1394
rect 1943 1339 1944 1386
rect 2018 1385 2019 1394
rect 1956 1339 1957 1388
rect 2000 1387 2001 1394
rect 1933 1339 1934 1390
rect 1956 1389 1957 1394
rect 1979 1339 1980 1390
rect 2021 1389 2022 1394
rect 2009 1391 2010 1394
rect 2041 1391 2042 1394
rect 1729 1398 1730 1401
rect 1736 1398 1737 1401
rect 1740 1400 1741 1477
rect 1761 1398 1762 1401
rect 1744 1402 1745 1477
rect 1793 1402 1794 1477
rect 1751 1404 1752 1477
rect 1843 1398 1844 1405
rect 1755 1398 1756 1407
rect 1808 1406 1809 1477
rect 1761 1408 1762 1477
rect 1828 1398 1829 1409
rect 1764 1398 1765 1411
rect 1780 1398 1781 1411
rect 1767 1398 1768 1413
rect 1837 1398 1838 1413
rect 1768 1414 1769 1477
rect 1831 1398 1832 1415
rect 1778 1416 1779 1477
rect 1790 1398 1791 1417
rect 1800 1398 1801 1417
rect 1849 1398 1850 1417
rect 1805 1418 1806 1477
rect 1819 1398 1820 1419
rect 1831 1418 1832 1477
rect 1852 1398 1853 1419
rect 1834 1420 1835 1477
rect 1840 1398 1841 1421
rect 1840 1422 1841 1477
rect 1858 1422 1859 1477
rect 1843 1424 1844 1477
rect 1855 1398 1856 1425
rect 1852 1426 1853 1477
rect 1864 1398 1865 1427
rect 1855 1428 1856 1477
rect 1867 1398 1868 1429
rect 1861 1430 1862 1477
rect 1879 1398 1880 1431
rect 1867 1432 1868 1477
rect 1885 1398 1886 1433
rect 1870 1434 1871 1477
rect 1886 1434 1887 1477
rect 1873 1436 1874 1477
rect 1888 1398 1889 1437
rect 1882 1398 1883 1439
rect 1962 1398 1963 1439
rect 1821 1440 1822 1477
rect 1882 1440 1883 1477
rect 1894 1398 1895 1441
rect 1971 1398 1972 1441
rect 1898 1442 1899 1477
rect 1935 1398 1936 1443
rect 1901 1444 1902 1477
rect 1938 1398 1939 1445
rect 1904 1446 1905 1477
rect 1923 1398 1924 1447
rect 1907 1398 1908 1449
rect 1947 1398 1948 1449
rect 1928 1450 1929 1477
rect 1953 1398 1954 1451
rect 1931 1452 1932 1477
rect 1956 1398 1957 1453
rect 1934 1454 1935 1477
rect 1949 1454 1950 1477
rect 1937 1456 1938 1477
rect 1965 1398 1966 1457
rect 1940 1458 1941 1477
rect 1968 1398 1969 1459
rect 1943 1460 1944 1477
rect 2024 1398 2025 1461
rect 1972 1462 1973 1477
rect 1997 1398 1998 1463
rect 1975 1464 1976 1477
rect 2000 1398 2001 1465
rect 1978 1466 1979 1477
rect 2041 1466 2042 1477
rect 1987 1468 1988 1477
rect 2038 1398 2039 1469
rect 2008 1470 2009 1477
rect 2009 1398 2010 1471
rect 2018 1398 2019 1471
rect 2034 1398 2035 1471
rect 2005 1472 2006 1477
rect 2035 1472 2036 1477
rect 2021 1398 2022 1475
rect 2031 1398 2032 1475
rect 1696 1483 1697 1538
rect 1870 1481 1871 1484
rect 1723 1481 1724 1486
rect 1733 1481 1734 1486
rect 1730 1481 1731 1488
rect 1737 1481 1738 1488
rect 1723 1489 1724 1538
rect 1730 1489 1731 1538
rect 1744 1481 1745 1490
rect 1808 1481 1809 1490
rect 1744 1491 1745 1538
rect 1793 1481 1794 1492
rect 1747 1493 1748 1538
rect 1805 1481 1806 1494
rect 1751 1495 1752 1538
rect 1788 1495 1789 1538
rect 1765 1481 1766 1498
rect 1804 1497 1805 1538
rect 1764 1499 1765 1538
rect 1778 1481 1779 1500
rect 1791 1499 1792 1538
rect 1831 1481 1832 1500
rect 1799 1481 1800 1502
rect 1801 1501 1802 1538
rect 1811 1481 1812 1502
rect 1953 1481 1954 1502
rect 1813 1503 1814 1538
rect 1825 1481 1826 1504
rect 1816 1505 1817 1538
rect 1834 1481 1835 1506
rect 1819 1507 1820 1538
rect 1849 1507 1850 1538
rect 1825 1509 1826 1538
rect 1843 1481 1844 1510
rect 1831 1511 1832 1538
rect 1834 1511 1835 1538
rect 1846 1511 1847 1538
rect 1852 1481 1853 1512
rect 1855 1481 1856 1512
rect 1861 1511 1862 1538
rect 1858 1511 1859 1538
rect 1858 1481 1859 1512
rect 1867 1481 1868 1512
rect 1882 1481 1883 1512
rect 1870 1513 1871 1538
rect 1873 1481 1874 1514
rect 1876 1513 1877 1538
rect 1922 1481 1923 1514
rect 1894 1515 1895 1538
rect 1904 1481 1905 1516
rect 1898 1481 1899 1518
rect 1912 1517 1913 1538
rect 1901 1481 1902 1520
rect 1915 1519 1916 1538
rect 1900 1521 1901 1538
rect 1931 1481 1932 1522
rect 1928 1481 1929 1524
rect 1948 1523 1949 1538
rect 1934 1481 1935 1526
rect 1961 1525 1962 1538
rect 1945 1527 1946 1538
rect 1963 1481 1964 1528
rect 1975 1481 1976 1528
rect 1989 1527 1990 1538
rect 1977 1529 1978 1538
rect 1978 1481 1979 1530
rect 1987 1481 1988 1530
rect 2001 1529 2002 1538
rect 1972 1481 1973 1532
rect 1986 1531 1987 1538
rect 1998 1531 1999 1538
rect 2008 1481 2009 1532
rect 2005 1481 2006 1534
rect 2028 1481 2029 1534
rect 2021 1535 2022 1538
rect 2025 1535 2026 1538
rect 2028 1535 2029 1538
rect 2032 1535 2033 1538
rect 1693 1542 1694 1545
rect 1861 1542 1862 1545
rect 1706 1546 1707 1611
rect 1719 1546 1720 1611
rect 1728 1546 1729 1611
rect 1764 1542 1765 1547
rect 1730 1542 1731 1549
rect 1737 1542 1738 1549
rect 1738 1550 1739 1611
rect 1748 1550 1749 1611
rect 1745 1552 1746 1611
rect 1759 1552 1760 1611
rect 1779 1552 1780 1611
rect 1804 1542 1805 1553
rect 1791 1554 1792 1611
rect 1801 1542 1802 1555
rect 1795 1542 1796 1557
rect 1813 1542 1814 1557
rect 1810 1542 1811 1559
rect 1825 1542 1826 1559
rect 1813 1560 1814 1611
rect 1822 1542 1823 1561
rect 1816 1542 1817 1563
rect 1837 1562 1838 1611
rect 1816 1564 1817 1611
rect 1849 1542 1850 1565
rect 1822 1566 1823 1611
rect 1834 1542 1835 1567
rect 1825 1568 1826 1611
rect 1858 1542 1859 1569
rect 1828 1570 1829 1611
rect 1864 1542 1865 1571
rect 1831 1572 1832 1611
rect 1876 1542 1877 1573
rect 1844 1574 1845 1611
rect 1945 1542 1946 1575
rect 1846 1542 1847 1577
rect 1972 1576 1973 1611
rect 1856 1578 1857 1611
rect 1965 1542 1966 1579
rect 1870 1542 1871 1581
rect 1933 1542 1934 1581
rect 1871 1582 1872 1611
rect 1912 1542 1913 1583
rect 1874 1584 1875 1611
rect 1915 1542 1916 1585
rect 1883 1586 1884 1611
rect 1948 1542 1949 1587
rect 1886 1588 1887 1611
rect 1900 1542 1901 1589
rect 1894 1542 1895 1591
rect 1921 1590 1922 1611
rect 1895 1592 1896 1611
rect 1979 1592 1980 1611
rect 1898 1594 1899 1611
rect 1939 1542 1940 1595
rect 1901 1596 1902 1611
rect 1942 1542 1943 1597
rect 1931 1598 1932 1611
rect 1977 1542 1978 1599
rect 1934 1600 1935 1611
rect 1986 1542 1987 1601
rect 1936 1542 1937 1603
rect 2018 1542 2019 1603
rect 1949 1604 1950 1611
rect 1998 1542 1999 1605
rect 1952 1606 1953 1611
rect 2001 1542 2002 1607
rect 1989 1542 1990 1609
rect 2007 1542 2008 1609
rect 1699 1615 1700 1618
rect 1706 1615 1707 1618
rect 1713 1615 1714 1618
rect 1719 1615 1720 1618
rect 1725 1615 1726 1618
rect 1738 1615 1739 1618
rect 1728 1615 1729 1620
rect 1748 1619 1749 1656
rect 1752 1615 1753 1620
rect 1782 1615 1783 1620
rect 1722 1615 1723 1622
rect 1751 1621 1752 1656
rect 1755 1615 1756 1622
rect 1764 1621 1765 1656
rect 1762 1615 1763 1624
rect 1769 1615 1770 1624
rect 1779 1615 1780 1624
rect 1794 1623 1795 1656
rect 1785 1615 1786 1626
rect 1828 1615 1829 1626
rect 1791 1615 1792 1628
rect 1809 1627 1810 1656
rect 1801 1615 1802 1630
rect 1816 1615 1817 1630
rect 1776 1615 1777 1632
rect 1800 1631 1801 1656
rect 1775 1633 1776 1656
rect 1797 1633 1798 1656
rect 1813 1615 1814 1634
rect 1819 1615 1820 1634
rect 1825 1615 1826 1634
rect 1911 1615 1912 1634
rect 1831 1615 1832 1636
rect 1860 1635 1861 1656
rect 1871 1615 1872 1636
rect 1907 1615 1908 1636
rect 1874 1615 1875 1638
rect 1880 1615 1881 1638
rect 1883 1615 1884 1638
rect 1912 1637 1913 1656
rect 1886 1615 1887 1640
rect 1888 1639 1889 1656
rect 1895 1615 1896 1640
rect 1914 1615 1915 1640
rect 1894 1641 1895 1656
rect 1944 1641 1945 1656
rect 1901 1615 1902 1644
rect 1903 1643 1904 1656
rect 1898 1615 1899 1646
rect 1900 1645 1901 1656
rect 1856 1615 1857 1648
rect 1897 1647 1898 1656
rect 1915 1647 1916 1656
rect 1928 1615 1929 1648
rect 1928 1649 1929 1656
rect 1949 1615 1950 1650
rect 1931 1615 1932 1652
rect 1957 1651 1958 1656
rect 1934 1615 1935 1654
rect 1938 1653 1939 1656
rect 1952 1615 1953 1654
rect 1954 1653 1955 1656
rect 1711 1662 1712 1699
rect 1748 1660 1749 1663
rect 1723 1664 1724 1699
rect 1751 1660 1752 1665
rect 1757 1660 1758 1665
rect 1764 1660 1765 1665
rect 1759 1666 1760 1699
rect 1761 1660 1762 1667
rect 1763 1666 1764 1699
rect 1797 1660 1798 1667
rect 1766 1668 1767 1699
rect 1809 1660 1810 1669
rect 1778 1660 1779 1671
rect 1800 1660 1801 1671
rect 1794 1660 1795 1673
rect 1815 1660 1816 1673
rect 1801 1674 1802 1699
rect 1957 1660 1958 1675
rect 1804 1676 1805 1699
rect 1822 1660 1823 1677
rect 1826 1660 1827 1677
rect 1833 1660 1834 1677
rect 1841 1676 1842 1699
rect 1860 1660 1861 1677
rect 1857 1678 1858 1699
rect 1903 1660 1904 1679
rect 1863 1680 1864 1699
rect 1897 1660 1898 1681
rect 1878 1682 1879 1699
rect 1915 1660 1916 1683
rect 1881 1684 1882 1699
rect 1888 1660 1889 1685
rect 1884 1686 1885 1699
rect 1918 1660 1919 1687
rect 1887 1688 1888 1699
rect 1900 1660 1901 1689
rect 1894 1660 1895 1691
rect 1935 1660 1936 1691
rect 1910 1692 1911 1699
rect 1938 1660 1939 1693
rect 1912 1660 1913 1695
rect 1948 1660 1949 1695
rect 1941 1660 1942 1697
rect 1954 1660 1955 1697
rect 1969 1660 1970 1697
rect 1976 1660 1977 1697
rect 1711 1703 1712 1706
rect 1717 1705 1718 1720
rect 1720 1705 1721 1720
rect 1723 1703 1724 1706
rect 1759 1703 1760 1706
rect 1763 1703 1764 1706
rect 1804 1705 1805 1720
rect 1804 1703 1805 1706
rect 1834 1705 1835 1720
rect 1847 1705 1848 1720
rect 1837 1707 1838 1720
rect 1841 1703 1842 1708
rect 1857 1703 1858 1708
rect 1913 1703 1914 1708
rect 1863 1703 1864 1710
rect 1904 1703 1905 1710
rect 1872 1711 1873 1720
rect 1884 1703 1885 1712
rect 1875 1713 1876 1720
rect 1887 1703 1888 1714
rect 1878 1703 1879 1716
rect 1907 1703 1908 1716
rect 1878 1717 1879 1720
rect 1900 1703 1901 1718
rect 1881 1717 1882 1720
rect 1881 1703 1882 1718
rect 1904 1717 1905 1720
rect 1910 1703 1911 1718
rect 1916 1703 1917 1718
rect 1937 1703 1938 1718
rect 1711 1724 1712 1727
rect 1717 1724 1718 1727
rect 1720 1724 1721 1727
rect 1749 1724 1750 1727
rect 1770 1726 1771 1745
rect 1784 1726 1785 1745
rect 1804 1724 1805 1727
rect 1831 1724 1832 1727
rect 1780 1724 1781 1729
rect 1804 1728 1805 1745
rect 1780 1730 1781 1745
rect 1791 1730 1792 1745
rect 1831 1730 1832 1745
rect 1881 1724 1882 1731
rect 1834 1724 1835 1733
rect 1843 1724 1844 1733
rect 1834 1734 1835 1745
rect 1840 1734 1841 1745
rect 1837 1724 1838 1737
rect 1907 1724 1908 1737
rect 1847 1724 1848 1739
rect 1857 1724 1858 1739
rect 1863 1738 1864 1745
rect 1872 1724 1873 1739
rect 1866 1740 1867 1745
rect 1875 1724 1876 1741
rect 1869 1742 1870 1745
rect 1878 1724 1879 1743
rect 1892 1742 1893 1745
rect 1904 1724 1905 1743
rect 1681 1749 1682 1752
rect 1688 1749 1689 1752
rect 1780 1749 1781 1752
rect 1784 1749 1785 1752
rect 1801 1749 1802 1752
rect 1804 1749 1805 1752
rect 1810 1749 1811 1752
rect 1811 1751 1812 1758
rect 1827 1751 1828 1758
rect 1831 1749 1832 1752
rect 1834 1749 1835 1752
rect 1836 1751 1837 1758
rect 1869 1749 1870 1752
rect 1871 1751 1872 1758
rect 1866 1749 1867 1754
rect 1868 1753 1869 1758
rect 1863 1749 1864 1756
rect 1865 1755 1866 1758
rect 1892 1749 1893 1756
rect 1898 1749 1899 1756
rect 1811 1764 1812 1767
rect 1811 1762 1812 1765
rect 1827 1764 1828 1767
rect 1827 1762 1828 1765
rect 1836 1764 1837 1767
rect 1836 1762 1837 1765
rect 1865 1764 1866 1767
rect 1865 1762 1866 1765
rect 1868 1764 1869 1767
rect 1868 1762 1869 1765
rect 1871 1764 1872 1767
rect 1871 1762 1872 1765
rect 1811 1773 1812 1776
rect 1811 1771 1812 1774
rect 1827 1773 1828 1776
rect 1827 1771 1828 1774
rect 1836 1773 1837 1776
rect 1836 1771 1837 1774
rect 1865 1773 1866 1776
rect 1865 1771 1866 1774
rect 1868 1773 1869 1776
rect 1868 1771 1869 1774
rect 1871 1773 1872 1776
rect 1871 1771 1872 1774
rect 1714 1782 1715 1795
rect 1868 1780 1869 1783
rect 1801 1784 1802 1795
rect 1811 1780 1812 1785
rect 1810 1786 1811 1795
rect 1827 1780 1828 1787
rect 1819 1788 1820 1795
rect 1836 1780 1837 1789
rect 1837 1790 1838 1795
rect 1865 1780 1866 1791
rect 1840 1792 1841 1795
rect 1871 1780 1872 1793
rect 1714 1799 1715 1802
rect 1718 1799 1719 1802
rect 1762 1799 1763 1802
rect 1840 1799 1841 1802
rect 1774 1799 1775 1804
rect 1801 1799 1802 1804
rect 1795 1799 1796 1806
rect 1837 1799 1838 1806
rect 1810 1799 1811 1808
rect 1813 1799 1814 1808
rect 1819 1799 1820 1808
rect 1822 1799 1823 1808
<< via >>
rect 1783 833 1784 834
rect 1786 833 1787 834
rect 1813 833 1814 834
rect 1819 833 1820 834
rect 1822 833 1823 834
rect 1828 833 1829 834
rect 1753 843 1754 844
rect 1755 843 1756 844
rect 1783 843 1784 844
rect 1808 843 1809 844
rect 1792 845 1793 846
rect 1817 845 1818 846
rect 1766 847 1767 848
rect 1792 847 1793 848
rect 1813 847 1814 848
rect 1833 847 1834 848
rect 1822 849 1823 850
rect 1842 849 1843 850
rect 1717 876 1718 877
rect 1865 876 1866 877
rect 1919 876 1920 877
rect 1926 876 1927 877
rect 1720 885 1721 886
rect 1892 885 1893 886
rect 1721 887 1722 888
rect 1724 887 1725 888
rect 1755 887 1756 888
rect 1757 887 1758 888
rect 1727 889 1728 890
rect 1754 889 1755 890
rect 1770 889 1771 890
rect 1794 889 1795 890
rect 1792 891 1793 892
rect 1797 891 1798 892
rect 1808 891 1809 892
rect 1813 891 1814 892
rect 1817 891 1818 892
rect 1822 891 1823 892
rect 1842 891 1843 892
rect 1845 891 1846 892
rect 1833 893 1834 894
rect 1842 893 1843 894
rect 1865 893 1866 894
rect 1873 893 1874 894
rect 1876 893 1877 894
rect 1915 893 1916 894
rect 1878 895 1879 896
rect 1895 895 1896 896
rect 1912 895 1913 896
rect 1925 895 1926 896
rect 1922 897 1923 898
rect 1931 897 1932 898
rect 1711 906 1712 907
rect 1724 906 1725 907
rect 1735 906 1736 907
rect 1841 906 1842 907
rect 1745 908 1746 909
rect 1752 908 1753 909
rect 1803 908 1804 909
rect 1820 908 1821 909
rect 1792 910 1793 911
rect 1804 910 1805 911
rect 1822 910 1823 911
rect 1832 910 1833 911
rect 1813 912 1814 913
rect 1823 912 1824 913
rect 1845 912 1846 913
rect 1851 912 1852 913
rect 1873 912 1874 913
rect 1885 912 1886 913
rect 1876 914 1877 915
rect 1888 914 1889 915
rect 1895 914 1896 915
rect 1914 914 1915 915
rect 1912 916 1913 917
rect 1920 916 1921 917
rect 1892 918 1893 919
rect 1911 918 1912 919
rect 1857 920 1858 921
rect 1891 920 1892 921
rect 1925 920 1926 921
rect 1938 920 1939 921
rect 1737 922 1738 923
rect 1938 922 1939 923
rect 1738 924 1739 925
rect 1754 924 1755 925
rect 1727 926 1728 927
rect 1755 926 1756 927
rect 1721 935 1722 936
rect 1725 935 1726 936
rect 1737 935 1738 936
rect 1755 935 1756 936
rect 1753 937 1754 938
rect 1758 937 1759 938
rect 1776 937 1777 938
rect 1795 937 1796 938
rect 1785 939 1786 940
rect 1798 939 1799 940
rect 1795 941 1796 942
rect 1823 941 1824 942
rect 1801 943 1802 944
rect 1820 943 1821 944
rect 1811 945 1812 946
rect 1832 945 1833 946
rect 1817 947 1818 948
rect 1860 947 1861 948
rect 1826 949 1827 950
rect 1841 949 1842 950
rect 1829 951 1830 952
rect 1841 951 1842 952
rect 1838 953 1839 954
rect 1857 953 1858 954
rect 1847 955 1848 956
rect 1894 955 1895 956
rect 1854 957 1855 958
rect 1872 957 1873 958
rect 1866 959 1867 960
rect 1888 959 1889 960
rect 1882 961 1883 962
rect 1944 961 1945 962
rect 1881 963 1882 964
rect 1959 963 1960 964
rect 1885 965 1886 966
rect 1890 965 1891 966
rect 1893 965 1894 966
rect 1938 965 1939 966
rect 1896 967 1897 968
rect 1921 967 1922 968
rect 1908 969 1909 970
rect 1914 969 1915 970
rect 1966 969 1967 970
rect 1973 969 1974 970
rect 1714 978 1715 979
rect 1718 978 1719 979
rect 1729 978 1730 979
rect 1771 978 1772 979
rect 1737 980 1738 981
rect 1749 980 1750 981
rect 1746 982 1747 983
rect 1758 982 1759 983
rect 1753 984 1754 985
rect 1761 984 1762 985
rect 1764 984 1765 985
rect 1803 984 1804 985
rect 1801 986 1802 987
rect 1822 986 1823 987
rect 1826 986 1827 987
rect 1849 986 1850 987
rect 1829 988 1830 989
rect 1852 988 1853 989
rect 1828 990 1829 991
rect 1840 990 1841 991
rect 1838 992 1839 993
rect 1860 992 1861 993
rect 1817 994 1818 995
rect 1837 994 1838 995
rect 1809 996 1810 997
rect 1816 996 1817 997
rect 1861 996 1862 997
rect 1874 996 1875 997
rect 1866 998 1867 999
rect 1884 998 1885 999
rect 1872 1000 1873 1001
rect 1941 1000 1942 1001
rect 1881 1002 1882 1003
rect 1928 1002 1929 1003
rect 1807 1004 1808 1005
rect 1929 1004 1930 1005
rect 1785 1006 1786 1007
rect 1806 1006 1807 1007
rect 1776 1008 1777 1009
rect 1784 1008 1785 1009
rect 1847 1008 1848 1009
rect 1881 1008 1882 1009
rect 1800 1010 1801 1011
rect 1846 1010 1847 1011
rect 1890 1010 1891 1011
rect 1948 1010 1949 1011
rect 1856 1012 1857 1013
rect 1890 1012 1891 1013
rect 1893 1012 1894 1013
rect 1920 1012 1921 1013
rect 1896 1014 1897 1015
rect 1923 1014 1924 1015
rect 1899 1016 1900 1017
rect 1926 1016 1927 1017
rect 1899 1018 1900 1019
rect 1902 1018 1903 1019
rect 1908 1018 1909 1019
rect 1932 1018 1933 1019
rect 1911 1020 1912 1021
rect 1935 1020 1936 1021
rect 1914 1022 1915 1023
rect 1917 1022 1918 1023
rect 1938 1022 1939 1023
rect 1993 1022 1994 1023
rect 1743 1031 1744 1032
rect 1770 1031 1771 1032
rect 1732 1033 1733 1034
rect 1742 1033 1743 1034
rect 1749 1033 1750 1034
rect 1764 1033 1765 1034
rect 1748 1035 1749 1036
rect 1752 1035 1753 1036
rect 1758 1035 1759 1036
rect 1767 1035 1768 1036
rect 1758 1037 1759 1038
rect 1761 1037 1762 1038
rect 1790 1037 1791 1038
rect 2032 1037 2033 1038
rect 1819 1039 1820 1040
rect 1828 1039 1829 1040
rect 1806 1041 1807 1042
rect 1829 1041 1830 1042
rect 1784 1043 1785 1044
rect 1807 1043 1808 1044
rect 1822 1043 1823 1044
rect 1856 1043 1857 1044
rect 1837 1045 1838 1046
rect 1847 1045 1848 1046
rect 1852 1045 1853 1046
rect 1886 1045 1887 1046
rect 1803 1047 1804 1048
rect 1853 1047 1854 1048
rect 1804 1049 1805 1050
rect 1838 1049 1839 1050
rect 1858 1049 1859 1050
rect 1892 1049 1893 1050
rect 1810 1051 1811 1052
rect 1859 1051 1860 1052
rect 1861 1051 1862 1052
rect 1867 1051 1868 1052
rect 1840 1053 1841 1054
rect 1868 1053 1869 1054
rect 1864 1055 1865 1056
rect 1901 1055 1902 1056
rect 1871 1057 1872 1058
rect 1878 1057 1879 1058
rect 1890 1057 1891 1058
rect 1944 1057 1945 1058
rect 1849 1059 1850 1060
rect 1889 1059 1890 1060
rect 1797 1061 1798 1062
rect 1850 1061 1851 1062
rect 1797 1063 1798 1064
rect 1800 1063 1801 1064
rect 1899 1063 1900 1064
rect 1948 1063 1949 1064
rect 1917 1065 1918 1066
rect 1972 1065 1973 1066
rect 1884 1067 1885 1068
rect 1917 1067 1918 1068
rect 1920 1067 1921 1068
rect 1975 1067 1976 1068
rect 1926 1069 1927 1070
rect 1981 1069 1982 1070
rect 1929 1071 1930 1072
rect 1984 1071 1985 1072
rect 1929 1073 1930 1074
rect 1938 1073 1939 1074
rect 1932 1075 1933 1076
rect 1986 1075 1987 1076
rect 1932 1077 1933 1078
rect 2025 1077 2026 1078
rect 1935 1079 1936 1080
rect 1979 1079 1980 1080
rect 1923 1081 1924 1082
rect 1978 1081 1979 1082
rect 1923 1083 1924 1084
rect 1994 1083 1995 1084
rect 1954 1085 1955 1086
rect 1990 1085 1991 1086
rect 2004 1085 2005 1086
rect 2008 1085 2009 1086
rect 1729 1094 1730 1095
rect 1739 1094 1740 1095
rect 1729 1096 1730 1097
rect 1847 1096 1848 1097
rect 1742 1098 1743 1099
rect 1745 1098 1746 1099
rect 1743 1100 1744 1101
rect 1750 1100 1751 1101
rect 1758 1100 1759 1101
rect 1789 1100 1790 1101
rect 1767 1102 1768 1103
rect 1783 1102 1784 1103
rect 1767 1104 1768 1105
rect 1838 1104 1839 1105
rect 1773 1106 1774 1107
rect 1780 1106 1781 1107
rect 1776 1108 1777 1109
rect 1826 1108 1827 1109
rect 1802 1110 1803 1111
rect 1880 1110 1881 1111
rect 1807 1112 1808 1113
rect 1838 1112 1839 1113
rect 1820 1114 1821 1115
rect 1874 1114 1875 1115
rect 1823 1116 1824 1117
rect 1871 1116 1872 1117
rect 1853 1118 1854 1119
rect 1862 1118 1863 1119
rect 1856 1120 1857 1121
rect 1883 1120 1884 1121
rect 1868 1122 1869 1123
rect 1895 1122 1896 1123
rect 1886 1124 1887 1125
rect 1968 1124 1969 1125
rect 1859 1126 1860 1127
rect 1886 1126 1887 1127
rect 1829 1128 1830 1129
rect 1859 1128 1860 1129
rect 1792 1130 1793 1131
rect 1829 1130 1830 1131
rect 1889 1130 1890 1131
rect 1919 1130 1920 1131
rect 1889 1132 1890 1133
rect 1925 1132 1926 1133
rect 1917 1134 1918 1135
rect 1934 1134 1935 1135
rect 1898 1136 1899 1137
rect 1916 1136 1917 1137
rect 1844 1138 1845 1139
rect 1898 1138 1899 1139
rect 1923 1138 1924 1139
rect 1940 1138 1941 1139
rect 1901 1140 1902 1141
rect 1922 1140 1923 1141
rect 1877 1142 1878 1143
rect 1901 1142 1902 1143
rect 1850 1144 1851 1145
rect 1877 1144 1878 1145
rect 1770 1146 1771 1147
rect 1850 1146 1851 1147
rect 1929 1146 1930 1147
rect 2047 1146 2048 1147
rect 1932 1148 1933 1149
rect 1959 1148 1960 1149
rect 1904 1150 1905 1151
rect 1931 1150 1932 1151
rect 1892 1152 1893 1153
rect 1904 1152 1905 1153
rect 1948 1152 1949 1153
rect 1962 1152 1963 1153
rect 1975 1152 1976 1153
rect 2004 1152 2005 1153
rect 1954 1154 1955 1155
rect 1974 1154 1975 1155
rect 1978 1154 1979 1155
rect 2010 1154 2011 1155
rect 1981 1156 1982 1157
rect 2013 1156 2014 1157
rect 1984 1158 1985 1159
rect 2007 1158 2008 1159
rect 1986 1160 1987 1161
rect 2068 1160 2069 1161
rect 1994 1162 1995 1163
rect 2001 1162 2002 1163
rect 1972 1164 1973 1165
rect 2001 1164 2002 1165
rect 2040 1164 2041 1165
rect 2054 1164 2055 1165
rect 2051 1166 2052 1167
rect 2065 1166 2066 1167
rect 1743 1175 1744 1176
rect 1847 1175 1848 1176
rect 1746 1177 1747 1178
rect 1826 1177 1827 1178
rect 1755 1179 1756 1180
rect 1789 1179 1790 1180
rect 1757 1181 1758 1182
rect 1785 1181 1786 1182
rect 1761 1183 1762 1184
rect 1768 1183 1769 1184
rect 1764 1185 1765 1186
rect 1850 1185 1851 1186
rect 1765 1187 1766 1188
rect 1783 1187 1784 1188
rect 1771 1189 1772 1190
rect 1821 1189 1822 1190
rect 1775 1191 1776 1192
rect 1782 1191 1783 1192
rect 1779 1193 1780 1194
rect 1880 1193 1881 1194
rect 1788 1195 1789 1196
rect 1827 1195 1828 1196
rect 1806 1197 1807 1198
rect 1824 1197 1825 1198
rect 1806 1199 1807 1200
rect 1829 1199 1830 1200
rect 1812 1201 1813 1202
rect 1862 1201 1863 1202
rect 1816 1203 1817 1204
rect 1883 1203 1884 1204
rect 1818 1205 1819 1206
rect 1859 1205 1860 1206
rect 1830 1207 1831 1208
rect 1857 1207 1858 1208
rect 1838 1209 1839 1210
rect 2061 1209 2062 1210
rect 1839 1211 1840 1212
rect 1877 1211 1878 1212
rect 1841 1213 1842 1214
rect 1889 1213 1890 1214
rect 1842 1215 1843 1216
rect 1944 1215 1945 1216
rect 1844 1217 1845 1218
rect 1901 1217 1902 1218
rect 1845 1219 1846 1220
rect 1886 1219 1887 1220
rect 1860 1221 1861 1222
rect 1874 1221 1875 1222
rect 1866 1223 1867 1224
rect 1895 1223 1896 1224
rect 1875 1225 1876 1226
rect 1904 1225 1905 1226
rect 1887 1227 1888 1228
rect 1981 1227 1982 1228
rect 1893 1229 1894 1230
rect 1916 1229 1917 1230
rect 1896 1231 1897 1232
rect 1919 1231 1920 1232
rect 1911 1233 1912 1234
rect 1931 1233 1932 1234
rect 1914 1235 1915 1236
rect 1946 1235 1947 1236
rect 1917 1237 1918 1238
rect 1934 1237 1935 1238
rect 1922 1239 1923 1240
rect 1953 1239 1954 1240
rect 1923 1241 1924 1242
rect 1940 1241 1941 1242
rect 1928 1243 1929 1244
rect 1932 1243 1933 1244
rect 1935 1243 1936 1244
rect 2019 1243 2020 1244
rect 1959 1245 1960 1246
rect 1978 1245 1979 1246
rect 1960 1247 1961 1248
rect 2058 1247 2059 1248
rect 1962 1249 1963 1250
rect 2016 1249 2017 1250
rect 1863 1251 1864 1252
rect 2017 1251 2018 1252
rect 1963 1253 1964 1254
rect 2068 1253 2069 1254
rect 1972 1255 1973 1256
rect 2004 1255 2005 1256
rect 1986 1257 1987 1258
rect 2044 1257 2045 1258
rect 1991 1259 1992 1260
rect 2007 1259 2008 1260
rect 1995 1261 1996 1262
rect 2001 1261 2002 1262
rect 1994 1263 1995 1264
rect 2010 1263 2011 1264
rect 1997 1265 1998 1266
rect 2013 1265 2014 1266
rect 1717 1274 1718 1275
rect 1724 1274 1725 1275
rect 1748 1274 1749 1275
rect 1752 1274 1753 1275
rect 1755 1274 1756 1275
rect 1758 1274 1759 1275
rect 1761 1274 1762 1275
rect 1797 1274 1798 1275
rect 1768 1276 1769 1277
rect 1821 1276 1822 1277
rect 1767 1278 1768 1279
rect 1785 1278 1786 1279
rect 1782 1280 1783 1281
rect 1824 1280 1825 1281
rect 1788 1282 1789 1283
rect 1842 1282 1843 1283
rect 1791 1284 1792 1285
rect 1830 1284 1831 1285
rect 1812 1286 1813 1287
rect 1833 1286 1834 1287
rect 1812 1288 1813 1289
rect 1818 1288 1819 1289
rect 1815 1290 1816 1291
rect 1981 1290 1982 1291
rect 1836 1292 1837 1293
rect 1860 1292 1861 1293
rect 1839 1294 1840 1295
rect 1872 1294 1873 1295
rect 1842 1296 1843 1297
rect 1863 1296 1864 1297
rect 1845 1298 1846 1299
rect 1866 1298 1867 1299
rect 1857 1300 1858 1301
rect 1948 1300 1949 1301
rect 1860 1302 1861 1303
rect 1896 1302 1897 1303
rect 1863 1304 1864 1305
rect 1875 1304 1876 1305
rect 1878 1304 1879 1305
rect 1978 1304 1979 1305
rect 1881 1306 1882 1307
rect 1911 1306 1912 1307
rect 1884 1308 1885 1309
rect 1887 1308 1888 1309
rect 1893 1308 1894 1309
rect 2010 1308 2011 1309
rect 1900 1310 1901 1311
rect 1917 1310 1918 1311
rect 1914 1312 1915 1313
rect 1929 1312 1930 1313
rect 1923 1314 1924 1315
rect 1933 1314 1934 1315
rect 1924 1316 1925 1317
rect 1975 1316 1976 1317
rect 1927 1318 1928 1319
rect 1935 1318 1936 1319
rect 1930 1320 1931 1321
rect 1997 1320 1998 1321
rect 1946 1322 1947 1323
rect 1972 1322 1973 1323
rect 1951 1324 1952 1325
rect 1963 1324 1964 1325
rect 1950 1326 1951 1327
rect 1979 1326 1980 1327
rect 1956 1328 1957 1329
rect 1991 1328 1992 1329
rect 1960 1330 1961 1331
rect 2035 1330 2036 1331
rect 1982 1332 1983 1333
rect 1994 1332 1995 1333
rect 1741 1341 1742 1342
rect 1764 1341 1765 1342
rect 1748 1343 1749 1344
rect 1761 1343 1762 1344
rect 1752 1345 1753 1346
rect 1784 1345 1785 1346
rect 1767 1347 1768 1348
rect 1790 1347 1791 1348
rect 1758 1349 1759 1350
rect 1767 1349 1768 1350
rect 1773 1349 1774 1350
rect 1997 1349 1998 1350
rect 1793 1351 1794 1352
rect 1840 1351 1841 1352
rect 1797 1353 1798 1354
rect 1819 1353 1820 1354
rect 1812 1355 1813 1356
rect 1828 1355 1829 1356
rect 1824 1357 1825 1358
rect 1881 1357 1882 1358
rect 1830 1359 1831 1360
rect 1843 1359 1844 1360
rect 1815 1361 1816 1362
rect 1831 1361 1832 1362
rect 1833 1361 1834 1362
rect 1852 1361 1853 1362
rect 1836 1363 1837 1364
rect 1855 1363 1856 1364
rect 1849 1365 1850 1366
rect 1887 1365 1888 1366
rect 1863 1367 1864 1368
rect 1882 1367 1883 1368
rect 1845 1369 1846 1370
rect 1864 1369 1865 1370
rect 1875 1369 1876 1370
rect 1935 1369 1936 1370
rect 1878 1371 1879 1372
rect 1894 1371 1895 1372
rect 1860 1373 1861 1374
rect 1879 1373 1880 1374
rect 1888 1373 1889 1374
rect 1939 1373 1940 1374
rect 1915 1375 1916 1376
rect 1938 1375 1939 1376
rect 1914 1377 1915 1378
rect 1950 1377 1951 1378
rect 1924 1379 1925 1380
rect 1965 1379 1966 1380
rect 1900 1381 1901 1382
rect 1923 1381 1924 1382
rect 1927 1381 1928 1382
rect 1968 1381 1969 1382
rect 1930 1383 1931 1384
rect 1953 1383 1954 1384
rect 1943 1385 1944 1386
rect 2018 1385 2019 1386
rect 1956 1387 1957 1388
rect 2000 1387 2001 1388
rect 1933 1389 1934 1390
rect 1956 1389 1957 1390
rect 1979 1389 1980 1390
rect 2021 1389 2022 1390
rect 2009 1391 2010 1392
rect 2041 1391 2042 1392
rect 1729 1400 1730 1401
rect 1736 1400 1737 1401
rect 1740 1400 1741 1401
rect 1761 1400 1762 1401
rect 1744 1402 1745 1403
rect 1793 1402 1794 1403
rect 1751 1404 1752 1405
rect 1843 1404 1844 1405
rect 1755 1406 1756 1407
rect 1808 1406 1809 1407
rect 1761 1408 1762 1409
rect 1828 1408 1829 1409
rect 1764 1410 1765 1411
rect 1780 1410 1781 1411
rect 1767 1412 1768 1413
rect 1837 1412 1838 1413
rect 1768 1414 1769 1415
rect 1831 1414 1832 1415
rect 1778 1416 1779 1417
rect 1790 1416 1791 1417
rect 1800 1416 1801 1417
rect 1849 1416 1850 1417
rect 1805 1418 1806 1419
rect 1819 1418 1820 1419
rect 1831 1418 1832 1419
rect 1852 1418 1853 1419
rect 1834 1420 1835 1421
rect 1840 1420 1841 1421
rect 1840 1422 1841 1423
rect 1858 1422 1859 1423
rect 1843 1424 1844 1425
rect 1855 1424 1856 1425
rect 1852 1426 1853 1427
rect 1864 1426 1865 1427
rect 1855 1428 1856 1429
rect 1867 1428 1868 1429
rect 1861 1430 1862 1431
rect 1879 1430 1880 1431
rect 1867 1432 1868 1433
rect 1885 1432 1886 1433
rect 1870 1434 1871 1435
rect 1886 1434 1887 1435
rect 1873 1436 1874 1437
rect 1888 1436 1889 1437
rect 1882 1438 1883 1439
rect 1962 1438 1963 1439
rect 1821 1440 1822 1441
rect 1882 1440 1883 1441
rect 1894 1440 1895 1441
rect 1971 1440 1972 1441
rect 1898 1442 1899 1443
rect 1935 1442 1936 1443
rect 1901 1444 1902 1445
rect 1938 1444 1939 1445
rect 1904 1446 1905 1447
rect 1923 1446 1924 1447
rect 1907 1448 1908 1449
rect 1947 1448 1948 1449
rect 1928 1450 1929 1451
rect 1953 1450 1954 1451
rect 1931 1452 1932 1453
rect 1956 1452 1957 1453
rect 1934 1454 1935 1455
rect 1949 1454 1950 1455
rect 1937 1456 1938 1457
rect 1965 1456 1966 1457
rect 1940 1458 1941 1459
rect 1968 1458 1969 1459
rect 1943 1460 1944 1461
rect 2024 1460 2025 1461
rect 1972 1462 1973 1463
rect 1997 1462 1998 1463
rect 1975 1464 1976 1465
rect 2000 1464 2001 1465
rect 1978 1466 1979 1467
rect 2041 1466 2042 1467
rect 1987 1468 1988 1469
rect 2038 1468 2039 1469
rect 2018 1470 2019 1471
rect 2034 1470 2035 1471
rect 2005 1472 2006 1473
rect 2035 1472 2036 1473
rect 2021 1474 2022 1475
rect 2031 1474 2032 1475
rect 1696 1483 1697 1484
rect 1870 1483 1871 1484
rect 1723 1485 1724 1486
rect 1733 1485 1734 1486
rect 1730 1487 1731 1488
rect 1737 1487 1738 1488
rect 1723 1489 1724 1490
rect 1730 1489 1731 1490
rect 1744 1489 1745 1490
rect 1808 1489 1809 1490
rect 1744 1491 1745 1492
rect 1793 1491 1794 1492
rect 1747 1493 1748 1494
rect 1805 1493 1806 1494
rect 1751 1495 1752 1496
rect 1788 1495 1789 1496
rect 1765 1497 1766 1498
rect 1804 1497 1805 1498
rect 1764 1499 1765 1500
rect 1778 1499 1779 1500
rect 1791 1499 1792 1500
rect 1831 1499 1832 1500
rect 1799 1501 1800 1502
rect 1801 1501 1802 1502
rect 1811 1501 1812 1502
rect 1953 1501 1954 1502
rect 1813 1503 1814 1504
rect 1825 1503 1826 1504
rect 1816 1505 1817 1506
rect 1834 1505 1835 1506
rect 1819 1507 1820 1508
rect 1849 1507 1850 1508
rect 1825 1509 1826 1510
rect 1843 1509 1844 1510
rect 1831 1511 1832 1512
rect 1834 1511 1835 1512
rect 1846 1511 1847 1512
rect 1852 1511 1853 1512
rect 1855 1511 1856 1512
rect 1861 1511 1862 1512
rect 1867 1511 1868 1512
rect 1882 1511 1883 1512
rect 1870 1513 1871 1514
rect 1873 1513 1874 1514
rect 1876 1513 1877 1514
rect 1922 1513 1923 1514
rect 1894 1515 1895 1516
rect 1904 1515 1905 1516
rect 1898 1517 1899 1518
rect 1912 1517 1913 1518
rect 1901 1519 1902 1520
rect 1915 1519 1916 1520
rect 1900 1521 1901 1522
rect 1931 1521 1932 1522
rect 1928 1523 1929 1524
rect 1948 1523 1949 1524
rect 1934 1525 1935 1526
rect 1961 1525 1962 1526
rect 1945 1527 1946 1528
rect 1963 1527 1964 1528
rect 1975 1527 1976 1528
rect 1989 1527 1990 1528
rect 1987 1529 1988 1530
rect 2001 1529 2002 1530
rect 1972 1531 1973 1532
rect 1986 1531 1987 1532
rect 1998 1531 1999 1532
rect 2008 1531 2009 1532
rect 2005 1533 2006 1534
rect 2028 1533 2029 1534
rect 2021 1535 2022 1536
rect 2025 1535 2026 1536
rect 2028 1535 2029 1536
rect 2032 1535 2033 1536
rect 1693 1544 1694 1545
rect 1861 1544 1862 1545
rect 1706 1546 1707 1547
rect 1719 1546 1720 1547
rect 1728 1546 1729 1547
rect 1764 1546 1765 1547
rect 1730 1548 1731 1549
rect 1737 1548 1738 1549
rect 1738 1550 1739 1551
rect 1748 1550 1749 1551
rect 1745 1552 1746 1553
rect 1759 1552 1760 1553
rect 1779 1552 1780 1553
rect 1804 1552 1805 1553
rect 1791 1554 1792 1555
rect 1801 1554 1802 1555
rect 1795 1556 1796 1557
rect 1813 1556 1814 1557
rect 1810 1558 1811 1559
rect 1825 1558 1826 1559
rect 1813 1560 1814 1561
rect 1822 1560 1823 1561
rect 1816 1562 1817 1563
rect 1837 1562 1838 1563
rect 1816 1564 1817 1565
rect 1849 1564 1850 1565
rect 1822 1566 1823 1567
rect 1834 1566 1835 1567
rect 1825 1568 1826 1569
rect 1858 1568 1859 1569
rect 1828 1570 1829 1571
rect 1864 1570 1865 1571
rect 1831 1572 1832 1573
rect 1876 1572 1877 1573
rect 1844 1574 1845 1575
rect 1945 1574 1946 1575
rect 1846 1576 1847 1577
rect 1972 1576 1973 1577
rect 1856 1578 1857 1579
rect 1965 1578 1966 1579
rect 1870 1580 1871 1581
rect 1933 1580 1934 1581
rect 1871 1582 1872 1583
rect 1912 1582 1913 1583
rect 1874 1584 1875 1585
rect 1915 1584 1916 1585
rect 1883 1586 1884 1587
rect 1948 1586 1949 1587
rect 1886 1588 1887 1589
rect 1900 1588 1901 1589
rect 1894 1590 1895 1591
rect 1921 1590 1922 1591
rect 1895 1592 1896 1593
rect 1979 1592 1980 1593
rect 1898 1594 1899 1595
rect 1939 1594 1940 1595
rect 1901 1596 1902 1597
rect 1942 1596 1943 1597
rect 1931 1598 1932 1599
rect 1977 1598 1978 1599
rect 1934 1600 1935 1601
rect 1986 1600 1987 1601
rect 1936 1602 1937 1603
rect 2018 1602 2019 1603
rect 1949 1604 1950 1605
rect 1998 1604 1999 1605
rect 1952 1606 1953 1607
rect 2001 1606 2002 1607
rect 1989 1608 1990 1609
rect 2007 1608 2008 1609
rect 1699 1617 1700 1618
rect 1706 1617 1707 1618
rect 1713 1617 1714 1618
rect 1719 1617 1720 1618
rect 1725 1617 1726 1618
rect 1738 1617 1739 1618
rect 1728 1619 1729 1620
rect 1748 1619 1749 1620
rect 1752 1619 1753 1620
rect 1782 1619 1783 1620
rect 1722 1621 1723 1622
rect 1751 1621 1752 1622
rect 1755 1621 1756 1622
rect 1764 1621 1765 1622
rect 1762 1623 1763 1624
rect 1769 1623 1770 1624
rect 1779 1623 1780 1624
rect 1794 1623 1795 1624
rect 1785 1625 1786 1626
rect 1828 1625 1829 1626
rect 1791 1627 1792 1628
rect 1809 1627 1810 1628
rect 1801 1629 1802 1630
rect 1816 1629 1817 1630
rect 1776 1631 1777 1632
rect 1800 1631 1801 1632
rect 1775 1633 1776 1634
rect 1797 1633 1798 1634
rect 1813 1633 1814 1634
rect 1819 1633 1820 1634
rect 1825 1633 1826 1634
rect 1911 1633 1912 1634
rect 1831 1635 1832 1636
rect 1860 1635 1861 1636
rect 1871 1635 1872 1636
rect 1907 1635 1908 1636
rect 1874 1637 1875 1638
rect 1880 1637 1881 1638
rect 1883 1637 1884 1638
rect 1912 1637 1913 1638
rect 1886 1639 1887 1640
rect 1888 1639 1889 1640
rect 1895 1639 1896 1640
rect 1914 1639 1915 1640
rect 1894 1641 1895 1642
rect 1944 1641 1945 1642
rect 1901 1643 1902 1644
rect 1903 1643 1904 1644
rect 1898 1645 1899 1646
rect 1900 1645 1901 1646
rect 1856 1647 1857 1648
rect 1897 1647 1898 1648
rect 1915 1647 1916 1648
rect 1928 1647 1929 1648
rect 1928 1649 1929 1650
rect 1949 1649 1950 1650
rect 1931 1651 1932 1652
rect 1957 1651 1958 1652
rect 1934 1653 1935 1654
rect 1938 1653 1939 1654
rect 1952 1653 1953 1654
rect 1954 1653 1955 1654
rect 1711 1662 1712 1663
rect 1748 1662 1749 1663
rect 1723 1664 1724 1665
rect 1751 1664 1752 1665
rect 1757 1664 1758 1665
rect 1764 1664 1765 1665
rect 1759 1666 1760 1667
rect 1761 1666 1762 1667
rect 1763 1666 1764 1667
rect 1797 1666 1798 1667
rect 1766 1668 1767 1669
rect 1809 1668 1810 1669
rect 1778 1670 1779 1671
rect 1800 1670 1801 1671
rect 1794 1672 1795 1673
rect 1815 1672 1816 1673
rect 1801 1674 1802 1675
rect 1957 1674 1958 1675
rect 1804 1676 1805 1677
rect 1822 1676 1823 1677
rect 1826 1676 1827 1677
rect 1833 1676 1834 1677
rect 1841 1676 1842 1677
rect 1860 1676 1861 1677
rect 1857 1678 1858 1679
rect 1903 1678 1904 1679
rect 1863 1680 1864 1681
rect 1897 1680 1898 1681
rect 1878 1682 1879 1683
rect 1915 1682 1916 1683
rect 1881 1684 1882 1685
rect 1888 1684 1889 1685
rect 1884 1686 1885 1687
rect 1918 1686 1919 1687
rect 1887 1688 1888 1689
rect 1900 1688 1901 1689
rect 1894 1690 1895 1691
rect 1935 1690 1936 1691
rect 1910 1692 1911 1693
rect 1938 1692 1939 1693
rect 1912 1694 1913 1695
rect 1948 1694 1949 1695
rect 1941 1696 1942 1697
rect 1954 1696 1955 1697
rect 1969 1696 1970 1697
rect 1976 1696 1977 1697
rect 1711 1705 1712 1706
rect 1717 1705 1718 1706
rect 1720 1705 1721 1706
rect 1723 1705 1724 1706
rect 1759 1705 1760 1706
rect 1763 1705 1764 1706
rect 1834 1705 1835 1706
rect 1847 1705 1848 1706
rect 1837 1707 1838 1708
rect 1841 1707 1842 1708
rect 1857 1707 1858 1708
rect 1913 1707 1914 1708
rect 1863 1709 1864 1710
rect 1904 1709 1905 1710
rect 1872 1711 1873 1712
rect 1884 1711 1885 1712
rect 1875 1713 1876 1714
rect 1887 1713 1888 1714
rect 1878 1715 1879 1716
rect 1907 1715 1908 1716
rect 1878 1717 1879 1718
rect 1900 1717 1901 1718
rect 1904 1717 1905 1718
rect 1910 1717 1911 1718
rect 1916 1717 1917 1718
rect 1937 1717 1938 1718
rect 1711 1726 1712 1727
rect 1717 1726 1718 1727
rect 1720 1726 1721 1727
rect 1749 1726 1750 1727
rect 1770 1726 1771 1727
rect 1784 1726 1785 1727
rect 1804 1726 1805 1727
rect 1831 1726 1832 1727
rect 1780 1728 1781 1729
rect 1804 1728 1805 1729
rect 1780 1730 1781 1731
rect 1791 1730 1792 1731
rect 1831 1730 1832 1731
rect 1881 1730 1882 1731
rect 1834 1732 1835 1733
rect 1843 1732 1844 1733
rect 1834 1734 1835 1735
rect 1840 1734 1841 1735
rect 1837 1736 1838 1737
rect 1907 1736 1908 1737
rect 1847 1738 1848 1739
rect 1857 1738 1858 1739
rect 1863 1738 1864 1739
rect 1872 1738 1873 1739
rect 1866 1740 1867 1741
rect 1875 1740 1876 1741
rect 1869 1742 1870 1743
rect 1878 1742 1879 1743
rect 1892 1742 1893 1743
rect 1904 1742 1905 1743
rect 1681 1751 1682 1752
rect 1688 1751 1689 1752
rect 1780 1751 1781 1752
rect 1784 1751 1785 1752
rect 1801 1751 1802 1752
rect 1804 1751 1805 1752
rect 1827 1751 1828 1752
rect 1831 1751 1832 1752
rect 1834 1751 1835 1752
rect 1836 1751 1837 1752
rect 1869 1751 1870 1752
rect 1871 1751 1872 1752
rect 1866 1753 1867 1754
rect 1868 1753 1869 1754
rect 1863 1755 1864 1756
rect 1865 1755 1866 1756
rect 1892 1755 1893 1756
rect 1898 1755 1899 1756
rect 1714 1782 1715 1783
rect 1868 1782 1869 1783
rect 1801 1784 1802 1785
rect 1811 1784 1812 1785
rect 1810 1786 1811 1787
rect 1827 1786 1828 1787
rect 1819 1788 1820 1789
rect 1836 1788 1837 1789
rect 1837 1790 1838 1791
rect 1865 1790 1866 1791
rect 1840 1792 1841 1793
rect 1871 1792 1872 1793
rect 1714 1801 1715 1802
rect 1718 1801 1719 1802
rect 1762 1801 1763 1802
rect 1840 1801 1841 1802
rect 1774 1803 1775 1804
rect 1801 1803 1802 1804
rect 1795 1805 1796 1806
rect 1837 1805 1838 1806
rect 1810 1807 1811 1808
rect 1813 1807 1814 1808
rect 1819 1807 1820 1808
rect 1822 1807 1823 1808
<< end >>
