magic
tech scmos
timestamp 1395743121
<< m1p >>
use CELL  1
transform -1 0 3179 0 1 2132
box 0 0 6 6
use CELL  2
transform -1 0 3114 0 1 1818
box 0 0 6 6
use CELL  3
transform -1 0 2619 0 1 5265
box 0 0 6 6
use CELL  4
transform -1 0 3264 0 1 3348
box 0 0 6 6
use CELL  5
transform 1 0 3112 0 -1 5078
box 0 0 6 6
use CELL  6
transform -1 0 2764 0 1 2663
box 0 0 6 6
use CELL  7
transform -1 0 2724 0 1 3543
box 0 0 6 6
use CELL  8
transform -1 0 2814 0 1 4421
box 0 0 6 6
use CELL  9
transform -1 0 2580 0 1 1818
box 0 0 6 6
use CELL  10
transform -1 0 2661 0 1 4666
box 0 0 6 6
use CELL  11
transform -1 0 2676 0 1 5442
box 0 0 6 6
use CELL  12
transform -1 0 3396 0 1 3107
box 0 0 6 6
use CELL  13
transform -1 0 2562 0 1 4212
box 0 0 6 6
use CELL  14
transform -1 0 2568 0 1 5442
box 0 0 6 6
use CELL  15
transform -1 0 3152 0 1 1967
box 0 0 6 6
use CELL  16
transform -1 0 2712 0 1 5265
box 0 0 6 6
use CELL  17
transform -1 0 3397 0 1 2876
box 0 0 6 6
use CELL  18
transform -1 0 2607 0 1 3543
box 0 0 6 6
use CELL  19
transform -1 0 2599 0 1 4421
box 0 0 6 6
use CELL  20
transform 1 0 2781 0 -1 1483
box 0 0 6 6
use CELL  21
transform 1 0 3107 0 1 2132
box 0 0 6 6
use CELL  22
transform -1 0 2654 0 1 1477
box 0 0 6 6
use CELL  23
transform -1 0 2986 0 1 5265
box 0 0 6 6
use CELL  24
transform -1 0 2718 0 -1 4893
box 0 0 6 6
use CELL  25
transform 1 0 2637 0 -1 3354
box 0 0 6 6
use CELL  26
transform 1 0 2568 0 1 5265
box 0 0 6 6
use CELL  27
transform -1 0 3196 0 1 2876
box 0 0 6 6
use CELL  28
transform 1 0 2886 0 1 3543
box 0 0 6 6
use CELL  29
transform -1 0 3307 0 1 2876
box 0 0 6 6
use CELL  30
transform -1 0 3088 0 1 5265
box 0 0 6 6
use CELL  31
transform -1 0 2635 0 1 1331
box 0 0 6 6
use CELL  32
transform -1 0 3263 0 1 2876
box 0 0 6 6
use CELL  33
transform 1 0 3098 0 -1 5271
box 0 0 6 6
use CELL  34
transform 1 0 2551 0 1 4017
box 0 0 6 6
use CELL  35
transform 1 0 3101 0 1 1967
box 0 0 6 6
use CELL  36
transform 1 0 2592 0 1 5442
box 0 0 6 6
use CELL  37
transform -1 0 3151 0 1 5072
box 0 0 6 6
use CELL  38
transform -1 0 3257 0 1 3796
box 0 0 6 6
use CELL  39
transform -1 0 2626 0 1 4017
box 0 0 6 6
use CELL  40
transform 1 0 3044 0 1 1574
box 0 0 6 6
use CELL  41
transform -1 0 3277 0 1 2876
box 0 0 6 6
use CELL  42
transform 1 0 3091 0 1 5265
box 0 0 6 6
use CELL  43
transform -1 0 2586 0 1 2876
box 0 0 6 6
use CELL  44
transform -1 0 2982 0 1 1574
box 0 0 6 6
use CELL  45
transform 1 0 2650 0 -1 2669
box 0 0 6 6
use CELL  46
transform -1 0 2833 0 1 1574
box 0 0 6 6
use CELL  47
transform 1 0 3232 0 1 2293
box 0 0 6 6
use CELL  48
transform -1 0 2608 0 1 4887
box 0 0 6 6
use CELL  49
transform 1 0 3113 0 1 5265
box 0 0 6 6
use CELL  50
transform -1 0 3153 0 1 2293
box 0 0 6 6
use CELL  51
transform -1 0 3057 0 -1 5271
box 0 0 6 6
use CELL  52
transform 1 0 2575 0 -1 5078
box 0 0 6 6
use CELL  53
transform 1 0 2960 0 1 1967
box 0 0 6 6
use CELL  54
transform -1 0 3299 0 1 3796
box 0 0 6 6
use CELL  55
transform -1 0 2688 0 1 1967
box 0 0 6 6
use CELL  56
transform 1 0 2663 0 -1 1685
box 0 0 6 6
use CELL  57
transform -1 0 2669 0 1 5442
box 0 0 6 6
use CELL  58
transform -1 0 2987 0 1 2132
box 0 0 6 6
use CELL  59
transform 1 0 2638 0 -1 1973
box 0 0 6 6
use CELL  60
transform 1 0 3185 0 1 5072
box 0 0 6 6
use CELL  61
transform -1 0 3143 0 1 2132
box 0 0 6 6
use CELL  62
transform -1 0 3243 0 1 4421
box 0 0 6 6
use CELL  63
transform -1 0 2690 0 -1 5078
box 0 0 6 6
use CELL  64
transform 1 0 3284 0 1 3348
box 0 0 6 6
use CELL  65
transform -1 0 3064 0 1 2462
box 0 0 6 6
use CELL  66
transform 1 0 3384 0 -1 2882
box 0 0 6 6
use CELL  67
transform -1 0 2685 0 1 5442
box 0 0 6 6
use CELL  68
transform 1 0 3071 0 1 5442
box 0 0 6 6
use CELL  69
transform -1 0 2580 0 1 3107
box 0 0 6 6
use CELL  70
transform -1 0 2592 0 1 2132
box 0 0 6 6
use CELL  71
transform -1 0 3317 0 1 4421
box 0 0 6 6
use CELL  72
transform 1 0 2634 0 -1 5271
box 0 0 6 6
use CELL  73
transform 1 0 2667 0 1 2132
box 0 0 6 6
use CELL  74
transform -1 0 2773 0 1 1574
box 0 0 6 6
use CELL  75
transform -1 0 2658 0 1 4017
box 0 0 6 6
use CELL  76
transform -1 0 3304 0 1 4017
box 0 0 6 6
use CELL  77
transform 1 0 2986 0 1 1679
box 0 0 6 6
use CELL  78
transform -1 0 3046 0 1 4017
box 0 0 6 6
use CELL  79
transform -1 0 3002 0 -1 4672
box 0 0 6 6
use CELL  80
transform 1 0 2545 0 -1 3113
box 0 0 6 6
use CELL  81
transform -1 0 2685 0 -1 1337
box 0 0 6 6
use CELL  82
transform -1 0 3044 0 1 1967
box 0 0 6 6
use CELL  83
transform -1 0 2737 0 1 2132
box 0 0 6 6
use CELL  84
transform -1 0 2569 0 1 4212
box 0 0 6 6
use CELL  85
transform -1 0 2593 0 1 3543
box 0 0 6 6
use CELL  86
transform -1 0 2592 0 1 1818
box 0 0 6 6
use CELL  87
transform -1 0 3292 0 -1 3802
box 0 0 6 6
use CELL  88
transform -1 0 2615 0 1 4887
box 0 0 6 6
use CELL  89
transform -1 0 2617 0 1 4212
box 0 0 6 6
use CELL  90
transform 1 0 3092 0 1 1818
box 0 0 6 6
use CELL  91
transform 1 0 2655 0 1 1384
box 0 0 6 6
use CELL  92
transform -1 0 2933 0 1 2132
box 0 0 6 6
use CELL  93
transform -1 0 2638 0 1 2132
box 0 0 6 6
use CELL  94
transform -1 0 2601 0 -1 1390
box 0 0 6 6
use CELL  95
transform -1 0 2676 0 1 5265
box 0 0 6 6
use CELL  96
transform -1 0 2617 0 -1 2138
box 0 0 6 6
use CELL  97
transform -1 0 3337 0 1 4212
box 0 0 6 6
use CELL  98
transform -1 0 3324 0 1 3107
box 0 0 6 6
use CELL  99
transform 1 0 3233 0 1 4017
box 0 0 6 6
use CELL  100
transform -1 0 3310 0 1 3543
box 0 0 6 6
use CELL  101
transform -1 0 2635 0 1 2293
box 0 0 6 6
use CELL  102
transform -1 0 2566 0 1 3796
box 0 0 6 6
use CELL  103
transform -1 0 2955 0 1 4212
box 0 0 6 6
use CELL  104
transform -1 0 3288 0 1 3107
box 0 0 6 6
use CELL  105
transform -1 0 3329 0 1 2663
box 0 0 6 6
use CELL  106
transform 1 0 3103 0 1 1679
box 0 0 6 6
use CELL  107
transform -1 0 2833 0 1 2663
box 0 0 6 6
use CELL  108
transform -1 0 3232 0 1 2462
box 0 0 6 6
use CELL  109
transform 1 0 3246 0 1 4887
box 0 0 6 6
use CELL  110
transform -1 0 2735 0 1 1818
box 0 0 6 6
use CELL  111
transform -1 0 2681 0 1 5599
box 0 0 6 6
use CELL  112
transform -1 0 3206 0 1 4666
box 0 0 6 6
use CELL  113
transform -1 0 2631 0 1 4212
box 0 0 6 6
use CELL  114
transform -1 0 2986 0 1 2462
box 0 0 6 6
use CELL  115
transform -1 0 2635 0 1 2876
box 0 0 6 6
use CELL  116
transform -1 0 2592 0 1 1384
box 0 0 6 6
use CELL  117
transform 1 0 3010 0 1 5599
box 0 0 6 6
use CELL  118
transform -1 0 2551 0 -1 1483
box 0 0 6 6
use CELL  119
transform -1 0 2591 0 1 4212
box 0 0 6 6
use CELL  120
transform -1 0 2621 0 1 2876
box 0 0 6 6
use CELL  121
transform 1 0 2977 0 1 5599
box 0 0 6 6
use CELL  122
transform -1 0 3205 0 1 2663
box 0 0 6 6
use CELL  123
transform -1 0 3206 0 1 2293
box 0 0 6 6
use CELL  124
transform -1 0 2992 0 1 4017
box 0 0 6 6
use CELL  125
transform -1 0 3194 0 1 4666
box 0 0 6 6
use CELL  126
transform -1 0 2606 0 1 2293
box 0 0 6 6
use CELL  127
transform 1 0 2615 0 1 4666
box 0 0 6 6
use CELL  128
transform 1 0 2891 0 1 1384
box 0 0 6 6
use CELL  129
transform 1 0 3160 0 -1 5271
box 0 0 6 6
use CELL  130
transform -1 0 3036 0 1 1818
box 0 0 6 6
use CELL  131
transform -1 0 2729 0 -1 5448
box 0 0 6 6
use CELL  132
transform -1 0 2586 0 1 3543
box 0 0 6 6
use CELL  133
transform -1 0 3136 0 1 4887
box 0 0 6 6
use CELL  134
transform -1 0 2624 0 1 2132
box 0 0 6 6
use CELL  135
transform 1 0 2984 0 1 5442
box 0 0 6 6
use CELL  136
transform -1 0 2737 0 1 1967
box 0 0 6 6
use CELL  137
transform -1 0 2672 0 1 3543
box 0 0 6 6
use CELL  138
transform -1 0 2634 0 1 5442
box 0 0 6 6
use CELL  139
transform -1 0 2649 0 -1 2669
box 0 0 6 6
use CELL  140
transform -1 0 2642 0 1 3107
box 0 0 6 6
use CELL  141
transform -1 0 3012 0 1 2293
box 0 0 6 6
use CELL  142
transform -1 0 2584 0 -1 4218
box 0 0 6 6
use CELL  143
transform -1 0 2712 0 -1 5783
box 0 0 6 6
use CELL  144
transform 1 0 2659 0 1 4017
box 0 0 6 6
use CELL  145
transform -1 0 3063 0 -1 5448
box 0 0 6 6
use CELL  146
transform -1 0 3271 0 1 4017
box 0 0 6 6
use CELL  147
transform -1 0 3383 0 1 2876
box 0 0 6 6
use CELL  148
transform 1 0 2813 0 1 1818
box 0 0 6 6
use CELL  149
transform -1 0 2719 0 1 5265
box 0 0 6 6
use CELL  150
transform -1 0 3345 0 -1 4427
box 0 0 6 6
use CELL  151
transform -1 0 3297 0 1 3348
box 0 0 6 6
use CELL  152
transform -1 0 2989 0 1 1574
box 0 0 6 6
use CELL  153
transform -1 0 2631 0 1 2132
box 0 0 6 6
use CELL  154
transform -1 0 2784 0 1 3543
box 0 0 6 6
use CELL  155
transform -1 0 2950 0 1 4017
box 0 0 6 6
use CELL  156
transform 1 0 3297 0 1 3543
box 0 0 6 6
use CELL  157
transform 1 0 3146 0 -1 5271
box 0 0 6 6
use CELL  158
transform -1 0 3318 0 1 4212
box 0 0 6 6
use CELL  159
transform 1 0 2607 0 1 4421
box 0 0 6 6
use CELL  160
transform -1 0 2699 0 1 4421
box 0 0 6 6
use CELL  161
transform -1 0 3121 0 -1 1824
box 0 0 6 6
use CELL  162
transform -1 0 2663 0 1 2462
box 0 0 6 6
use CELL  163
transform -1 0 3193 0 1 4212
box 0 0 6 6
use CELL  164
transform -1 0 2641 0 1 3543
box 0 0 6 6
use CELL  165
transform -1 0 2780 0 -1 1337
box 0 0 6 6
use CELL  166
transform -1 0 2647 0 1 5706
box 0 0 6 6
use CELL  167
transform 1 0 3078 0 1 5442
box 0 0 6 6
use CELL  168
transform -1 0 2787 0 1 2462
box 0 0 6 6
use CELL  169
transform 1 0 2607 0 -1 5448
box 0 0 6 6
use CELL  170
transform -1 0 2667 0 1 5599
box 0 0 6 6
use CELL  171
transform -1 0 2628 0 1 1574
box 0 0 6 6
use CELL  172
transform -1 0 3375 0 1 3543
box 0 0 6 6
use CELL  173
transform -1 0 2658 0 1 2293
box 0 0 6 6
use CELL  174
transform 1 0 3160 0 -1 1973
box 0 0 6 6
use CELL  175
transform 1 0 2781 0 1 5706
box 0 0 6 6
use CELL  176
transform 1 0 2610 0 -1 2468
box 0 0 6 6
use CELL  177
transform 1 0 2547 0 1 3796
box 0 0 6 6
use CELL  178
transform 1 0 2574 0 1 5706
box 0 0 6 6
use CELL  179
transform -1 0 2928 0 -1 5605
box 0 0 6 6
use CELL  180
transform -1 0 3223 0 1 4212
box 0 0 6 6
use CELL  181
transform -1 0 3078 0 1 3107
box 0 0 6 6
use CELL  182
transform -1 0 2851 0 1 2876
box 0 0 6 6
use CELL  183
transform -1 0 2654 0 1 4666
box 0 0 6 6
use CELL  184
transform -1 0 2660 0 1 3543
box 0 0 6 6
use CELL  185
transform -1 0 2803 0 1 5599
box 0 0 6 6
use CELL  186
transform -1 0 2980 0 1 5072
box 0 0 6 6
use CELL  187
transform -1 0 3159 0 1 1967
box 0 0 6 6
use CELL  188
transform -1 0 3319 0 1 2876
box 0 0 6 6
use CELL  189
transform -1 0 3213 0 1 3107
box 0 0 6 6
use CELL  190
transform -1 0 2811 0 1 5706
box 0 0 6 6
use CELL  191
transform 1 0 2532 0 -1 1824
box 0 0 6 6
use CELL  192
transform -1 0 3171 0 1 2293
box 0 0 6 6
use CELL  193
transform -1 0 2595 0 1 2462
box 0 0 6 6
use CELL  194
transform -1 0 2646 0 1 1280
box 0 0 6 6
use CELL  195
transform 1 0 3246 0 1 3348
box 0 0 6 6
use CELL  196
transform -1 0 2739 0 1 5777
box 0 0 6 6
use CELL  197
transform -1 0 2823 0 -1 5712
box 0 0 6 6
use CELL  198
transform 1 0 3266 0 1 2293
box 0 0 6 6
use CELL  199
transform -1 0 2607 0 1 4666
box 0 0 6 6
use CELL  200
transform 1 0 3311 0 -1 3802
box 0 0 6 6
use CELL  201
transform 1 0 2648 0 -1 5712
box 0 0 6 6
use CELL  202
transform 1 0 2632 0 1 3796
box 0 0 6 6
use CELL  203
transform -1 0 2707 0 1 2876
box 0 0 6 6
use CELL  204
transform -1 0 2669 0 1 3796
box 0 0 6 6
use CELL  205
transform -1 0 3218 0 1 2462
box 0 0 6 6
use CELL  206
transform -1 0 3264 0 1 3796
box 0 0 6 6
use CELL  207
transform -1 0 2587 0 -1 5605
box 0 0 6 6
use CELL  208
transform -1 0 3271 0 -1 2669
box 0 0 6 6
use CELL  209
transform -1 0 2575 0 1 5072
box 0 0 6 6
use CELL  210
transform -1 0 2896 0 1 5599
box 0 0 6 6
use CELL  211
transform 1 0 2932 0 1 1477
box 0 0 6 6
use CELL  212
transform 1 0 3325 0 1 3796
box 0 0 6 6
use CELL  213
transform 1 0 2616 0 -1 1390
box 0 0 6 6
use CELL  214
transform -1 0 3024 0 1 2293
box 0 0 6 6
use CELL  215
transform 1 0 2695 0 -1 1337
box 0 0 6 6
use CELL  216
transform 1 0 3313 0 -1 4672
box 0 0 6 6
use CELL  217
transform 1 0 2740 0 -1 4893
box 0 0 6 6
use CELL  218
transform -1 0 2601 0 1 4887
box 0 0 6 6
use CELL  219
transform 1 0 2969 0 1 1477
box 0 0 6 6
use CELL  220
transform -1 0 2544 0 1 4421
box 0 0 6 6
use CELL  221
transform -1 0 2730 0 1 2132
box 0 0 6 6
use CELL  222
transform -1 0 2592 0 1 3796
box 0 0 6 6
use CELL  223
transform -1 0 2725 0 1 4017
box 0 0 6 6
use CELL  224
transform 1 0 2540 0 -1 3802
box 0 0 6 6
use CELL  225
transform -1 0 2793 0 1 2293
box 0 0 6 6
use CELL  226
transform -1 0 2899 0 1 3543
box 0 0 6 6
use CELL  227
transform -1 0 3368 0 1 3543
box 0 0 6 6
use CELL  228
transform 1 0 2638 0 1 1574
box 0 0 6 6
use CELL  229
transform -1 0 3074 0 -1 1685
box 0 0 6 6
use CELL  230
transform -1 0 2644 0 -1 2468
box 0 0 6 6
use CELL  231
transform 1 0 2775 0 -1 5783
box 0 0 6 6
use CELL  232
transform 1 0 2614 0 -1 3802
box 0 0 6 6
use CELL  233
transform 1 0 3037 0 1 1574
box 0 0 6 6
use CELL  234
transform -1 0 2605 0 1 4212
box 0 0 6 6
use CELL  235
transform -1 0 3278 0 1 4017
box 0 0 6 6
use CELL  236
transform -1 0 2725 0 1 4887
box 0 0 6 6
use CELL  237
transform -1 0 3232 0 1 3543
box 0 0 6 6
use CELL  238
transform -1 0 3103 0 -1 5448
box 0 0 6 6
use CELL  239
transform -1 0 2709 0 1 3107
box 0 0 6 6
use CELL  240
transform -1 0 2877 0 1 3796
box 0 0 6 6
use CELL  241
transform -1 0 2764 0 1 3348
box 0 0 6 6
use CELL  242
transform -1 0 2657 0 1 3796
box 0 0 6 6
use CELL  243
transform 1 0 3346 0 -1 4672
box 0 0 6 6
use CELL  244
transform -1 0 2725 0 -1 5712
box 0 0 6 6
use CELL  245
transform 1 0 2785 0 1 1384
box 0 0 6 6
use CELL  246
transform -1 0 2694 0 1 1331
box 0 0 6 6
use CELL  247
transform 1 0 3238 0 1 5072
box 0 0 6 6
use CELL  248
transform 1 0 2636 0 1 4017
box 0 0 6 6
use CELL  249
transform 1 0 2669 0 -1 4427
box 0 0 6 6
use CELL  250
transform -1 0 3216 0 1 5072
box 0 0 6 6
use CELL  251
transform 1 0 2678 0 1 1679
box 0 0 6 6
use CELL  252
transform -1 0 3290 0 -1 4218
box 0 0 6 6
use CELL  253
transform -1 0 2660 0 1 1967
box 0 0 6 6
use CELL  254
transform 1 0 3330 0 -1 3113
box 0 0 6 6
use CELL  255
transform 1 0 3258 0 1 5072
box 0 0 6 6
use CELL  256
transform -1 0 3234 0 1 3348
box 0 0 6 6
use CELL  257
transform -1 0 3184 0 1 4887
box 0 0 6 6
use CELL  258
transform 1 0 2735 0 1 4421
box 0 0 6 6
use CELL  259
transform -1 0 2616 0 1 5072
box 0 0 6 6
use CELL  260
transform -1 0 3237 0 1 5072
box 0 0 6 6
use CELL  261
transform -1 0 2580 0 1 4887
box 0 0 6 6
use CELL  262
transform 1 0 3075 0 1 1679
box 0 0 6 6
use CELL  263
transform -1 0 3162 0 1 4212
box 0 0 6 6
use CELL  264
transform -1 0 2605 0 1 2663
box 0 0 6 6
use CELL  265
transform 1 0 2532 0 -1 1390
box 0 0 6 6
use CELL  266
transform 1 0 3330 0 1 3348
box 0 0 6 6
use CELL  267
transform 1 0 3144 0 1 4421
box 0 0 6 6
use CELL  268
transform -1 0 2586 0 1 2462
box 0 0 6 6
use CELL  269
transform -1 0 2810 0 1 1331
box 0 0 6 6
use CELL  270
transform -1 0 2755 0 1 2663
box 0 0 6 6
use CELL  271
transform -1 0 2672 0 1 5777
box 0 0 6 6
use CELL  272
transform -1 0 2653 0 1 3543
box 0 0 6 6
use CELL  273
transform -1 0 2616 0 1 3107
box 0 0 6 6
use CELL  274
transform -1 0 2684 0 1 5777
box 0 0 6 6
use CELL  275
transform -1 0 2610 0 -1 1483
box 0 0 6 6
use CELL  276
transform 1 0 3166 0 -1 4023
box 0 0 6 6
use CELL  277
transform -1 0 2864 0 -1 5712
box 0 0 6 6
use CELL  278
transform 1 0 3082 0 1 1679
box 0 0 6 6
use CELL  279
transform -1 0 2772 0 1 3796
box 0 0 6 6
use CELL  280
transform -1 0 2687 0 1 2462
box 0 0 6 6
use CELL  281
transform 1 0 3132 0 1 5265
box 0 0 6 6
use CELL  282
transform 1 0 2662 0 -1 5712
box 0 0 6 6
use CELL  283
transform -1 0 2985 0 1 1679
box 0 0 6 6
use CELL  284
transform 1 0 3173 0 1 1967
box 0 0 6 6
use CELL  285
transform -1 0 3192 0 1 4421
box 0 0 6 6
use CELL  286
transform -1 0 3308 0 1 2663
box 0 0 6 6
use CELL  287
transform -1 0 2610 0 1 1679
box 0 0 6 6
use CELL  288
transform -1 0 3317 0 1 3543
box 0 0 6 6
use CELL  289
transform -1 0 3104 0 1 2132
box 0 0 6 6
use CELL  290
transform 1 0 3085 0 -1 1973
box 0 0 6 6
use CELL  291
transform -1 0 2720 0 1 4212
box 0 0 6 6
use CELL  292
transform 1 0 3125 0 1 5265
box 0 0 6 6
use CELL  293
transform 1 0 3171 0 1 4887
box 0 0 6 6
use CELL  294
transform 1 0 3339 0 -1 4672
box 0 0 6 6
use CELL  295
transform 1 0 2618 0 1 5599
box 0 0 6 6
use CELL  296
transform 1 0 2602 0 1 3348
box 0 0 6 6
use CELL  297
transform 1 0 3164 0 1 4666
box 0 0 6 6
use CELL  298
transform -1 0 3243 0 -1 2669
box 0 0 6 6
use CELL  299
transform -1 0 2643 0 1 5442
box 0 0 6 6
use CELL  300
transform 1 0 3020 0 1 2132
box 0 0 6 6
use CELL  301
transform -1 0 3164 0 1 3348
box 0 0 6 6
use CELL  302
transform 1 0 3319 0 -1 4218
box 0 0 6 6
use CELL  303
transform -1 0 3259 0 1 4421
box 0 0 6 6
use CELL  304
transform 1 0 2972 0 1 1679
box 0 0 6 6
use CELL  305
transform 1 0 3291 0 1 4212
box 0 0 6 6
use CELL  306
transform 1 0 3221 0 1 3348
box 0 0 6 6
use CELL  307
transform -1 0 3157 0 1 3348
box 0 0 6 6
use CELL  308
transform -1 0 2659 0 -1 1824
box 0 0 6 6
use CELL  309
transform -1 0 3100 0 1 1967
box 0 0 6 6
use CELL  310
transform -1 0 2634 0 1 4421
box 0 0 6 6
use CELL  311
transform -1 0 3265 0 -1 2299
box 0 0 6 6
use CELL  312
transform -1 0 3322 0 -1 2669
box 0 0 6 6
use CELL  313
transform -1 0 2728 0 1 1818
box 0 0 6 6
use CELL  314
transform -1 0 2791 0 1 2876
box 0 0 6 6
use CELL  315
transform -1 0 2776 0 1 4017
box 0 0 6 6
use CELL  316
transform -1 0 2683 0 -1 4218
box 0 0 6 6
use CELL  317
transform -1 0 3344 0 1 2876
box 0 0 6 6
use CELL  318
transform 1 0 2629 0 1 1967
box 0 0 6 6
use CELL  319
transform -1 0 3292 0 1 4017
box 0 0 6 6
use CELL  320
transform 1 0 2763 0 -1 2299
box 0 0 6 6
use CELL  321
transform -1 0 3250 0 1 2462
box 0 0 6 6
use CELL  322
transform 1 0 2905 0 1 1574
box 0 0 6 6
use CELL  323
transform -1 0 2621 0 1 2663
box 0 0 6 6
use CELL  324
transform 1 0 2709 0 -1 5448
box 0 0 6 6
use CELL  325
transform -1 0 3057 0 1 1574
box 0 0 6 6
use CELL  326
transform -1 0 2643 0 1 1679
box 0 0 6 6
use CELL  327
transform -1 0 3145 0 1 4887
box 0 0 6 6
use CELL  328
transform -1 0 2681 0 -1 1973
box 0 0 6 6
use CELL  329
transform -1 0 2652 0 1 2132
box 0 0 6 6
use CELL  330
transform -1 0 2636 0 1 1679
box 0 0 6 6
use CELL  331
transform -1 0 2799 0 1 3796
box 0 0 6 6
use CELL  332
transform 1 0 2710 0 1 1384
box 0 0 6 6
use CELL  333
transform -1 0 2628 0 1 3107
box 0 0 6 6
use CELL  334
transform -1 0 2704 0 1 2663
box 0 0 6 6
use CELL  335
transform 1 0 3345 0 1 2876
box 0 0 6 6
use CELL  336
transform -1 0 2712 0 -1 3354
box 0 0 6 6
use CELL  337
transform -1 0 2796 0 1 1331
box 0 0 6 6
use CELL  338
transform -1 0 3043 0 -1 5271
box 0 0 6 6
use CELL  339
transform 1 0 2538 0 -1 3113
box 0 0 6 6
use CELL  340
transform -1 0 3073 0 1 1818
box 0 0 6 6
use CELL  341
transform 1 0 2982 0 1 2293
box 0 0 6 6
use CELL  342
transform 1 0 2741 0 1 1477
box 0 0 6 6
use CELL  343
transform -1 0 2667 0 1 1331
box 0 0 6 6
use CELL  344
transform -1 0 3285 0 1 3796
box 0 0 6 6
use CELL  345
transform 1 0 2778 0 1 3107
box 0 0 6 6
use CELL  346
transform -1 0 2613 0 -1 3802
box 0 0 6 6
use CELL  347
transform 1 0 2656 0 1 1679
box 0 0 6 6
use CELL  348
transform -1 0 2990 0 1 1967
box 0 0 6 6
use CELL  349
transform 1 0 3218 0 1 4887
box 0 0 6 6
use CELL  350
transform -1 0 2866 0 -1 1483
box 0 0 6 6
use CELL  351
transform -1 0 2557 0 -1 1824
box 0 0 6 6
use CELL  352
transform -1 0 2684 0 1 4887
box 0 0 6 6
use CELL  353
transform -1 0 3382 0 1 3543
box 0 0 6 6
use CELL  354
transform 1 0 2925 0 1 1477
box 0 0 6 6
use CELL  355
transform -1 0 3329 0 1 3543
box 0 0 6 6
use CELL  356
transform -1 0 3014 0 1 2132
box 0 0 6 6
use CELL  357
transform -1 0 3339 0 1 4666
box 0 0 6 6
use CELL  358
transform -1 0 2538 0 1 1477
box 0 0 6 6
use CELL  359
transform -1 0 3200 0 1 5072
box 0 0 6 6
use CELL  360
transform -1 0 3192 0 1 2293
box 0 0 6 6
use CELL  361
transform -1 0 2752 0 1 2876
box 0 0 6 6
use CELL  362
transform 1 0 2639 0 1 2132
box 0 0 6 6
use CELL  363
transform -1 0 2702 0 1 3107
box 0 0 6 6
use CELL  364
transform 1 0 2721 0 -1 1685
box 0 0 6 6
use CELL  365
transform 1 0 2738 0 1 1967
box 0 0 6 6
use CELL  366
transform 1 0 3019 0 1 5442
box 0 0 6 6
use CELL  367
transform -1 0 2683 0 1 5265
box 0 0 6 6
use CELL  368
transform 1 0 3026 0 1 5442
box 0 0 6 6
use CELL  369
transform 1 0 2710 0 1 1818
box 0 0 6 6
use CELL  370
transform -1 0 3236 0 1 2663
box 0 0 6 6
use CELL  371
transform 1 0 2629 0 1 1477
box 0 0 6 6
use CELL  372
transform 1 0 3064 0 1 5442
box 0 0 6 6
use CELL  373
transform 1 0 2608 0 1 1967
box 0 0 6 6
use CELL  374
transform -1 0 2635 0 1 2663
box 0 0 6 6
use CELL  375
transform -1 0 2601 0 1 3348
box 0 0 6 6
use CELL  376
transform -1 0 3298 0 1 4666
box 0 0 6 6
use CELL  377
transform 1 0 2689 0 -1 2669
box 0 0 6 6
use CELL  378
transform 1 0 3323 0 -1 3354
box 0 0 6 6
use CELL  379
transform -1 0 2906 0 1 1967
box 0 0 6 6
use CELL  380
transform -1 0 3018 0 -1 5448
box 0 0 6 6
use CELL  381
transform 1 0 3129 0 1 1818
box 0 0 6 6
use CELL  382
transform 1 0 3091 0 -1 3549
box 0 0 6 6
use CELL  383
transform -1 0 2685 0 1 4666
box 0 0 6 6
use CELL  384
transform -1 0 2658 0 -1 1580
box 0 0 6 6
use CELL  385
transform -1 0 2622 0 1 2293
box 0 0 6 6
use CELL  386
transform -1 0 2698 0 1 1574
box 0 0 6 6
use CELL  387
transform -1 0 3050 0 1 4666
box 0 0 6 6
use CELL  388
transform 1 0 2645 0 -1 1580
box 0 0 6 6
use CELL  389
transform -1 0 2772 0 1 5777
box 0 0 6 6
use CELL  390
transform -1 0 2702 0 -1 1390
box 0 0 6 6
use CELL  391
transform -1 0 2739 0 1 3543
box 0 0 6 6
use CELL  392
transform 1 0 3316 0 -1 3354
box 0 0 6 6
use CELL  393
transform -1 0 3301 0 1 2663
box 0 0 6 6
use CELL  394
transform 1 0 3318 0 1 4421
box 0 0 6 6
use CELL  395
transform -1 0 2903 0 1 5599
box 0 0 6 6
use CELL  396
transform -1 0 3101 0 1 2462
box 0 0 6 6
use CELL  397
transform -1 0 2732 0 -1 5712
box 0 0 6 6
use CELL  398
transform 1 0 3099 0 1 1818
box 0 0 6 6
use CELL  399
transform 1 0 3089 0 1 1679
box 0 0 6 6
use CELL  400
transform -1 0 2628 0 1 1477
box 0 0 6 6
use CELL  401
transform 1 0 2801 0 1 1384
box 0 0 6 6
use CELL  402
transform 1 0 2588 0 1 4887
box 0 0 6 6
use CELL  403
transform -1 0 2729 0 1 4421
box 0 0 6 6
use CELL  404
transform -1 0 3048 0 1 2293
box 0 0 6 6
use CELL  405
transform -1 0 2604 0 1 5599
box 0 0 6 6
use CELL  406
transform -1 0 2649 0 -1 4023
box 0 0 6 6
use CELL  407
transform -1 0 2961 0 1 1477
box 0 0 6 6
use CELL  408
transform 1 0 2808 0 1 1384
box 0 0 6 6
use CELL  409
transform 1 0 2842 0 1 1384
box 0 0 6 6
use CELL  410
transform 1 0 3214 0 -1 2299
box 0 0 6 6
use CELL  411
transform -1 0 2664 0 1 3348
box 0 0 6 6
use CELL  412
transform -1 0 2658 0 1 5810
box 0 0 6 6
use CELL  413
transform 1 0 2622 0 -1 1337
box 0 0 6 6
use CELL  414
transform -1 0 3250 0 1 4421
box 0 0 6 6
use CELL  415
transform -1 0 3271 0 -1 3802
box 0 0 6 6
use CELL  416
transform 1 0 2849 0 1 1384
box 0 0 6 6
use CELL  417
transform 1 0 2856 0 1 1384
box 0 0 6 6
use CELL  418
transform 1 0 2648 0 1 5265
box 0 0 6 6
use CELL  419
transform 1 0 2756 0 -1 2299
box 0 0 6 6
use CELL  420
transform 1 0 3096 0 1 1679
box 0 0 6 6
use CELL  421
transform -1 0 3144 0 1 4212
box 0 0 6 6
use CELL  422
transform -1 0 2656 0 1 2876
box 0 0 6 6
use CELL  423
transform 1 0 3252 0 -1 5078
box 0 0 6 6
use CELL  424
transform 1 0 2868 0 1 1384
box 0 0 6 6
use CELL  425
transform -1 0 3156 0 1 1818
box 0 0 6 6
use CELL  426
transform -1 0 3094 0 1 2462
box 0 0 6 6
use CELL  427
transform -1 0 2649 0 1 3107
box 0 0 6 6
use CELL  428
transform -1 0 3181 0 1 2663
box 0 0 6 6
use CELL  429
transform -1 0 2671 0 -1 1824
box 0 0 6 6
use CELL  430
transform 1 0 2884 0 1 1384
box 0 0 6 6
use CELL  431
transform 1 0 2533 0 1 3796
box 0 0 6 6
use CELL  432
transform 1 0 3312 0 1 4017
box 0 0 6 6
use CELL  433
transform 1 0 3143 0 1 1818
box 0 0 6 6
use CELL  434
transform -1 0 3350 0 1 3543
box 0 0 6 6
use CELL  435
transform -1 0 2631 0 1 5599
box 0 0 6 6
use CELL  436
transform -1 0 2853 0 1 3107
box 0 0 6 6
use CELL  437
transform -1 0 2730 0 1 4666
box 0 0 6 6
use CELL  438
transform 1 0 3128 0 1 2132
box 0 0 6 6
use CELL  439
transform 1 0 3277 0 1 3348
box 0 0 6 6
use CELL  440
transform -1 0 2624 0 1 1818
box 0 0 6 6
use CELL  441
transform 1 0 2711 0 1 5072
box 0 0 6 6
use CELL  442
transform -1 0 3284 0 1 4421
box 0 0 6 6
use CELL  443
transform -1 0 3121 0 1 4887
box 0 0 6 6
use CELL  444
transform -1 0 2967 0 1 4212
box 0 0 6 6
use CELL  445
transform -1 0 2771 0 1 5442
box 0 0 6 6
use CELL  446
transform 1 0 3227 0 1 3796
box 0 0 6 6
use CELL  447
transform 1 0 3272 0 1 2462
box 0 0 6 6
use CELL  448
transform -1 0 2786 0 -1 2138
box 0 0 6 6
use CELL  449
transform 1 0 2920 0 -1 1685
box 0 0 6 6
use CELL  450
transform -1 0 2739 0 1 3796
box 0 0 6 6
use CELL  451
transform -1 0 3011 0 1 5442
box 0 0 6 6
use CELL  452
transform 1 0 2684 0 1 4212
box 0 0 6 6
use CELL  453
transform 1 0 3403 0 1 3107
box 0 0 6 6
use CELL  454
transform -1 0 2665 0 -1 2299
box 0 0 6 6
use CELL  455
transform -1 0 2650 0 1 5442
box 0 0 6 6
use CELL  456
transform -1 0 2799 0 1 2462
box 0 0 6 6
use CELL  457
transform -1 0 2760 0 1 5777
box 0 0 6 6
use CELL  458
transform -1 0 2683 0 -1 1286
box 0 0 6 6
use CELL  459
transform -1 0 2661 0 -1 2138
box 0 0 6 6
use CELL  460
transform -1 0 2622 0 1 4887
box 0 0 6 6
use CELL  461
transform -1 0 3046 0 1 3796
box 0 0 6 6
use CELL  462
transform -1 0 2649 0 1 2876
box 0 0 6 6
use CELL  463
transform -1 0 2953 0 1 2876
box 0 0 6 6
use CELL  464
transform -1 0 2580 0 1 3348
box 0 0 6 6
use CELL  465
transform -1 0 3324 0 1 3796
box 0 0 6 6
use CELL  466
transform -1 0 2730 0 1 2462
box 0 0 6 6
use CELL  467
transform -1 0 2688 0 1 5599
box 0 0 6 6
use CELL  468
transform -1 0 3269 0 -1 4218
box 0 0 6 6
use CELL  469
transform 1 0 3337 0 1 3107
box 0 0 6 6
use CELL  470
transform 1 0 2707 0 1 2293
box 0 0 6 6
use CELL  471
transform -1 0 3186 0 1 4212
box 0 0 6 6
use CELL  472
transform -1 0 2679 0 1 3543
box 0 0 6 6
use CELL  473
transform 1 0 3270 0 1 4212
box 0 0 6 6
use CELL  474
transform 1 0 3122 0 1 1818
box 0 0 6 6
use CELL  475
transform 1 0 2894 0 1 1818
box 0 0 6 6
use CELL  476
transform -1 0 3333 0 1 4666
box 0 0 6 6
use CELL  477
transform 1 0 3383 0 -1 3113
box 0 0 6 6
use CELL  478
transform 1 0 2520 0 1 1384
box 0 0 6 6
use CELL  479
transform 1 0 3337 0 1 3543
box 0 0 6 6
use CELL  480
transform -1 0 2580 0 1 3796
box 0 0 6 6
use CELL  481
transform -1 0 2631 0 1 1384
box 0 0 6 6
use CELL  482
transform -1 0 2630 0 1 2462
box 0 0 6 6
use CELL  483
transform 1 0 3166 0 1 5072
box 0 0 6 6
use CELL  484
transform -1 0 2838 0 1 5706
box 0 0 6 6
use CELL  485
transform 1 0 3137 0 1 1967
box 0 0 6 6
use CELL  486
transform -1 0 2652 0 1 5599
box 0 0 6 6
use CELL  487
transform -1 0 2744 0 1 4666
box 0 0 6 6
use CELL  488
transform -1 0 2578 0 1 4212
box 0 0 6 6
use CELL  489
transform 1 0 2631 0 -1 5078
box 0 0 6 6
use CELL  490
transform -1 0 2853 0 -1 1337
box 0 0 6 6
use CELL  491
transform -1 0 2633 0 1 1818
box 0 0 6 6
use CELL  492
transform -1 0 3311 0 1 4212
box 0 0 6 6
use CELL  493
transform 1 0 2593 0 -1 2138
box 0 0 6 6
use CELL  494
transform 1 0 2996 0 -1 2138
box 0 0 6 6
use CELL  495
transform 1 0 3058 0 -1 2669
box 0 0 6 6
use CELL  496
transform 1 0 3258 0 -1 4023
box 0 0 6 6
use CELL  497
transform -1 0 2918 0 1 1574
box 0 0 6 6
use CELL  498
transform -1 0 2893 0 1 2462
box 0 0 6 6
use CELL  499
transform -1 0 3220 0 1 3107
box 0 0 6 6
use CELL  500
transform -1 0 2780 0 1 1477
box 0 0 6 6
use CELL  501
transform 1 0 2743 0 1 4017
box 0 0 6 6
use CELL  502
transform 1 0 2997 0 -1 1580
box 0 0 6 6
use CELL  503
transform 1 0 3023 0 1 5599
box 0 0 6 6
use CELL  504
transform -1 0 3252 0 1 2293
box 0 0 6 6
use CELL  505
transform 1 0 3217 0 1 5072
box 0 0 6 6
use CELL  506
transform -1 0 2771 0 1 5706
box 0 0 6 6
use CELL  507
transform -1 0 3196 0 1 4887
box 0 0 6 6
use CELL  508
transform -1 0 3217 0 1 4887
box 0 0 6 6
use CELL  509
transform 1 0 3306 0 -1 4672
box 0 0 6 6
use CELL  510
transform 1 0 3194 0 1 2132
box 0 0 6 6
use CELL  511
transform -1 0 3023 0 1 5599
box 0 0 6 6
use CELL  512
transform -1 0 3206 0 1 2132
box 0 0 6 6
use CELL  513
transform -1 0 2949 0 1 5599
box 0 0 6 6
use CELL  514
transform -1 0 3166 0 1 3796
box 0 0 6 6
use CELL  515
transform -1 0 2598 0 1 4212
box 0 0 6 6
use CELL  516
transform 1 0 3273 0 -1 2299
box 0 0 6 6
use CELL  517
transform 1 0 2791 0 1 1574
box 0 0 6 6
use CELL  518
transform 1 0 2643 0 1 2293
box 0 0 6 6
use CELL  519
transform -1 0 2593 0 1 4017
box 0 0 6 6
use CELL  520
transform -1 0 2647 0 1 4666
box 0 0 6 6
use CELL  521
transform 1 0 3279 0 -1 2468
box 0 0 6 6
use CELL  522
transform -1 0 2669 0 1 1967
box 0 0 6 6
use CELL  523
transform -1 0 2628 0 1 2876
box 0 0 6 6
use CELL  524
transform 1 0 3167 0 -1 2468
box 0 0 6 6
use CELL  525
transform -1 0 2935 0 1 5599
box 0 0 6 6
use CELL  526
transform -1 0 2638 0 1 4212
box 0 0 6 6
use CELL  527
transform -1 0 2594 0 -1 3354
box 0 0 6 6
use CELL  528
transform 1 0 2720 0 -1 1337
box 0 0 6 6
use CELL  529
transform -1 0 2645 0 1 1818
box 0 0 6 6
use CELL  530
transform -1 0 3179 0 1 5072
box 0 0 6 6
use CELL  531
transform -1 0 2627 0 1 4421
box 0 0 6 6
use CELL  532
transform -1 0 3292 0 1 2462
box 0 0 6 6
use CELL  533
transform -1 0 3283 0 1 2663
box 0 0 6 6
use CELL  534
transform -1 0 2532 0 1 3107
box 0 0 6 6
use CELL  535
transform -1 0 2676 0 1 5810
box 0 0 6 6
use CELL  536
transform 1 0 2919 0 1 1574
box 0 0 6 6
use CELL  537
transform -1 0 2731 0 1 5072
box 0 0 6 6
use CELL  538
transform 1 0 2562 0 -1 5078
box 0 0 6 6
use CELL  539
transform 1 0 3104 0 -1 5448
box 0 0 6 6
use CELL  540
transform -1 0 2623 0 1 2462
box 0 0 6 6
use CELL  541
transform 1 0 3258 0 1 2462
box 0 0 6 6
use CELL  542
transform 1 0 2990 0 1 1574
box 0 0 6 6
use CELL  543
transform 1 0 2685 0 1 1574
box 0 0 6 6
use CELL  544
transform 1 0 3078 0 1 1967
box 0 0 6 6
use CELL  545
transform -1 0 3170 0 1 4887
box 0 0 6 6
use CELL  546
transform -1 0 2592 0 -1 2299
box 0 0 6 6
use CELL  547
transform -1 0 2722 0 1 5442
box 0 0 6 6
use CELL  548
transform 1 0 3009 0 1 1574
box 0 0 6 6
use CELL  549
transform -1 0 2598 0 1 1967
box 0 0 6 6
use CELL  550
transform 1 0 2663 0 -1 5271
box 0 0 6 6
use CELL  551
transform -1 0 2886 0 -1 2468
box 0 0 6 6
use CELL  552
transform -1 0 2683 0 1 5072
box 0 0 6 6
use CELL  553
transform -1 0 2614 0 1 4017
box 0 0 6 6
use CELL  554
transform -1 0 2532 0 -1 1337
box 0 0 6 6
use CELL  555
transform -1 0 2614 0 1 4666
box 0 0 6 6
use CELL  556
transform 1 0 3016 0 1 1574
box 0 0 6 6
use CELL  557
transform -1 0 2628 0 1 2663
box 0 0 6 6
use CELL  558
transform -1 0 3273 0 1 4666
box 0 0 6 6
use CELL  559
transform 1 0 3023 0 1 1574
box 0 0 6 6
use CELL  560
transform -1 0 2808 0 1 3543
box 0 0 6 6
use CELL  561
transform 1 0 3030 0 1 1574
box 0 0 6 6
use CELL  562
transform 1 0 2611 0 -1 1824
box 0 0 6 6
use CELL  563
transform -1 0 3246 0 1 4017
box 0 0 6 6
use CELL  564
transform -1 0 2628 0 1 5265
box 0 0 6 6
use CELL  565
transform -1 0 2720 0 1 2293
box 0 0 6 6
use CELL  566
transform 1 0 2882 0 1 5706
box 0 0 6 6
use CELL  567
transform -1 0 2602 0 1 2462
box 0 0 6 6
use CELL  568
transform 1 0 2898 0 1 1384
box 0 0 6 6
use CELL  569
transform -1 0 3226 0 1 3796
box 0 0 6 6
use CELL  570
transform -1 0 2695 0 1 5599
box 0 0 6 6
use CELL  571
transform -1 0 2921 0 1 5599
box 0 0 6 6
use CELL  572
transform -1 0 3326 0 1 2876
box 0 0 6 6
use CELL  573
transform -1 0 2845 0 1 5706
box 0 0 6 6
use CELL  574
transform -1 0 2674 0 1 2663
box 0 0 6 6
use CELL  575
transform 1 0 3071 0 1 1967
box 0 0 6 6
use CELL  576
transform -1 0 2610 0 1 1818
box 0 0 6 6
use CELL  577
transform -1 0 2610 0 1 1331
box 0 0 6 6
use CELL  578
transform -1 0 2635 0 -1 1580
box 0 0 6 6
use CELL  579
transform -1 0 3039 0 -1 5448
box 0 0 6 6
use CELL  580
transform 1 0 2853 0 1 1477
box 0 0 6 6
use CELL  581
transform 1 0 3056 0 1 1679
box 0 0 6 6
use CELL  582
transform 1 0 3239 0 -1 2299
box 0 0 6 6
use CELL  583
transform -1 0 3205 0 1 4887
box 0 0 6 6
use CELL  584
transform -1 0 2627 0 1 5442
box 0 0 6 6
use CELL  585
transform -1 0 3225 0 1 2462
box 0 0 6 6
use CELL  586
transform -1 0 3237 0 1 4666
box 0 0 6 6
use CELL  587
transform -1 0 2718 0 1 5810
box 0 0 6 6
use CELL  588
transform 1 0 2773 0 1 1384
box 0 0 6 6
use CELL  589
transform -1 0 2839 0 1 2876
box 0 0 6 6
use CELL  590
transform 1 0 2692 0 -1 1286
box 0 0 6 6
use CELL  591
transform -1 0 3029 0 -1 1824
box 0 0 6 6
use CELL  592
transform -1 0 2876 0 1 5706
box 0 0 6 6
use CELL  593
transform 1 0 3207 0 -1 2299
box 0 0 6 6
use CELL  594
transform -1 0 2650 0 1 3796
box 0 0 6 6
use CELL  595
transform 1 0 3179 0 1 3348
box 0 0 6 6
use CELL  596
transform -1 0 2676 0 1 1574
box 0 0 6 6
use CELL  597
transform -1 0 3091 0 -1 1824
box 0 0 6 6
use CELL  598
transform -1 0 2737 0 1 4666
box 0 0 6 6
use CELL  599
transform 1 0 2641 0 1 4887
box 0 0 6 6
use CELL  600
transform -1 0 2972 0 1 1818
box 0 0 6 6
use CELL  601
transform -1 0 2588 0 1 5072
box 0 0 6 6
use CELL  602
transform -1 0 3066 0 1 1818
box 0 0 6 6
use CELL  603
transform -1 0 3264 0 1 2663
box 0 0 6 6
use CELL  604
transform -1 0 3197 0 1 3348
box 0 0 6 6
use CELL  605
transform -1 0 2607 0 1 4017
box 0 0 6 6
use CELL  606
transform 1 0 2703 0 -1 1390
box 0 0 6 6
use CELL  607
transform 1 0 2713 0 1 1331
box 0 0 6 6
use CELL  608
transform 1 0 3344 0 -1 3113
box 0 0 6 6
use CELL  609
transform 1 0 2669 0 -1 3113
box 0 0 6 6
use CELL  610
transform -1 0 3270 0 1 2876
box 0 0 6 6
use CELL  611
transform -1 0 2598 0 1 2663
box 0 0 6 6
use CELL  612
transform -1 0 2845 0 1 5599
box 0 0 6 6
use CELL  613
transform -1 0 2642 0 1 2876
box 0 0 6 6
use CELL  614
transform -1 0 3207 0 1 5072
box 0 0 6 6
use CELL  615
transform 1 0 2782 0 -1 5783
box 0 0 6 6
use CELL  616
transform 1 0 3272 0 1 3796
box 0 0 6 6
use CELL  617
transform -1 0 2767 0 1 5599
box 0 0 6 6
use CELL  618
transform -1 0 3064 0 1 3348
box 0 0 6 6
use CELL  619
transform 1 0 2574 0 -1 5605
box 0 0 6 6
use CELL  620
transform -1 0 2635 0 1 3107
box 0 0 6 6
use CELL  621
transform -1 0 2609 0 1 5072
box 0 0 6 6
use CELL  622
transform -1 0 3195 0 1 3107
box 0 0 6 6
use CELL  623
transform -1 0 2650 0 1 3348
box 0 0 6 6
use CELL  624
transform -1 0 2727 0 -1 4218
box 0 0 6 6
use CELL  625
transform -1 0 2724 0 1 5072
box 0 0 6 6
use CELL  626
transform -1 0 3193 0 1 2132
box 0 0 6 6
use CELL  627
transform -1 0 3145 0 1 5265
box 0 0 6 6
use CELL  628
transform -1 0 3336 0 1 3543
box 0 0 6 6
use CELL  629
transform -1 0 2647 0 1 5265
box 0 0 6 6
use CELL  630
transform 1 0 3299 0 1 4666
box 0 0 6 6
use CELL  631
transform -1 0 3283 0 1 4212
box 0 0 6 6
use CELL  632
transform -1 0 2931 0 1 4421
box 0 0 6 6
use CELL  633
transform -1 0 3161 0 1 2462
box 0 0 6 6
use CELL  634
transform -1 0 3081 0 1 5265
box 0 0 6 6
use CELL  635
transform -1 0 3106 0 1 2663
box 0 0 6 6
use CELL  636
transform -1 0 3227 0 1 2876
box 0 0 6 6
use CELL  637
transform -1 0 3271 0 1 2462
box 0 0 6 6
use CELL  638
transform 1 0 3031 0 1 1679
box 0 0 6 6
use CELL  639
transform -1 0 3296 0 1 3543
box 0 0 6 6
use CELL  640
transform -1 0 2600 0 -1 4023
box 0 0 6 6
use CELL  641
transform -1 0 2600 0 1 4666
box 0 0 6 6
use CELL  642
transform 1 0 3320 0 -1 4672
box 0 0 6 6
use CELL  643
transform 1 0 3298 0 -1 4218
box 0 0 6 6
use CELL  644
transform 1 0 2580 0 -1 4672
box 0 0 6 6
use CELL  645
transform -1 0 2788 0 1 3348
box 0 0 6 6
use CELL  646
transform -1 0 3227 0 1 3107
box 0 0 6 6
use CELL  647
transform 1 0 3157 0 1 4017
box 0 0 6 6
use CELL  648
transform 1 0 2622 0 1 1967
box 0 0 6 6
use CELL  649
transform -1 0 2654 0 1 4887
box 0 0 6 6
use CELL  650
transform -1 0 3160 0 1 5072
box 0 0 6 6
use CELL  651
transform -1 0 2606 0 1 3796
box 0 0 6 6
use CELL  652
transform -1 0 2762 0 -1 5712
box 0 0 6 6
use CELL  653
transform -1 0 2593 0 1 2876
box 0 0 6 6
use CELL  654
transform -1 0 2595 0 1 5072
box 0 0 6 6
use CELL  655
transform -1 0 2676 0 1 3796
box 0 0 6 6
use CELL  656
transform -1 0 2642 0 1 2663
box 0 0 6 6
use CELL  657
transform 1 0 3049 0 1 1679
box 0 0 6 6
use CELL  658
transform -1 0 2660 0 1 5777
box 0 0 6 6
use CELL  659
transform -1 0 2676 0 1 1280
box 0 0 6 6
use CELL  660
transform 1 0 2637 0 1 5599
box 0 0 6 6
use CELL  661
transform -1 0 2586 0 1 4017
box 0 0 6 6
use CELL  662
transform 1 0 3309 0 1 2663
box 0 0 6 6
use CELL  663
transform -1 0 2879 0 1 5442
box 0 0 6 6
use CELL  664
transform -1 0 2903 0 1 4666
box 0 0 6 6
use CELL  665
transform -1 0 2877 0 1 2293
box 0 0 6 6
use CELL  666
transform -1 0 3193 0 1 3543
box 0 0 6 6
use CELL  667
transform -1 0 2637 0 1 2462
box 0 0 6 6
use CELL  668
transform -1 0 2618 0 -1 5712
box 0 0 6 6
use CELL  669
transform 1 0 3245 0 1 5072
box 0 0 6 6
use CELL  670
transform 1 0 2976 0 1 1477
box 0 0 6 6
use CELL  671
transform 1 0 3271 0 1 4421
box 0 0 6 6
use CELL  672
transform -1 0 3142 0 1 5072
box 0 0 6 6
use CELL  673
transform 1 0 2877 0 1 1384
box 0 0 6 6
use CELL  674
transform 1 0 3011 0 -1 1973
box 0 0 6 6
use CELL  675
transform -1 0 2652 0 1 1818
box 0 0 6 6
use CELL  676
transform -1 0 2780 0 1 5706
box 0 0 6 6
use CELL  677
transform -1 0 2614 0 -1 2669
box 0 0 6 6
use CELL  678
transform -1 0 3208 0 1 2876
box 0 0 6 6
use CELL  679
transform -1 0 3212 0 1 2663
box 0 0 6 6
use CELL  680
transform -1 0 2744 0 1 2132
box 0 0 6 6
use CELL  681
transform -1 0 3039 0 1 3796
box 0 0 6 6
use CELL  682
transform -1 0 2700 0 1 2876
box 0 0 6 6
use CELL  683
transform 1 0 2835 0 1 1384
box 0 0 6 6
use CELL  684
transform -1 0 2719 0 1 3348
box 0 0 6 6
use CELL  685
transform 1 0 3119 0 1 2462
box 0 0 6 6
use CELL  686
transform -1 0 2657 0 1 3348
box 0 0 6 6
use CELL  687
transform -1 0 3173 0 1 3796
box 0 0 6 6
use CELL  688
transform -1 0 2873 0 1 1477
box 0 0 6 6
use CELL  689
transform -1 0 3172 0 1 5265
box 0 0 6 6
use CELL  690
transform -1 0 2806 0 -1 3354
box 0 0 6 6
use CELL  691
transform -1 0 2959 0 -1 1685
box 0 0 6 6
use CELL  692
transform -1 0 2817 0 -1 1337
box 0 0 6 6
use CELL  693
transform 1 0 2918 0 1 1477
box 0 0 6 6
use CELL  694
transform -1 0 3127 0 1 2132
box 0 0 6 6
use CELL  695
transform 1 0 3146 0 1 4887
box 0 0 6 6
use CELL  696
transform 1 0 2991 0 1 5599
box 0 0 6 6
use CELL  697
transform -1 0 3120 0 -1 2138
box 0 0 6 6
use CELL  698
transform -1 0 3130 0 1 4017
box 0 0 6 6
use CELL  699
transform -1 0 2817 0 1 1679
box 0 0 6 6
use CELL  700
transform 1 0 3359 0 1 4421
box 0 0 6 6
use CELL  701
transform -1 0 3262 0 1 4212
box 0 0 6 6
use CELL  702
transform -1 0 3031 0 -1 5271
box 0 0 6 6
use CELL  703
transform -1 0 2612 0 -1 5271
box 0 0 6 6
use CELL  704
transform -1 0 3050 0 1 5265
box 0 0 6 6
use CELL  705
transform -1 0 2670 0 1 2876
box 0 0 6 6
use CELL  706
transform -1 0 2602 0 1 5072
box 0 0 6 6
use CELL  707
transform 1 0 2985 0 1 4212
box 0 0 6 6
use CELL  708
transform -1 0 3155 0 1 2132
box 0 0 6 6
use CELL  709
transform 1 0 3188 0 1 2462
box 0 0 6 6
use CELL  710
transform 1 0 2965 0 1 1679
box 0 0 6 6
use CELL  711
transform 1 0 2647 0 1 1331
box 0 0 6 6
use CELL  712
transform -1 0 2681 0 1 1477
box 0 0 6 6
use CELL  713
transform -1 0 2600 0 1 3543
box 0 0 6 6
use CELL  714
transform -1 0 2761 0 1 4017
box 0 0 6 6
use CELL  715
transform -1 0 2705 0 1 5265
box 0 0 6 6
use CELL  716
transform -1 0 3258 0 1 4666
box 0 0 6 6
use CELL  717
transform -1 0 3289 0 1 3543
box 0 0 6 6
use CELL  718
transform 1 0 3214 0 1 2876
box 0 0 6 6
use CELL  719
transform -1 0 2972 0 -1 5448
box 0 0 6 6
use CELL  720
transform 1 0 3332 0 1 4421
box 0 0 6 6
use CELL  721
transform -1 0 2617 0 1 1679
box 0 0 6 6
use CELL  722
transform -1 0 3312 0 1 3107
box 0 0 6 6
use CELL  723
transform -1 0 2587 0 1 4887
box 0 0 6 6
use CELL  724
transform -1 0 2896 0 -1 1580
box 0 0 6 6
use CELL  725
transform 1 0 3112 0 -1 3802
box 0 0 6 6
use CELL  726
transform -1 0 2688 0 1 3348
box 0 0 6 6
use CELL  727
transform 1 0 3060 0 -1 4427
box 0 0 6 6
use CELL  728
transform -1 0 2897 0 1 1477
box 0 0 6 6
use CELL  729
transform -1 0 2628 0 1 2293
box 0 0 6 6
use CELL  730
transform 1 0 3199 0 1 3543
box 0 0 6 6
use CELL  731
transform 1 0 2783 0 -1 1337
box 0 0 6 6
use CELL  732
transform -1 0 2649 0 1 5072
box 0 0 6 6
use CELL  733
transform -1 0 2604 0 1 5706
box 0 0 6 6
use CELL  734
transform -1 0 3315 0 -1 3354
box 0 0 6 6
use CELL  735
transform -1 0 2689 0 1 1818
box 0 0 6 6
use CELL  736
transform -1 0 2620 0 1 5442
box 0 0 6 6
use CELL  737
transform 1 0 2936 0 1 5599
box 0 0 6 6
use CELL  738
transform -1 0 2748 0 1 4421
box 0 0 6 6
use CELL  739
transform -1 0 2640 0 1 4887
box 0 0 6 6
use CELL  740
transform -1 0 2636 0 1 3348
box 0 0 6 6
use CELL  741
transform -1 0 2656 0 1 5072
box 0 0 6 6
use CELL  742
transform -1 0 2700 0 1 4887
box 0 0 6 6
use CELL  743
transform 1 0 2962 0 1 5599
box 0 0 6 6
use CELL  744
transform -1 0 3331 0 1 4421
box 0 0 6 6
use CELL  745
transform -1 0 2692 0 1 5706
box 0 0 6 6
use CELL  746
transform -1 0 2663 0 1 2876
box 0 0 6 6
use CELL  747
transform -1 0 2660 0 -1 1337
box 0 0 6 6
use CELL  748
transform 1 0 3352 0 1 4421
box 0 0 6 6
use CELL  749
transform -1 0 2656 0 1 2462
box 0 0 6 6
use CELL  750
transform 1 0 2797 0 -1 1337
box 0 0 6 6
use CELL  751
transform 1 0 2599 0 -1 5271
box 0 0 6 6
use CELL  752
transform -1 0 2804 0 1 2132
box 0 0 6 6
use CELL  753
transform 1 0 3225 0 1 4887
box 0 0 6 6
use CELL  754
transform -1 0 2648 0 1 4421
box 0 0 6 6
use CELL  755
transform -1 0 3276 0 1 3348
box 0 0 6 6
use CELL  756
transform 1 0 2687 0 1 1679
box 0 0 6 6
use CELL  757
transform -1 0 2710 0 -1 1580
box 0 0 6 6
use CELL  758
transform -1 0 3172 0 -1 1973
box 0 0 6 6
use CELL  759
transform 1 0 2616 0 -1 5783
box 0 0 6 6
use CELL  760
transform -1 0 2838 0 -1 1337
box 0 0 6 6
use CELL  761
transform -1 0 3331 0 1 4212
box 0 0 6 6
use CELL  762
transform -1 0 2902 0 -1 4893
box 0 0 6 6
use CELL  763
transform 1 0 2688 0 1 4666
box 0 0 6 6
use CELL  764
transform 1 0 2694 0 1 1679
box 0 0 6 6
use CELL  765
transform -1 0 3352 0 1 4421
box 0 0 6 6
use CELL  766
transform -1 0 2609 0 1 2462
box 0 0 6 6
use CELL  767
transform -1 0 2754 0 1 4212
box 0 0 6 6
use CELL  768
transform -1 0 3180 0 1 3796
box 0 0 6 6
use CELL  769
transform 1 0 2575 0 -1 5271
box 0 0 6 6
use CELL  770
transform 1 0 3376 0 -1 3113
box 0 0 6 6
use CELL  771
transform 1 0 2605 0 1 5599
box 0 0 6 6
use CELL  772
transform -1 0 2895 0 1 5706
box 0 0 6 6
use CELL  773
transform 1 0 2818 0 1 1679
box 0 0 6 6
use CELL  774
transform -1 0 2532 0 1 3796
box 0 0 6 6
use CELL  775
transform 1 0 2651 0 1 5442
box 0 0 6 6
use CELL  776
transform -1 0 2817 0 1 3543
box 0 0 6 6
use CELL  777
transform -1 0 2841 0 1 1477
box 0 0 6 6
use CELL  778
transform -1 0 3186 0 1 2132
box 0 0 6 6
use CELL  779
transform -1 0 3115 0 -1 1685
box 0 0 6 6
use CELL  780
transform 1 0 2644 0 1 1679
box 0 0 6 6
use CELL  781
transform -1 0 3234 0 1 3107
box 0 0 6 6
use CELL  782
transform -1 0 3096 0 1 5442
box 0 0 6 6
use CELL  783
transform -1 0 2575 0 1 5442
box 0 0 6 6
use CELL  784
transform -1 0 3073 0 1 4887
box 0 0 6 6
use CELL  785
transform -1 0 3285 0 1 4017
box 0 0 6 6
use CELL  786
transform -1 0 3302 0 -1 4427
box 0 0 6 6
use CELL  787
transform -1 0 3211 0 1 4212
box 0 0 6 6
use CELL  788
transform -1 0 2663 0 1 3107
box 0 0 6 6
use CELL  789
transform -1 0 2614 0 1 3543
box 0 0 6 6
use CELL  790
transform -1 0 2642 0 -1 1483
box 0 0 6 6
use CELL  791
transform -1 0 3208 0 -1 4023
box 0 0 6 6
use CELL  792
transform 1 0 3211 0 1 3543
box 0 0 6 6
use CELL  793
transform -1 0 2718 0 1 5777
box 0 0 6 6
use CELL  794
transform -1 0 2653 0 1 5777
box 0 0 6 6
use CELL  795
transform 1 0 2962 0 1 1477
box 0 0 6 6
use CELL  796
transform -1 0 2606 0 1 4421
box 0 0 6 6
use CELL  797
transform -1 0 3213 0 -1 2138
box 0 0 6 6
use CELL  798
transform 1 0 3076 0 1 1818
box 0 0 6 6
use CELL  799
transform -1 0 2881 0 1 2663
box 0 0 6 6
use CELL  800
transform -1 0 3219 0 1 4421
box 0 0 6 6
use CELL  801
transform 1 0 2948 0 1 1477
box 0 0 6 6
use CELL  802
transform 1 0 2594 0 -1 2882
box 0 0 6 6
use CELL  803
transform -1 0 2559 0 1 3796
box 0 0 6 6
use CELL  804
transform 1 0 2684 0 1 5265
box 0 0 6 6
use CELL  805
transform -1 0 2800 0 1 1384
box 0 0 6 6
use CELL  806
transform -1 0 2615 0 1 2293
box 0 0 6 6
use CELL  807
transform -1 0 2710 0 1 1280
box 0 0 6 6
use CELL  808
transform -1 0 3403 0 1 3107
box 0 0 6 6
use CELL  809
transform -1 0 3199 0 1 2293
box 0 0 6 6
use CELL  810
transform -1 0 2695 0 1 1967
box 0 0 6 6
use CELL  811
transform -1 0 2550 0 1 4017
box 0 0 6 6
use CELL  812
transform -1 0 2611 0 1 5706
box 0 0 6 6
use CELL  813
transform 1 0 2593 0 1 2293
box 0 0 6 6
use CELL  814
transform -1 0 2668 0 1 5072
box 0 0 6 6
use CELL  815
transform -1 0 2642 0 1 2293
box 0 0 6 6
use CELL  816
transform -1 0 3180 0 1 2293
box 0 0 6 6
use CELL  817
transform -1 0 2640 0 -1 5712
box 0 0 6 6
use CELL  818
transform 1 0 3224 0 1 4666
box 0 0 6 6
use CELL  819
transform 1 0 2655 0 1 5706
box 0 0 6 6
use CELL  820
transform 1 0 2682 0 1 1384
box 0 0 6 6
use CELL  821
transform -1 0 3159 0 1 5265
box 0 0 6 6
use CELL  822
transform -1 0 2593 0 1 4666
box 0 0 6 6
use CELL  823
transform -1 0 2765 0 1 1477
box 0 0 6 6
use CELL  824
transform -1 0 2640 0 1 4666
box 0 0 6 6
use CELL  825
transform 1 0 3239 0 1 4887
box 0 0 6 6
use CELL  826
transform -1 0 2912 0 1 1477
box 0 0 6 6
use CELL  827
transform 1 0 3226 0 1 4017
box 0 0 6 6
use CELL  828
transform -1 0 2663 0 1 4887
box 0 0 6 6
use CELL  829
transform -1 0 2624 0 1 1679
box 0 0 6 6
use CELL  830
transform 1 0 2668 0 1 5599
box 0 0 6 6
use CELL  831
transform 1 0 3181 0 1 3796
box 0 0 6 6
use CELL  832
transform 1 0 2644 0 -1 4218
box 0 0 6 6
use CELL  833
transform -1 0 2607 0 1 1967
box 0 0 6 6
use CELL  834
transform -1 0 3291 0 1 4666
box 0 0 6 6
use CELL  835
transform 1 0 3251 0 1 2462
box 0 0 6 6
use CELL  836
transform -1 0 2624 0 1 4212
box 0 0 6 6
use CELL  837
transform -1 0 3142 0 -1 1824
box 0 0 6 6
use CELL  838
transform 1 0 2729 0 1 1477
box 0 0 6 6
use CELL  839
transform -1 0 2723 0 1 2462
box 0 0 6 6
use CELL  840
transform -1 0 3357 0 1 3107
box 0 0 6 6
use CELL  841
transform -1 0 3375 0 1 3107
box 0 0 6 6
use CELL  842
transform 1 0 2941 0 -1 1483
box 0 0 6 6
use CELL  843
transform -1 0 2852 0 -1 5712
box 0 0 6 6
use CELL  844
transform -1 0 2550 0 -1 1824
box 0 0 6 6
use CELL  845
transform -1 0 3238 0 1 4887
box 0 0 6 6
use CELL  846
transform -1 0 3004 0 1 5442
box 0 0 6 6
use CELL  847
transform -1 0 2651 0 1 1967
box 0 0 6 6
use CELL  848
transform -1 0 2587 0 1 3348
box 0 0 6 6
use CELL  849
transform -1 0 2633 0 1 4017
box 0 0 6 6
use CELL  850
transform -1 0 2679 0 1 1384
box 0 0 6 6
use CELL  851
transform -1 0 2604 0 1 3107
box 0 0 6 6
use CELL  852
transform -1 0 3311 0 1 4017
box 0 0 6 6
use CELL  853
transform -1 0 3259 0 1 2293
box 0 0 6 6
use CELL  854
transform 1 0 3112 0 1 2663
box 0 0 6 6
use CELL  855
transform -1 0 2592 0 1 3107
box 0 0 6 6
use CELL  856
transform -1 0 2619 0 1 1477
box 0 0 6 6
use CELL  857
transform 1 0 2725 0 1 5599
box 0 0 6 6
use CELL  858
transform -1 0 2870 0 1 1967
box 0 0 6 6
use CELL  859
transform 1 0 2539 0 1 1477
box 0 0 6 6
use CELL  860
transform -1 0 2997 0 1 5442
box 0 0 6 6
use CELL  861
transform 1 0 2648 0 1 1384
box 0 0 6 6
use CELL  862
transform -1 0 3246 0 1 4666
box 0 0 6 6
use CELL  863
transform -1 0 3154 0 -1 4023
box 0 0 6 6
use CELL  864
transform -1 0 2691 0 1 4887
box 0 0 6 6
use CELL  865
transform -1 0 3372 0 1 4421
box 0 0 6 6
use CELL  866
transform -1 0 2723 0 1 1477
box 0 0 6 6
use CELL  867
transform 1 0 3252 0 -1 4893
box 0 0 6 6
use CELL  868
transform 1 0 2622 0 1 5810
box 0 0 6 6
use CELL  869
transform 1 0 2615 0 -1 1973
box 0 0 6 6
use CELL  870
transform -1 0 3010 0 -1 5605
box 0 0 6 6
use CELL  871
transform 1 0 2984 0 1 5599
box 0 0 6 6
use CELL  872
transform -1 0 3206 0 1 2462
box 0 0 6 6
use CELL  873
transform -1 0 2599 0 1 3796
box 0 0 6 6
use CELL  874
transform -1 0 2641 0 1 4421
box 0 0 6 6
use CELL  875
transform -1 0 2847 0 -1 1337
box 0 0 6 6
use CELL  876
transform -1 0 3125 0 -1 1973
box 0 0 6 6
use CELL  877
transform -1 0 2625 0 1 5072
box 0 0 6 6
use CELL  878
transform 1 0 2997 0 -1 5605
box 0 0 6 6
use CELL  879
transform -1 0 2633 0 1 4666
box 0 0 6 6
use CELL  880
transform 1 0 3045 0 1 5442
box 0 0 6 6
use CELL  881
transform -1 0 2620 0 1 4421
box 0 0 6 6
use CELL  882
transform -1 0 2608 0 1 2132
box 0 0 6 6
use CELL  883
transform -1 0 2615 0 1 3348
box 0 0 6 6
use CELL  884
transform -1 0 2598 0 1 5265
box 0 0 6 6
use CELL  885
transform 1 0 2950 0 1 5599
box 0 0 6 6
use CELL  886
transform 1 0 2905 0 1 1384
box 0 0 6 6
use CELL  887
transform -1 0 2592 0 1 4421
box 0 0 6 6
use CELL  888
transform 1 0 2699 0 1 5777
box 0 0 6 6
use CELL  889
transform 1 0 3224 0 1 5072
box 0 0 6 6
use CELL  890
transform -1 0 2902 0 1 3348
box 0 0 6 6
use CELL  891
transform -1 0 2656 0 -1 3113
box 0 0 6 6
use CELL  892
transform 1 0 2689 0 1 1384
box 0 0 6 6
use CELL  893
transform -1 0 2754 0 1 3107
box 0 0 6 6
use CELL  894
transform 1 0 2729 0 -1 1337
box 0 0 6 6
use CELL  895
transform 1 0 2639 0 1 1384
box 0 0 6 6
use CELL  896
transform -1 0 2646 0 1 5777
box 0 0 6 6
use CELL  897
transform -1 0 3369 0 1 2876
box 0 0 6 6
use CELL  898
transform 1 0 2632 0 1 1384
box 0 0 6 6
use CELL  899
transform -1 0 2617 0 1 5599
box 0 0 6 6
use CELL  900
transform 1 0 3370 0 -1 2882
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 3155 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 3062 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 3003 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 2938 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 2862 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 3105 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 3091 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 2619 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 2616 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 2782 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 3312 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 3289 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 3218 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 3182 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 3252 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 2932 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 2882 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 3052 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 3027 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 3049 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 2730 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 2718 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 2707 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 2888 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 2917 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 2929 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 2904 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 2885 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 2890 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 2869 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 2662 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 2847 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 2696 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 2704 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 2715 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 2834 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 2794 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 2896 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 2691 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 2569 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 2562 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 2575 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 3167 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 3226 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 3238 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 3289 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 3357 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 3363 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 3303 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 3356 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 3305 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 3292 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 3131 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 3170 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 3229 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 3241 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 3292 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 3360 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 3366 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 3306 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 3359 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 3308 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 2864 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 2710 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 2914 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 2854 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 2626 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 2856 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 2906 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 2830 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 2880 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 2893 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 2838 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 2902 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 2848 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 2893 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 2924 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 2915 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 2954 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 2961 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 2977 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 3019 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 3172 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 3090 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 3103 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 3145 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 3139 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 3073 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 2705 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 2663 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 2719 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 2793 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 2780 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 2824 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 3076 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 2863 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 3079 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 2962 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 3023 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 3078 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 3036 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 2902 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 2849 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 2791 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 2981 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 3033 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 2982 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 2977 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-109
transform 1 0 3024 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-110
transform 1 0 2992 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-111
transform 1 0 2953 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-112
transform 1 0 2973 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-113
transform 1 0 2821 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-114
transform 1 0 2853 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-115
transform 1 0 2844 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-116
transform 1 0 2857 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-117
transform 1 0 2841 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-118
transform 1 0 2973 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-119
transform 1 0 2918 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-120
transform 1 0 2851 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-121
transform 1 0 2857 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-122
transform 1 0 2857 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-123
transform 1 0 2813 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-124
transform 1 0 2752 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-125
transform 1 0 2697 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-126
transform 1 0 2688 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-127
transform 1 0 3171 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-128
transform 1 0 3127 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-129
transform 1 0 3163 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-130
transform 1 0 3145 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-131
transform 1 0 3097 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-132
transform 1 0 3048 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-133
transform 1 0 3057 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-134
transform 1 0 3052 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-135
transform 1 0 3315 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-136
transform 1 0 3292 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-137
transform 1 0 3221 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-138
transform 1 0 3185 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-139
transform 1 0 3171 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-140
transform 1 0 3069 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-141
transform 1 0 3072 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-142
transform 1 0 2644 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-143
transform 1 0 2641 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-144
transform 1 0 3233 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-145
transform 1 0 3236 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-146
transform 1 0 3151 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-147
transform 1 0 2634 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-148
transform 1 0 2631 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-149
transform 1 0 2845 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-150
transform 1 0 3088 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-151
transform 1 0 3079 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-152
transform 1 0 3041 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-153
transform 1 0 3090 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-154
transform 1 0 3054 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-155
transform 1 0 3118 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-156
transform 1 0 3151 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-157
transform 1 0 3181 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-158
transform 1 0 3145 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-159
transform 1 0 3214 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-160
transform 1 0 3217 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-161
transform 1 0 2740 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-162
transform 1 0 2724 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-163
transform 1 0 2677 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-164
transform 1 0 2829 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-165
transform 1 0 2868 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-166
transform 1 0 2894 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-167
transform 1 0 2666 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-168
transform 1 0 3276 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-169
transform 1 0 3215 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-170
transform 1 0 3271 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-171
transform 1 0 3196 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-172
transform 1 0 3190 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-173
transform 1 0 3160 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-174
transform 1 0 3152 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-175
transform 1 0 3209 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-176
transform 1 0 3225 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-177
transform 1 0 3199 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-178
transform 1 0 3193 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-179
transform 1 0 3187 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-180
transform 1 0 3274 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-181
transform 1 0 3218 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-182
transform 1 0 3279 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-183
transform 1 0 3239 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-184
transform 1 0 3181 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-185
transform 1 0 3161 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-186
transform 1 0 3159 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-187
transform 1 0 3104 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-188
transform 1 0 3044 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-189
transform 1 0 3082 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-190
transform 1 0 2764 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-191
transform 1 0 2606 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-192
transform 1 0 2604 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-193
transform 1 0 2667 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-194
transform 1 0 2682 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-195
transform 1 0 2970 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-196
transform 1 0 2973 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-197
transform 1 0 2944 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-198
transform 1 0 2922 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-199
transform 1 0 2805 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-200
transform 1 0 2749 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-201
transform 1 0 2756 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-202
transform 1 0 2637 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-203
transform 1 0 3141 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-204
transform 1 0 3080 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-205
transform 1 0 3144 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-206
transform 1 0 3083 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-207
transform 1 0 3105 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-208
transform 1 0 3125 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-209
transform 1 0 3245 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-210
transform 1 0 3252 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-211
transform 1 0 3248 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-212
transform 1 0 2873 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-213
transform 1 0 2867 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-214
transform 1 0 2857 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-215
transform 1 0 2800 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-216
transform 1 0 2795 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-217
transform 1 0 2745 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-218
transform 1 0 2755 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-219
transform 1 0 2764 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-220
transform 1 0 2681 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-221
transform 1 0 2948 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-222
transform 1 0 3014 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-223
transform 1 0 2926 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-224
transform 1 0 2884 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-225
transform 1 0 2820 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-226
transform 1 0 2652 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-227
transform 1 0 2649 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-228
transform 1 0 2675 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-229
transform 1 0 2818 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-230
transform 1 0 2818 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-231
transform 1 0 2820 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-232
transform 1 0 2887 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-233
transform 1 0 2938 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-234
transform 1 0 2910 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-235
transform 1 0 2929 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-236
transform 1 0 2928 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-237
transform 1 0 2955 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-238
transform 1 0 2822 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-239
transform 1 0 2911 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-240
transform 1 0 3022 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-241
transform 1 0 2973 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-242
transform 1 0 2966 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-243
transform 1 0 2951 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-244
transform 1 0 3017 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-245
transform 1 0 3025 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-246
transform 1 0 2970 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-247
transform 1 0 2963 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-248
transform 1 0 3332 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-249
transform 1 0 3271 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-250
transform 1 0 3206 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-251
transform 1 0 2738 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-252
transform 1 0 2785 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-253
transform 1 0 2809 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-254
transform 1 0 2818 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-255
transform 1 0 2804 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-256
transform 1 0 2793 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-257
transform 1 0 2764 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-258
transform 1 0 2794 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-259
transform 1 0 2809 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-260
transform 1 0 2810 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-261
transform 1 0 2802 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-262
transform 1 0 2805 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-263
transform 1 0 2815 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-264
transform 1 0 2690 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-265
transform 1 0 2608 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-266
transform 1 0 3250 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-267
transform 1 0 3244 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-268
transform 1 0 3237 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-269
transform 1 0 3247 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-270
transform 1 0 3211 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-271
transform 1 0 3208 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-272
transform 1 0 2890 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-273
transform 1 0 2887 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-274
transform 1 0 2860 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-275
transform 1 0 2900 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-276
transform 1 0 2909 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-277
transform 1 0 2942 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-278
transform 1 0 3295 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-279
transform 1 0 3233 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-280
transform 1 0 3317 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-281
transform 1 0 3264 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-282
transform 1 0 3324 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-283
transform 1 0 3307 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-284
transform 1 0 3252 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-285
transform 1 0 3076 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-286
transform 1 0 3142 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-287
transform 1 0 2685 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-288
transform 1 0 2679 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-289
transform 1 0 2771 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-290
transform 1 0 2824 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-291
transform 1 0 2875 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-292
transform 1 0 2855 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-293
transform 1 0 2885 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-294
transform 1 0 2924 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-295
transform 1 0 2931 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-296
transform 1 0 2932 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-297
transform 1 0 2992 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-298
transform 1 0 2904 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-299
transform 1 0 2938 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-300
transform 1 0 2968 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-301
transform 1 0 3016 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-302
transform 1 0 2991 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-303
transform 1 0 2974 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-304
transform 1 0 2633 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-305
transform 1 0 2748 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-306
transform 1 0 2742 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-307
transform 1 0 2752 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-308
transform 1 0 2742 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-309
transform 1 0 2708 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-310
transform 1 0 2664 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-311
transform 1 0 2663 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-312
transform 1 0 2624 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-313
transform 1 0 3220 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-314
transform 1 0 2866 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-315
transform 1 0 2685 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-316
transform 1 0 2949 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-317
transform 1 0 2910 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-318
transform 1 0 2681 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-319
transform 1 0 2671 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-320
transform 1 0 2687 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-321
transform 1 0 3073 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-322
transform 1 0 3028 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-323
transform 1 0 2967 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-324
transform 1 0 2918 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-325
transform 1 0 2948 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-326
transform 1 0 2898 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-327
transform 1 0 2891 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-328
transform 1 0 2680 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-329
transform 1 0 2847 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-330
transform 1 0 2815 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-331
transform 1 0 2917 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-332
transform 1 0 2836 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-333
transform 1 0 2963 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-334
transform 1 0 2985 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-335
transform 1 0 2958 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-336
transform 1 0 2746 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-337
transform 1 0 2764 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-338
transform 1 0 2767 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-339
transform 1 0 2765 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-340
transform 1 0 2775 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-341
transform 1 0 2766 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-342
transform 1 0 2953 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-343
transform 1 0 2752 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-344
transform 1 0 2770 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-345
transform 1 0 2773 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-346
transform 1 0 2789 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-347
transform 1 0 2787 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-348
transform 1 0 2772 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-349
transform 1 0 2782 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-350
transform 1 0 2997 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-351
transform 1 0 3264 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-352
transform 1 0 3258 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-353
transform 1 0 3256 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-354
transform 1 0 3259 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-355
transform 1 0 3255 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-356
transform 1 0 3238 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-357
transform 1 0 2686 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-358
transform 1 0 2706 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-359
transform 1 0 2641 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-360
transform 1 0 2997 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-361
transform 1 0 3326 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-362
transform 1 0 2929 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-363
transform 1 0 2935 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-364
transform 1 0 3175 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-365
transform 1 0 3173 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-366
transform 1 0 3224 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-367
transform 1 0 3277 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-368
transform 1 0 3288 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-369
transform 1 0 3240 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-370
transform 1 0 3277 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-371
transform 1 0 2891 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-372
transform 1 0 2846 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-373
transform 1 0 2845 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-374
transform 1 0 2849 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-375
transform 1 0 2677 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-376
transform 1 0 2693 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-377
transform 1 0 2674 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-378
transform 1 0 2735 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-379
transform 1 0 2782 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-380
transform 1 0 2806 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-381
transform 1 0 2815 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-382
transform 1 0 2843 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-383
transform 1 0 2814 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-384
transform 1 0 2853 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-385
transform 1 0 2938 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-386
transform 1 0 3021 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-387
transform 1 0 2733 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-388
transform 1 0 3049 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-389
transform 1 0 3112 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-390
transform 1 0 3174 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-391
transform 1 0 3130 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-392
transform 1 0 3166 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-393
transform 1 0 3148 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-394
transform 1 0 2908 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-395
transform 1 0 2926 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-396
transform 1 0 2676 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-397
transform 1 0 2910 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-398
transform 1 0 2827 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-399
transform 1 0 2769 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-400
transform 1 0 2557 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-401
transform 1 0 2550 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-402
transform 1 0 2550 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-403
transform 1 0 2592 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-404
transform 1 0 2598 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-405
transform 1 0 2599 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-406
transform 1 0 2606 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-407
transform 1 0 2586 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-408
transform 1 0 2605 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-409
transform 1 0 2612 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-410
transform 1 0 2607 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-411
transform 1 0 2615 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-412
transform 1 0 2632 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-413
transform 1 0 2638 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-414
transform 1 0 2649 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-415
transform 1 0 2650 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-416
transform 1 0 2666 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-417
transform 1 0 2661 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-418
transform 1 0 2654 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-419
transform 1 0 2640 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-420
transform 1 0 2628 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-421
transform 1 0 2604 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-422
transform 1 0 2565 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-423
transform 1 0 2705 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-424
transform 1 0 2689 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-425
transform 1 0 2904 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-426
transform 1 0 2676 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-427
transform 1 0 2691 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-428
transform 1 0 2697 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-429
transform 1 0 2911 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-430
transform 1 0 3153 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-431
transform 1 0 3028 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-432
transform 1 0 3106 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-433
transform 1 0 3067 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-434
transform 1 0 3046 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-435
transform 1 0 3031 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-436
transform 1 0 3109 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-437
transform 1 0 3070 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-438
transform 1 0 3040 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-439
transform 1 0 2934 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-440
transform 1 0 3109 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-441
transform 1 0 3106 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-442
transform 1 0 3031 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-443
transform 1 0 2978 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-444
transform 1 0 3140 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-445
transform 1 0 3072 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-446
transform 1 0 3114 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-447
transform 1 0 3143 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-448
transform 1 0 3112 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-449
transform 1 0 3109 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-450
transform 1 0 2733 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-451
transform 1 0 2773 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-452
transform 1 0 2725 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-453
transform 1 0 2763 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-454
transform 1 0 2727 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-455
transform 1 0 2737 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-456
transform 1 0 2721 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-457
transform 1 0 2709 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-458
transform 1 0 2694 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-459
transform 1 0 2681 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-460
transform 1 0 2685 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-461
transform 1 0 2680 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-462
transform 1 0 2877 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-463
transform 1 0 2665 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-464
transform 1 0 2867 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-465
transform 1 0 2831 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-466
transform 1 0 2804 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-467
transform 1 0 2684 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-468
transform 1 0 2661 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-469
transform 1 0 2642 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-470
transform 1 0 2622 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-471
transform 1 0 2874 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-472
transform 1 0 3207 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-473
transform 1 0 3205 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-474
transform 1 0 3279 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-475
transform 1 0 3308 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-476
transform 1 0 2870 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-477
transform 1 0 2806 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-478
transform 1 0 2753 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-479
transform 1 0 2685 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-480
transform 1 0 2701 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-481
transform 1 0 2892 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-482
transform 1 0 2961 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-483
transform 1 0 2709 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-484
transform 1 0 2691 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-485
transform 1 0 2674 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-486
transform 1 0 2660 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-487
transform 1 0 2679 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-488
transform 1 0 2664 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-489
transform 1 0 3082 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-490
transform 1 0 3091 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-491
transform 1 0 2998 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-492
transform 1 0 2921 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-493
transform 1 0 2836 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-494
transform 1 0 2694 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-495
transform 1 0 2685 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-496
transform 1 0 2691 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-497
transform 1 0 2894 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-498
transform 1 0 2949 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-499
transform 1 0 2932 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-500
transform 1 0 2881 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-501
transform 1 0 2875 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-502
transform 1 0 2746 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-503
transform 1 0 2825 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-504
transform 1 0 2758 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-505
transform 1 0 2758 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-506
transform 1 0 2886 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-507
transform 1 0 2920 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-508
transform 1 0 2848 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-509
transform 1 0 2736 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-510
transform 1 0 2839 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-511
transform 1 0 2871 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-512
transform 1 0 2868 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-513
transform 1 0 2899 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-514
transform 1 0 2898 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-515
transform 1 0 2916 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-516
transform 1 0 2870 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-517
transform 1 0 2875 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-518
transform 1 0 2752 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-519
transform 1 0 2734 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-520
transform 1 0 2703 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-521
transform 1 0 2729 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-522
transform 1 0 2706 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-523
transform 1 0 2738 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-524
transform 1 0 2779 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-525
transform 1 0 2834 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-526
transform 1 0 2956 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-527
transform 1 0 2864 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-528
transform 1 0 3214 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-529
transform 1 0 3211 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-530
transform 1 0 3243 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-531
transform 1 0 2899 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-532
transform 1 0 2935 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-533
transform 1 0 2890 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-534
transform 1 0 2840 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-535
transform 1 0 2785 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-536
transform 1 0 2744 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-537
transform 1 0 3258 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-538
transform 1 0 3184 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-539
transform 1 0 3179 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-540
transform 1 0 3107 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-541
transform 1 0 3051 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-542
transform 1 0 2971 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-543
transform 1 0 2876 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-544
transform 1 0 2788 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-545
transform 1 0 3243 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-546
transform 1 0 3280 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-547
transform 1 0 3193 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-548
transform 1 0 3223 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-549
transform 1 0 3229 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-550
transform 1 0 3265 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-551
transform 1 0 3291 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-552
transform 1 0 2873 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-553
transform 1 0 2814 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-554
transform 1 0 2813 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-555
transform 1 0 2892 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-556
transform 1 0 2811 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-557
transform 1 0 2713 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-558
transform 1 0 2718 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-559
transform 1 0 2701 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-560
transform 1 0 2693 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-561
transform 1 0 2737 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-562
transform 1 0 2740 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-563
transform 1 0 2998 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-564
transform 1 0 2929 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-565
transform 1 0 2979 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-566
transform 1 0 2856 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-567
transform 1 0 3003 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-568
transform 1 0 2971 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-569
transform 1 0 2976 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-570
transform 1 0 3051 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-571
transform 1 0 2874 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-572
transform 1 0 3000 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-573
transform 1 0 2866 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-574
transform 1 0 3039 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-575
transform 1 0 2820 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-576
transform 1 0 2850 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-577
transform 1 0 2837 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-578
transform 1 0 2797 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-579
transform 1 0 2835 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-580
transform 1 0 2841 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-581
transform 1 0 2831 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-582
transform 1 0 2742 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-583
transform 1 0 2747 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-584
transform 1 0 2768 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-585
transform 1 0 2757 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-586
transform 1 0 2872 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-587
transform 1 0 3117 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-588
transform 1 0 2766 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-589
transform 1 0 2740 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-590
transform 1 0 2718 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-591
transform 1 0 2759 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-592
transform 1 0 2752 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-593
transform 1 0 2808 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-594
transform 1 0 2818 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-595
transform 1 0 2911 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-596
transform 1 0 2707 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-597
transform 1 0 2750 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-598
transform 1 0 2770 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-599
transform 1 0 2776 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-600
transform 1 0 2791 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-601
transform 1 0 2831 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-602
transform 1 0 2844 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-603
transform 1 0 2704 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-604
transform 1 0 2747 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-605
transform 1 0 2793 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-606
transform 1 0 2903 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-607
transform 1 0 2771 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-608
transform 1 0 2713 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-609
transform 1 0 2704 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-610
transform 1 0 2770 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-611
transform 1 0 2710 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-612
transform 1 0 2660 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-613
transform 1 0 2781 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-614
transform 1 0 2768 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-615
transform 1 0 2780 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-616
transform 1 0 2750 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-617
transform 1 0 2706 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-618
transform 1 0 2698 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-619
transform 1 0 2701 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-620
transform 1 0 2676 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-621
transform 1 0 2715 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-622
transform 1 0 2704 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-623
transform 1 0 3262 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-624
transform 1 0 2880 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-625
transform 1 0 2885 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-626
transform 1 0 2861 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-627
transform 1 0 2837 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-628
transform 1 0 2769 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-629
transform 1 0 2734 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-630
transform 1 0 2902 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-631
transform 1 0 2950 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-632
transform 1 0 2791 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-633
transform 1 0 2799 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-634
transform 1 0 2905 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-635
transform 1 0 2775 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-636
transform 1 0 2775 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-637
transform 1 0 2803 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-638
transform 1 0 2803 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-639
transform 1 0 2835 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-640
transform 1 0 2863 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-641
transform 1 0 2962 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-642
transform 1 0 2994 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-643
transform 1 0 2842 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-644
transform 1 0 3125 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-645
transform 1 0 3143 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-646
transform 1 0 3180 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-647
transform 1 0 3209 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-648
transform 1 0 3274 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-649
transform 1 0 3335 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-650
transform 1 0 3294 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-651
transform 1 0 3234 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-652
transform 1 0 3265 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-653
transform 1 0 3211 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-654
transform 1 0 3217 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-655
transform 1 0 3250 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-656
transform 1 0 3302 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-657
transform 1 0 3273 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-658
transform 1 0 3196 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-659
transform 1 0 3191 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-660
transform 1 0 3119 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-661
transform 1 0 2881 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-662
transform 1 0 2981 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-663
transform 1 0 2886 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-664
transform 1 0 2676 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-665
transform 1 0 2618 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-666
transform 1 0 2643 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-667
transform 1 0 2676 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-668
transform 1 0 2722 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-669
transform 1 0 2734 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-670
transform 1 0 2706 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-671
transform 1 0 2786 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-672
transform 1 0 2829 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-673
transform 1 0 2787 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-674
transform 1 0 2797 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-675
transform 1 0 2778 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-676
transform 1 0 2793 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-677
transform 1 0 2703 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-678
transform 1 0 2687 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-679
transform 1 0 2682 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-680
transform 1 0 2686 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-681
transform 1 0 2678 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-682
transform 1 0 2692 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-683
transform 1 0 2703 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-684
transform 1 0 2660 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-685
transform 1 0 2659 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-686
transform 1 0 2675 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-687
transform 1 0 2635 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-688
transform 1 0 2610 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-689
transform 1 0 2592 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-690
transform 1 0 2909 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-691
transform 1 0 3180 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-692
transform 1 0 3146 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-693
transform 1 0 3097 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-694
transform 1 0 3094 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-695
transform 1 0 3126 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-696
transform 1 0 3183 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-697
transform 1 0 3073 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-698
transform 1 0 3010 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-699
transform 1 0 2974 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-700
transform 1 0 2919 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-701
transform 1 0 3001 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-702
transform 1 0 2971 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-703
transform 1 0 2907 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-704
transform 1 0 2906 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-705
transform 1 0 2876 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-706
transform 1 0 2903 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-707
transform 1 0 3049 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-708
transform 1 0 3024 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-709
transform 1 0 3022 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-710
transform 1 0 3007 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-711
transform 1 0 3058 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-712
transform 1 0 2819 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-713
transform 1 0 2838 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-714
transform 1 0 2790 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-715
transform 1 0 2817 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-716
transform 1 0 2788 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-717
transform 1 0 2784 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-718
transform 1 0 2767 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-719
transform 1 0 2776 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-720
transform 1 0 2821 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-721
transform 1 0 2909 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-722
transform 1 0 2959 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-723
transform 1 0 3022 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-724
transform 1 0 3031 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-725
transform 1 0 2920 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-726
transform 1 0 2926 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-727
transform 1 0 2993 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-728
transform 1 0 3021 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-729
transform 1 0 3009 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-730
transform 1 0 3010 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-731
transform 1 0 2932 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-732
transform 1 0 2896 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-733
transform 1 0 2855 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-734
transform 1 0 2929 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-735
transform 1 0 2990 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-736
transform 1 0 3018 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-737
transform 1 0 3006 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-738
transform 1 0 3113 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-739
transform 1 0 3116 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-740
transform 1 0 3134 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-741
transform 1 0 3234 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-742
transform 1 0 3164 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-743
transform 1 0 3205 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-744
transform 1 0 3193 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-745
transform 1 0 3149 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-746
transform 1 0 3135 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-747
transform 1 0 3092 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-748
transform 1 0 3065 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-749
transform 1 0 3054 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-750
transform 1 0 3019 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-751
transform 1 0 2952 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-752
transform 1 0 2885 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-753
transform 1 0 2829 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-754
transform 1 0 2823 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-755
transform 1 0 3196 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-756
transform 1 0 3152 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-757
transform 1 0 3138 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-758
transform 1 0 3095 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-759
transform 1 0 3068 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-760
transform 1 0 3057 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-761
transform 1 0 3022 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-762
transform 1 0 2955 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-763
transform 1 0 2888 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-764
transform 1 0 2832 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-765
transform 1 0 2826 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-766
transform 1 0 2736 0 1 1280
box 0 0 3 6
use FEEDTHRU  F-767
transform 1 0 3120 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-768
transform 1 0 3103 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-769
transform 1 0 3123 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-770
transform 1 0 3148 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-771
transform 1 0 3184 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-772
transform 1 0 2760 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-773
transform 1 0 2653 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-774
transform 1 0 2562 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-775
transform 1 0 2563 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-776
transform 1 0 3162 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-777
transform 1 0 3081 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-778
transform 1 0 3164 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-779
transform 1 0 3184 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-780
transform 1 0 3242 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-781
transform 1 0 3201 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-782
transform 1 0 3139 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-783
transform 1 0 3169 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-784
transform 1 0 2914 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-785
transform 1 0 2890 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-786
transform 1 0 2853 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-787
transform 1 0 2725 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-788
transform 1 0 2722 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-789
transform 1 0 2733 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-790
transform 1 0 2737 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-791
transform 1 0 2739 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-792
transform 1 0 2711 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-793
transform 1 0 2731 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-794
transform 1 0 2728 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-795
transform 1 0 2730 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-796
transform 1 0 2734 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-797
transform 1 0 2745 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-798
transform 1 0 2739 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-799
transform 1 0 2749 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-800
transform 1 0 2739 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-801
transform 1 0 2676 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-802
transform 1 0 2670 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-803
transform 1 0 2684 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-804
transform 1 0 2710 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-805
transform 1 0 2757 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-806
transform 1 0 2747 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-807
transform 1 0 2750 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-808
transform 1 0 2792 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-809
transform 1 0 2646 0 1 1280
box 0 0 3 6
use FEEDTHRU  F-810
transform 1 0 2673 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-811
transform 1 0 2667 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-812
transform 1 0 2702 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-813
transform 1 0 2716 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-814
transform 1 0 2763 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-815
transform 1 0 2718 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-816
transform 1 0 2924 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-817
transform 1 0 2777 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-818
transform 1 0 3196 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-819
transform 1 0 3223 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-820
transform 1 0 3259 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-821
transform 1 0 3261 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-822
transform 1 0 3187 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-823
transform 1 0 2811 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-824
transform 1 0 2968 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-825
transform 1 0 2851 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-826
transform 1 0 2907 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-827
transform 1 0 2832 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-828
transform 1 0 2830 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-829
transform 1 0 2805 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-830
transform 1 0 2815 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-831
transform 1 0 2815 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-832
transform 1 0 2895 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-833
transform 1 0 2838 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-834
transform 1 0 2845 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-835
transform 1 0 2817 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-836
transform 1 0 2889 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-837
transform 1 0 2836 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-838
transform 1 0 2811 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-839
transform 1 0 2859 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-840
transform 1 0 3131 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-841
transform 1 0 3111 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-842
transform 1 0 3136 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-843
transform 1 0 3154 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-844
transform 1 0 3137 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-845
transform 1 0 3156 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-846
transform 1 0 2702 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-847
transform 1 0 2696 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-848
transform 1 0 2685 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-849
transform 1 0 2884 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-850
transform 1 0 2939 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-851
transform 1 0 3034 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-852
transform 1 0 3070 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-853
transform 1 0 2863 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-854
transform 1 0 2933 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-855
transform 1 0 2986 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-856
transform 1 0 3055 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-857
transform 1 0 3046 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-858
transform 1 0 3050 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-859
transform 1 0 2851 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-860
transform 1 0 2645 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-861
transform 1 0 2711 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-862
transform 1 0 3052 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-863
transform 1 0 3088 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-864
transform 1 0 3148 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-865
transform 1 0 3132 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-866
transform 1 0 3076 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-867
transform 1 0 3103 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-868
transform 1 0 3100 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-869
transform 1 0 3079 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-870
transform 1 0 3102 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-871
transform 1 0 3120 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-872
transform 1 0 2710 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-873
transform 1 0 2707 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-874
transform 1 0 2914 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-875
transform 1 0 2749 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-876
transform 1 0 2740 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-877
transform 1 0 2748 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-878
transform 1 0 2699 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-879
transform 1 0 2710 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-880
transform 1 0 2694 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-881
transform 1 0 2715 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-882
transform 1 0 2700 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-883
transform 1 0 2693 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-884
transform 1 0 2691 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-885
transform 1 0 2695 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-886
transform 1 0 2669 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-887
transform 1 0 2668 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-888
transform 1 0 2679 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-889
transform 1 0 2635 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-890
transform 1 0 2633 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-891
transform 1 0 2789 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-892
transform 1 0 2819 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-893
transform 1 0 2824 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-894
transform 1 0 2902 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-895
transform 1 0 2901 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-896
transform 1 0 2886 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-897
transform 1 0 2861 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-898
transform 1 0 2833 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-899
transform 1 0 2812 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-900
transform 1 0 2812 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-901
transform 1 0 2816 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-902
transform 1 0 2767 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-903
transform 1 0 2920 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-904
transform 1 0 2937 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-905
transform 1 0 2898 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-906
transform 1 0 3025 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-907
transform 1 0 3217 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-908
transform 1 0 3185 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-909
transform 1 0 3246 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-910
transform 1 0 3245 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-911
transform 1 0 3065 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-912
transform 1 0 3006 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-913
transform 1 0 2896 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-914
transform 1 0 2896 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-915
transform 1 0 2811 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-916
transform 1 0 2991 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-917
transform 1 0 2798 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-918
transform 1 0 2916 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-919
transform 1 0 2788 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-920
transform 1 0 2781 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-921
transform 1 0 2784 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-922
transform 1 0 2767 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-923
transform 1 0 2760 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-924
transform 1 0 2800 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-925
transform 1 0 2787 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-926
transform 1 0 2796 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-927
transform 1 0 2776 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-928
transform 1 0 3193 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-929
transform 1 0 3231 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-930
transform 1 0 3215 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-931
transform 1 0 3127 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-932
transform 1 0 2911 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-933
transform 1 0 2914 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-934
transform 1 0 2846 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-935
transform 1 0 2939 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-936
transform 1 0 2994 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-937
transform 1 0 3106 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-938
transform 1 0 3079 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-939
transform 1 0 3135 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-940
transform 1 0 3151 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-941
transform 1 0 3091 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-942
transform 1 0 3055 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-943
transform 1 0 2994 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-944
transform 1 0 2987 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-945
transform 1 0 2954 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-946
transform 1 0 2951 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-947
transform 1 0 3087 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-948
transform 1 0 2980 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-949
transform 1 0 2988 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-950
transform 1 0 3016 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-951
transform 1 0 2991 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-952
transform 1 0 2983 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-953
transform 1 0 2935 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-954
transform 1 0 2946 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-955
transform 1 0 2886 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-956
transform 1 0 2860 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-957
transform 1 0 2844 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-958
transform 1 0 3142 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-959
transform 1 0 2823 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-960
transform 1 0 2844 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-961
transform 1 0 2812 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-962
transform 1 0 3103 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-963
transform 1 0 3194 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-964
transform 1 0 3201 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-965
transform 1 0 3162 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-966
transform 1 0 3142 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-967
transform 1 0 3168 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-968
transform 1 0 2765 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-969
transform 1 0 3104 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-970
transform 1 0 3082 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-971
transform 1 0 3115 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-972
transform 1 0 3212 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-973
transform 1 0 3228 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-974
transform 1 0 3202 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-975
transform 1 0 3112 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-976
transform 1 0 3070 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-977
transform 1 0 3118 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-978
transform 1 0 3097 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-979
transform 1 0 3156 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-980
transform 1 0 2940 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-981
transform 1 0 2967 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-982
transform 1 0 2956 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-983
transform 1 0 2946 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-984
transform 1 0 2941 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-985
transform 1 0 2950 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-986
transform 1 0 2779 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-987
transform 1 0 2825 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-988
transform 1 0 2865 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-989
transform 1 0 2826 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-990
transform 1 0 3130 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-991
transform 1 0 3133 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-992
transform 1 0 3121 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-993
transform 1 0 3206 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-994
transform 1 0 3268 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-995
transform 1 0 3232 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-996
transform 1 0 3118 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-997
transform 1 0 3063 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-998
transform 1 0 2731 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-999
transform 1 0 2719 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1000
transform 1 0 2783 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1001
transform 1 0 2826 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1002
transform 1 0 2784 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1003
transform 1 0 2794 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1004
transform 1 0 2775 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1005
transform 1 0 2790 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1006
transform 1 0 3042 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1007
transform 1 0 3029 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1008
transform 1 0 3034 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1009
transform 1 0 3051 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1010
transform 1 0 3054 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1011
transform 1 0 3026 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1012
transform 1 0 2989 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1013
transform 1 0 3025 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1014
transform 1 0 2902 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1015
transform 1 0 2766 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1016
transform 1 0 2770 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1017
transform 1 0 2779 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1018
transform 1 0 2772 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1019
transform 1 0 2794 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1020
transform 1 0 2826 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1021
transform 1 0 2805 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1022
transform 1 0 2830 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1023
transform 1 0 2730 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1024
transform 1 0 2732 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1025
transform 1 0 2744 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1026
transform 1 0 2713 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1027
transform 1 0 2541 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1028
transform 1 0 2560 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1029
transform 1 0 2559 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1030
transform 1 0 2650 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1031
transform 1 0 2636 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1032
transform 1 0 2651 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1033
transform 1 0 2682 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1034
transform 1 0 2671 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1035
transform 1 0 2672 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1036
transform 1 0 2704 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1037
transform 1 0 2713 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1038
transform 1 0 2709 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1039
transform 1 0 2725 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1040
transform 1 0 2757 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1041
transform 1 0 2763 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1042
transform 1 0 2761 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1043
transform 1 0 2745 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1044
transform 1 0 2799 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1045
transform 1 0 2756 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1046
transform 1 0 2709 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1047
transform 1 0 3237 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1048
transform 1 0 3297 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1049
transform 1 0 3251 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1050
transform 1 0 2755 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1051
transform 1 0 2761 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1052
transform 1 0 2791 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1053
transform 1 0 2847 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1054
transform 1 0 2899 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1055
transform 1 0 2959 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1056
transform 1 0 2957 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1057
transform 1 0 3043 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1058
transform 1 0 3018 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1059
transform 1 0 2992 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1060
transform 1 0 2980 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1061
transform 1 0 3046 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1062
transform 1 0 3021 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1063
transform 1 0 2947 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1064
transform 1 0 2667 0 1 5810
box 0 0 3 6
use FEEDTHRU  F-1065
transform 1 0 2850 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1066
transform 1 0 2818 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1067
transform 1 0 2841 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1068
transform 1 0 2854 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1069
transform 1 0 2838 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1070
transform 1 0 2892 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1071
transform 1 0 2849 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1072
transform 1 0 2803 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1073
transform 1 0 2696 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-1074
transform 1 0 2676 0 1 5810
box 0 0 3 6
use FEEDTHRU  F-1075
transform 1 0 2660 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1076
transform 1 0 2782 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1077
transform 1 0 2830 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1078
transform 1 0 2810 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1079
transform 1 0 2837 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1080
transform 1 0 2879 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1081
transform 1 0 2741 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1082
transform 1 0 2865 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1083
transform 1 0 2902 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1084
transform 1 0 2800 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1085
transform 1 0 3105 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1086
transform 1 0 3123 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1087
transform 1 0 3086 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1088
transform 1 0 3064 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1089
transform 1 0 3046 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1090
transform 1 0 2814 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1091
transform 1 0 2826 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1092
transform 1 0 2857 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1093
transform 1 0 3143 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1094
transform 1 0 2733 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1095
transform 1 0 2978 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1096
transform 1 0 2981 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1097
transform 1 0 2963 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1098
transform 1 0 3074 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1099
transform 1 0 2713 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1100
transform 1 0 2759 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1101
transform 1 0 2776 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1102
transform 1 0 2788 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1103
transform 1 0 3001 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1104
transform 1 0 3013 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1105
transform 1 0 3001 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1106
transform 1 0 2924 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1107
transform 1 0 2833 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1108
transform 1 0 2809 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1109
transform 1 0 2884 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1110
transform 1 0 2881 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1111
transform 1 0 2957 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1112
transform 1 0 3015 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1113
transform 1 0 2871 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1114
transform 1 0 2884 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1115
transform 1 0 2993 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1116
transform 1 0 3000 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1117
transform 1 0 3046 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1118
transform 1 0 3154 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1119
transform 1 0 3124 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1120
transform 1 0 3085 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1121
transform 1 0 3154 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1122
transform 1 0 3121 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1123
transform 1 0 3084 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1124
transform 1 0 3106 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1125
transform 1 0 3034 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1126
transform 1 0 3004 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1127
transform 1 0 2964 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1128
transform 1 0 2957 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1129
transform 1 0 2921 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1130
transform 1 0 2918 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1131
transform 1 0 3163 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1132
transform 1 0 3116 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1133
transform 1 0 2954 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1134
transform 1 0 2957 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1135
transform 1 0 2990 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1136
transform 1 0 2997 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1137
transform 1 0 3016 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1138
transform 1 0 3028 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1139
transform 1 0 3036 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1140
transform 1 0 3115 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1141
transform 1 0 2777 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1142
transform 1 0 2790 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1143
transform 1 0 3014 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1144
transform 1 0 3114 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1145
transform 1 0 3134 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1146
transform 1 0 3127 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1147
transform 1 0 2907 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1148
transform 1 0 2865 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1149
transform 1 0 2878 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1150
transform 1 0 2867 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1151
transform 1 0 2810 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1152
transform 1 0 2846 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1153
transform 1 0 2844 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1154
transform 1 0 2935 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1155
transform 1 0 2965 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1156
transform 1 0 2822 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1157
transform 1 0 2858 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1158
transform 1 0 2859 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1159
transform 1 0 3013 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1160
transform 1 0 2946 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1161
transform 1 0 2980 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1162
transform 1 0 2952 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1163
transform 1 0 2983 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1164
transform 1 0 2977 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1165
transform 1 0 2940 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1166
transform 1 0 3007 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1167
transform 1 0 2959 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1168
transform 1 0 2905 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1169
transform 1 0 2865 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1170
transform 1 0 2870 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1171
transform 1 0 2846 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1172
transform 1 0 2919 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1173
transform 1 0 3154 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1174
transform 1 0 3118 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1175
transform 1 0 3140 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1176
transform 1 0 3030 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1177
transform 1 0 3017 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1178
transform 1 0 2990 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1179
transform 1 0 3011 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1180
transform 1 0 3118 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1181
transform 1 0 3175 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1182
transform 1 0 3121 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1183
transform 1 0 3183 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1184
transform 1 0 3184 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1185
transform 1 0 3145 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1186
transform 1 0 3085 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1187
transform 1 0 3072 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1188
transform 1 0 3158 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1189
transform 1 0 3035 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1190
transform 1 0 3020 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1191
transform 1 0 3025 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1192
transform 1 0 2964 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1193
transform 1 0 2913 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1194
transform 1 0 2912 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1195
transform 1 0 2894 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1196
transform 1 0 2876 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1197
transform 1 0 2866 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1198
transform 1 0 2836 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1199
transform 1 0 3148 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1200
transform 1 0 3187 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1201
transform 1 0 3186 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1202
transform 1 0 3124 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1203
transform 1 0 3075 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1204
transform 1 0 3026 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1205
transform 1 0 2920 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1206
transform 1 0 2871 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1207
transform 1 0 3043 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1208
transform 1 0 3042 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1209
transform 1 0 3128 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1210
transform 1 0 3146 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1211
transform 1 0 3183 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1212
transform 1 0 3107 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1213
transform 1 0 3163 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1214
transform 1 0 3196 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1215
transform 1 0 3195 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1216
transform 1 0 3133 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1217
transform 1 0 3268 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1218
transform 1 0 3046 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1219
transform 1 0 3045 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1220
transform 1 0 3047 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1221
transform 1 0 3062 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1222
transform 1 0 3087 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1223
transform 1 0 3101 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1224
transform 1 0 3157 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1225
transform 1 0 2825 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1226
transform 1 0 2855 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1227
transform 1 0 2836 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1228
transform 1 0 2771 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1229
transform 1 0 3019 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1230
transform 1 0 2820 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1231
transform 1 0 2832 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1232
transform 1 0 2869 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1233
transform 1 0 2828 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1234
transform 1 0 2838 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1235
transform 1 0 2772 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1236
transform 1 0 2778 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1237
transform 1 0 2765 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1238
transform 1 0 2777 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1239
transform 1 0 2810 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1240
transform 1 0 2808 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1241
transform 1 0 2808 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1242
transform 1 0 2845 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1243
transform 1 0 2839 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1244
transform 1 0 2829 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1245
transform 1 0 2836 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1246
transform 1 0 2868 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1247
transform 1 0 2865 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1248
transform 1 0 2896 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1249
transform 1 0 2895 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1250
transform 1 0 2913 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1251
transform 1 0 2931 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1252
transform 1 0 2965 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1253
transform 1 0 2824 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1254
transform 1 0 2811 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1255
transform 1 0 2821 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1256
transform 1 0 2917 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1257
transform 1 0 2901 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1258
transform 1 0 2900 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1259
transform 1 0 2870 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1260
transform 1 0 2858 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1261
transform 1 0 2848 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1262
transform 1 0 2773 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1263
transform 1 0 2756 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1264
transform 1 0 2877 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1265
transform 1 0 2929 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1266
transform 1 0 2887 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1267
transform 1 0 2917 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1268
transform 1 0 2767 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1269
transform 1 0 2768 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-1270
transform 1 0 2770 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1271
transform 1 0 2817 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1272
transform 1 0 2863 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1273
transform 1 0 2771 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-1274
transform 1 0 2755 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1275
transform 1 0 3094 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1276
transform 1 0 3151 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1277
transform 1 0 3097 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1278
transform 1 0 3082 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1279
transform 1 0 3136 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1280
transform 1 0 2862 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1281
transform 1 0 2917 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1282
transform 1 0 2859 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1283
transform 1 0 2936 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1284
transform 1 0 2944 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1285
transform 1 0 2818 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1286
transform 1 0 3124 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1287
transform 1 0 3091 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1288
transform 1 0 3144 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1289
transform 1 0 3142 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1290
transform 1 0 3130 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1291
transform 1 0 2975 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1292
transform 1 0 2933 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1293
transform 1 0 2930 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1294
transform 1 0 2947 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1295
transform 1 0 2875 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1296
transform 1 0 3264 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1297
transform 1 0 3290 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1298
transform 1 0 3235 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1299
transform 1 0 3208 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1300
transform 1 0 3157 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1301
transform 1 0 3223 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1302
transform 1 0 3176 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1303
transform 1 0 3293 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1304
transform 1 0 2977 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1305
transform 1 0 2986 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1306
transform 1 0 2926 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1307
transform 1 0 2953 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1308
transform 1 0 2913 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1309
transform 1 0 2925 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1310
transform 1 0 2926 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1311
transform 1 0 2869 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1312
transform 1 0 2902 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1313
transform 1 0 2908 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1314
transform 1 0 2987 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1315
transform 1 0 2899 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1316
transform 1 0 2902 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1317
transform 1 0 3040 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1318
transform 1 0 2738 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1319
transform 1 0 2788 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1320
transform 1 0 2796 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1321
transform 1 0 2783 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1322
transform 1 0 2792 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1323
transform 1 0 2834 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1324
transform 1 0 2826 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1325
transform 1 0 2696 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1326
transform 1 0 2728 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1327
transform 1 0 2805 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1328
transform 1 0 2789 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1329
transform 1 0 2798 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1330
transform 1 0 2840 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1331
transform 1 0 2832 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1332
transform 1 0 2838 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1333
transform 1 0 2881 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1334
transform 1 0 2869 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1335
transform 1 0 2874 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1336
transform 1 0 2892 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1337
transform 1 0 2884 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1338
transform 1 0 2908 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1339
transform 1 0 2799 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1340
transform 1 0 2799 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1341
transform 1 0 3218 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1342
transform 1 0 3176 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1343
transform 1 0 3234 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1344
transform 1 0 3196 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1345
transform 1 0 3139 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1346
transform 1 0 3076 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1347
transform 1 0 3154 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1348
transform 1 0 3094 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1349
transform 1 0 2906 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1350
transform 1 0 2929 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1351
transform 1 0 2887 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1352
transform 1 0 2957 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1353
transform 1 0 3010 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1354
transform 1 0 3163 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1355
transform 1 0 3155 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1356
transform 1 0 3128 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1357
transform 1 0 3148 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1358
transform 1 0 3106 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1359
transform 1 0 3093 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1360
transform 1 0 3037 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1361
transform 1 0 2995 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1362
transform 1 0 2953 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1363
transform 1 0 2934 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1364
transform 1 0 2960 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1365
transform 1 0 2964 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1366
transform 1 0 2982 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1367
transform 1 0 2761 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1368
transform 1 0 2820 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1369
transform 1 0 2863 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1370
transform 1 0 2851 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1371
transform 1 0 2797 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1372
transform 1 0 2854 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1373
transform 1 0 2864 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1374
transform 1 0 2753 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1375
transform 1 0 2977 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1376
transform 1 0 2995 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1377
transform 1 0 2962 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1378
transform 1 0 2912 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1379
transform 1 0 2763 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-1380
transform 1 0 2739 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-1381
transform 1 0 2799 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1382
transform 1 0 2765 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1383
transform 1 0 2809 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1384
transform 1 0 2947 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1385
transform 1 0 3165 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1386
transform 1 0 3163 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1387
transform 1 0 3121 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1388
transform 1 0 3070 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1389
transform 1 0 3066 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1390
transform 1 0 3032 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1391
transform 1 0 3134 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1392
transform 1 0 2999 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1393
transform 1 0 2998 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1394
transform 1 0 2943 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1395
transform 1 0 2903 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1396
transform 1 0 2826 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1397
transform 1 0 2838 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-1398
transform 1 0 2848 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1399
transform 1 0 2802 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1400
transform 1 0 3043 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1401
transform 1 0 3067 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1402
transform 1 0 3066 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1403
transform 1 0 3034 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1404
transform 1 0 3079 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1405
transform 1 0 3103 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1406
transform 1 0 3082 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1407
transform 1 0 3060 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1408
transform 1 0 3093 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1409
transform 1 0 3089 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1410
transform 1 0 2986 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1411
transform 1 0 2750 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1412
transform 1 0 2803 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1413
transform 1 0 2867 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1414
transform 1 0 2966 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1415
transform 1 0 3002 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1416
transform 1 0 3012 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1417
transform 1 0 3028 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1418
transform 1 0 3082 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1419
transform 1 0 3109 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1420
transform 1 0 3237 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1421
transform 1 0 3167 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1422
transform 1 0 3208 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1423
transform 1 0 3046 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1424
transform 1 0 3145 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1425
transform 1 0 3165 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1426
transform 1 0 3204 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1427
transform 1 0 3197 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1428
transform 1 0 3106 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1429
transform 1 0 3067 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1430
transform 1 0 3016 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1431
transform 1 0 2963 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1432
transform 1 0 2887 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1433
transform 1 0 2829 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1434
transform 1 0 2772 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-1435
transform 1 0 2736 0 1 5810
box 0 0 3 6
use FEEDTHRU  F-1436
transform 1 0 2714 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1437
transform 1 0 2701 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1438
transform 1 0 3036 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1439
transform 1 0 2923 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1440
transform 1 0 2884 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1441
transform 1 0 2935 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1442
transform 1 0 2877 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1443
transform 1 0 2926 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1444
transform 1 0 2925 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1445
transform 1 0 2952 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1446
transform 1 0 3105 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1447
transform 1 0 3111 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1448
transform 1 0 3149 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1449
transform 1 0 3100 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1450
transform 1 0 3097 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1451
transform 1 0 3129 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1452
transform 1 0 3052 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1453
transform 1 0 3006 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1454
transform 1 0 3049 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1455
transform 1 0 3085 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1456
transform 1 0 3108 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1457
transform 1 0 3156 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1458
transform 1 0 3002 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1459
transform 1 0 2993 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1460
transform 1 0 3039 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1461
transform 1 0 3004 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1462
transform 1 0 2875 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1463
transform 1 0 2893 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1464
transform 1 0 2844 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1465
transform 1 0 2865 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1466
transform 1 0 2869 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1467
transform 1 0 2929 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1468
transform 1 0 2893 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1469
transform 1 0 3208 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1470
transform 1 0 3282 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1471
transform 1 0 3005 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1472
transform 1 0 3023 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1473
transform 1 0 3044 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1474
transform 1 0 3060 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1475
transform 1 0 2871 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1476
transform 1 0 2878 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1477
transform 1 0 3049 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1478
transform 1 0 3003 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1479
transform 1 0 2828 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1480
transform 1 0 2840 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1481
transform 1 0 2882 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1482
transform 1 0 2877 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1483
transform 1 0 2899 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1484
transform 1 0 2947 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1485
transform 1 0 2941 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1486
transform 1 0 2919 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1487
transform 1 0 2902 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1488
transform 1 0 2959 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1489
transform 1 0 2901 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1490
transform 1 0 2950 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1491
transform 1 0 2955 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1492
transform 1 0 2760 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1493
transform 1 0 3253 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1494
transform 1 0 3305 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1495
transform 1 0 3178 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1496
transform 1 0 3085 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1497
transform 1 0 3138 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1498
transform 1 0 3136 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1499
transform 1 0 3127 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1500
transform 1 0 3052 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1501
transform 1 0 2743 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1502
transform 1 0 2786 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1503
transform 1 0 2800 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1504
transform 1 0 2824 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1505
transform 1 0 2842 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1506
transform 1 0 2740 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1507
transform 1 0 2783 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1508
transform 1 0 2806 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1509
transform 1 0 2830 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1510
transform 1 0 2854 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1511
transform 1 0 2909 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1512
transform 1 0 2976 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1513
transform 1 0 2931 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1514
transform 1 0 2932 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1515
transform 1 0 2883 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1516
transform 1 0 2982 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1517
transform 1 0 2986 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1518
transform 1 0 2978 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1519
transform 1 0 3030 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1520
transform 1 0 2979 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1521
transform 1 0 2974 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1522
transform 1 0 2802 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1523
transform 1 0 2746 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1524
transform 1 0 2708 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1525
transform 1 0 3110 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1526
transform 1 0 3037 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1527
transform 1 0 2986 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1528
transform 1 0 2935 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1529
transform 1 0 2897 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1530
transform 1 0 2991 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1531
transform 1 0 2917 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1532
transform 1 0 2938 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1533
transform 1 0 2965 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1534
transform 1 0 3133 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1535
transform 1 0 3329 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1536
transform 1 0 3162 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1537
transform 1 0 3169 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1538
transform 1 0 3142 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1539
transform 1 0 2819 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1540
transform 1 0 2860 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1541
transform 1 0 2860 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1542
transform 1 0 2925 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1543
transform 1 0 2918 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1544
transform 1 0 2888 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1545
transform 1 0 2950 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1546
transform 1 0 2977 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1547
transform 1 0 2686 0 1 1280
box 0 0 3 6
use FEEDTHRU  F-1548
transform 1 0 2858 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1549
transform 1 0 2834 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1550
transform 1 0 2891 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1551
transform 1 0 2911 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1552
transform 1 0 2917 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1553
transform 1 0 2883 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1554
transform 1 0 3006 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1555
transform 1 0 2794 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1556
transform 1 0 3126 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1557
transform 1 0 3098 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1558
transform 1 0 3013 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1559
transform 1 0 3057 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1560
transform 1 0 3022 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1561
transform 1 0 2982 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1562
transform 1 0 3061 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1563
transform 1 0 3010 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1564
transform 1 0 3024 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1565
transform 1 0 3087 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1566
transform 1 0 3038 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1567
transform 1 0 2968 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1568
transform 1 0 2980 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1569
transform 1 0 2947 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1570
transform 1 0 3276 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1571
transform 1 0 2538 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1572
transform 1 0 2619 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1573
transform 1 0 2658 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1574
transform 1 0 2712 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1575
transform 1 0 2695 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1576
transform 1 0 2716 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1577
transform 1 0 2747 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1578
transform 1 0 2753 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1579
transform 1 0 2754 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1580
transform 1 0 2800 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1581
transform 1 0 2797 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1582
transform 1 0 2790 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1583
transform 1 0 2764 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1584
transform 1 0 2808 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1585
transform 1 0 2757 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1586
transform 1 0 2812 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1587
transform 1 0 2796 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1588
transform 1 0 2856 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1589
transform 1 0 2795 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1590
transform 1 0 2731 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1591
transform 1 0 2856 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1592
transform 1 0 2850 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1593
transform 1 0 2868 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1594
transform 1 0 2917 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1595
transform 1 0 2912 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1596
transform 1 0 2716 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1597
transform 1 0 2663 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-1598
transform 1 0 2850 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1599
transform 1 0 2818 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1600
transform 1 0 2789 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1601
transform 1 0 2755 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1602
transform 1 0 3255 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1603
transform 1 0 3067 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1604
transform 1 0 3072 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1605
transform 1 0 2872 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1606
transform 1 0 2832 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1607
transform 1 0 3004 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1608
transform 1 0 2965 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1609
transform 1 0 2952 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1610
transform 1 0 2945 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1611
transform 1 0 2912 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1612
transform 1 0 2927 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1613
transform 1 0 2890 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1614
transform 1 0 2845 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1615
transform 1 0 2799 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1616
transform 1 0 2722 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1617
transform 1 0 3063 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1618
transform 1 0 3055 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1619
transform 1 0 3040 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1620
transform 1 0 3060 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1621
transform 1 0 2833 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1622
transform 1 0 2884 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1623
transform 1 0 2882 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1624
transform 1 0 2906 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1625
transform 1 0 2939 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1626
transform 1 0 2946 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1627
transform 1 0 3084 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1628
transform 1 0 3122 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1629
transform 1 0 3151 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1630
transform 1 0 3136 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1631
transform 1 0 3221 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1632
transform 1 0 2762 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1633
transform 1 0 2824 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1634
transform 1 0 2885 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1635
transform 1 0 2923 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1636
transform 1 0 2956 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1637
transform 1 0 2950 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1638
transform 1 0 3019 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1639
transform 1 0 3017 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1640
transform 1 0 2993 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1641
transform 1 0 3013 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1642
transform 1 0 2958 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1643
transform 1 0 2912 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1644
transform 1 0 2968 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1645
transform 1 0 2877 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1646
transform 1 0 2931 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1647
transform 1 0 2873 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1648
transform 1 0 2890 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1649
transform 1 0 2835 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1650
transform 1 0 2933 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1651
transform 1 0 2860 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1652
transform 1 0 3076 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1653
transform 1 0 2899 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1654
transform 1 0 2862 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1655
transform 1 0 2853 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1656
transform 1 0 2960 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1657
transform 1 0 3013 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1658
transform 1 0 3007 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1659
transform 1 0 2995 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1660
transform 1 0 3080 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1661
transform 1 0 2852 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1662
transform 1 0 2888 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1663
transform 1 0 2895 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1664
transform 1 0 2822 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1665
transform 1 0 2833 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1666
transform 1 0 2785 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1667
transform 1 0 2735 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1668
transform 1 0 2965 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1669
transform 1 0 3078 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1670
transform 1 0 3227 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1671
transform 1 0 3280 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1672
transform 1 0 2773 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1673
transform 1 0 2817 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1674
transform 1 0 2772 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1675
transform 1 0 2827 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1676
transform 1 0 2817 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1677
transform 1 0 2871 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1678
transform 1 0 2816 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1679
transform 1 0 2746 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1680
transform 1 0 2737 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1681
transform 1 0 2731 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1682
transform 1 0 2694 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1683
transform 1 0 2652 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1684
transform 1 0 2580 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1685
transform 1 0 2664 0 1 5810
box 0 0 3 6
use FEEDTHRU  F-1686
transform 1 0 2684 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-1687
transform 1 0 2690 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-1688
transform 1 0 2926 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1689
transform 1 0 2908 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1690
transform 1 0 2861 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1691
transform 1 0 2773 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1692
transform 1 0 3042 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1693
transform 1 0 3088 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1694
transform 1 0 2874 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1695
transform 1 0 2923 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1696
transform 1 0 2905 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1697
transform 1 0 2907 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1698
transform 1 0 2850 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1699
transform 1 0 2893 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1700
transform 1 0 2532 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-1701
transform 1 0 2544 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1702
transform 1 0 2645 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1703
transform 1 0 2946 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1704
transform 1 0 2907 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1705
transform 1 0 2914 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1706
transform 1 0 2859 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1707
transform 1 0 2956 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1708
transform 1 0 3138 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1709
transform 1 0 3066 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1710
transform 1 0 3061 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1711
transform 1 0 3092 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1712
transform 1 0 2977 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1713
transform 1 0 2938 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1714
transform 1 0 2970 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1715
transform 1 0 2971 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1716
transform 1 0 2830 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1717
transform 1 0 2848 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1718
transform 1 0 2848 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1719
transform 1 0 2915 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1720
transform 1 0 2970 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1721
transform 1 0 2879 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1722
transform 1 0 2974 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1723
transform 1 0 3054 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1724
transform 1 0 3110 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1725
transform 1 0 3182 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1726
transform 1 0 3040 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1727
transform 1 0 3122 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1728
transform 1 0 3262 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1729
transform 1 0 3226 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1730
transform 1 0 3091 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1731
transform 1 0 2845 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1732
transform 1 0 2814 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1733
transform 1 0 2745 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-1734
transform 1 0 3145 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1735
transform 1 0 3076 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1736
transform 1 0 3147 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1737
transform 1 0 3091 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1738
transform 1 0 3102 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1739
transform 1 0 2953 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1740
transform 1 0 2958 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1741
transform 1 0 2908 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1742
transform 1 0 2816 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1743
transform 1 0 2852 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1744
transform 1 0 2945 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1745
transform 1 0 2740 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1746
transform 1 0 2750 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-1747
transform 1 0 2698 0 1 1280
box 0 0 3 6
use FEEDTHRU  F-1748
transform 1 0 2795 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1749
transform 1 0 2836 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1750
transform 1 0 2801 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1751
transform 1 0 2854 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1752
transform 1 0 2854 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1753
transform 1 0 2810 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1754
transform 1 0 2749 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1755
transform 1 0 2695 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1756
transform 1 0 2706 0 1 5810
box 0 0 3 6
use FEEDTHRU  F-1757
transform 1 0 2727 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-1758
transform 1 0 2771 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1759
transform 1 0 2827 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1760
transform 1 0 2709 0 1 5810
box 0 0 3 6
use FEEDTHRU  F-1761
transform 1 0 2730 0 1 5777
box 0 0 3 6
use FEEDTHRU  F-1762
transform 1 0 3001 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1763
transform 1 0 2989 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1764
transform 1 0 2994 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1765
transform 1 0 2995 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1766
transform 1 0 3022 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1767
transform 1 0 2937 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1768
transform 1 0 2983 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1769
transform 1 0 2689 0 1 1280
box 0 0 3 6
use FEEDTHRU  F-1770
transform 1 0 2726 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-1771
transform 1 0 2725 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1772
transform 1 0 2802 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1773
transform 1 0 2839 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1774
transform 1 0 2914 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1775
transform 1 0 2857 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1776
transform 1 0 2823 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1777
transform 1 0 2743 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1778
transform 1 0 2753 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-1779
transform 1 0 2867 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1780
transform 1 0 2959 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1781
transform 1 0 2954 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1782
transform 1 0 3066 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1783
transform 1 0 3034 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1784
transform 1 0 3124 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1785
transform 1 0 2950 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1786
transform 1 0 2896 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1787
transform 1 0 2876 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1788
transform 1 0 2908 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1789
transform 1 0 2998 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1790
transform 1 0 3042 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1791
transform 1 0 2683 0 1 1280
box 0 0 3 6
use FEEDTHRU  F-1792
transform 1 0 3055 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1793
transform 1 0 3128 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1794
transform 1 0 2905 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1795
transform 1 0 2881 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1796
transform 1 0 2889 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1797
transform 1 0 2842 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1798
transform 1 0 2899 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1799
transform 1 0 2891 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1800
transform 1 0 2941 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1801
transform 1 0 2968 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1802
transform 1 0 2956 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1803
transform 1 0 3032 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1804
transform 1 0 3081 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1805
transform 1 0 3018 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1806
transform 1 0 3016 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1807
transform 1 0 2970 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1808
transform 1 0 3049 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1809
transform 1 0 2980 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1810
transform 1 0 2879 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1811
transform 1 0 2929 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1812
transform 1 0 2944 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1813
transform 1 0 2938 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1814
transform 1 0 3020 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1815
transform 1 0 3066 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1816
transform 1 0 2962 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1817
transform 1 0 2851 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1818
transform 1 0 2807 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1819
transform 1 0 2737 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1820
transform 1 0 2680 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1821
transform 1 0 2999 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1822
transform 1 0 2972 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1823
transform 1 0 2881 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1824
transform 1 0 2866 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1825
transform 1 0 2942 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1826
transform 1 0 3000 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1827
transform 1 0 2943 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1828
transform 1 0 3132 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1829
transform 1 0 3058 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1830
transform 1 0 3037 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1831
transform 1 0 3019 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1832
transform 1 0 3030 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1833
transform 1 0 3054 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1834
transform 1 0 3038 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1835
transform 1 0 3005 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1836
transform 1 0 2975 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1837
transform 1 0 3001 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1838
transform 1 0 2961 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1839
transform 1 0 2915 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1840
transform 1 0 2823 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1841
transform 1 0 2829 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-1842
transform 1 0 2903 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1843
transform 1 0 2827 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1844
transform 1 0 2842 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1845
transform 1 0 2948 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1846
transform 1 0 3012 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1847
transform 1 0 2853 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1848
transform 1 0 2911 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1849
transform 1 0 2851 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1850
transform 1 0 2901 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1851
transform 1 0 2899 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1852
transform 1 0 2887 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1853
transform 1 0 2911 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1854
transform 1 0 2883 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1855
transform 1 0 2958 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1856
transform 1 0 2889 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1857
transform 1 0 3043 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1858
transform 1 0 2958 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1859
transform 1 0 2889 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1860
transform 1 0 2692 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1861
transform 1 0 2746 0 1 5599
box 0 0 3 6
use FEEDTHRU  F-1862
transform 1 0 2962 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1863
transform 1 0 2939 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1864
transform 1 0 2960 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1865
transform 1 0 2962 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1866
transform 1 0 2902 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1867
transform 1 0 2850 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1868
transform 1 0 3019 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1869
transform 1 0 2746 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1870
transform 1 0 2747 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-1871
transform 1 0 2701 0 1 1280
box 0 0 3 6
use FEEDTHRU  F-1872
transform 1 0 3192 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1873
transform 1 0 3117 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1874
transform 1 0 3119 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1875
transform 1 0 2974 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1876
transform 1 0 2992 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1877
transform 1 0 2848 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1878
transform 1 0 2863 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1879
transform 1 0 2839 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1880
transform 1 0 2921 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1881
transform 1 0 2988 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1882
transform 1 0 2913 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1883
transform 1 0 2908 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1884
transform 1 0 2919 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1885
transform 1 0 2989 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1886
transform 1 0 2914 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1887
transform 1 0 2964 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1888
transform 1 0 2959 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1889
transform 1 0 2983 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1890
transform 1 0 2923 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1891
transform 1 0 2911 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1892
transform 1 0 3113 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1893
transform 1 0 2801 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1894
transform 1 0 2828 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1895
transform 1 0 2864 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1896
transform 1 0 3054 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1897
transform 1 0 2878 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1898
transform 1 0 2954 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1899
transform 1 0 2683 0 1 5706
box 0 0 3 6
use FEEDTHRU  F-1900
transform 1 0 2951 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1901
transform 1 0 2958 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1902
transform 1 0 2959 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1903
transform 1 0 3016 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1904
transform 1 0 2995 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1905
transform 1 0 3012 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1906
transform 1 0 2956 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1907
transform 1 0 3031 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1908
transform 1 0 2940 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1909
transform 1 0 2998 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1910
transform 1 0 3000 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1911
transform 1 0 3075 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1912
transform 1 0 3014 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1913
transform 1 0 2932 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1914
transform 1 0 2950 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1915
transform 1 0 2984 0 1 4666
box 0 0 3 6
use FEEDTHRU  F-1916
transform 1 0 3048 0 1 4421
box 0 0 3 6
use FEEDTHRU  F-1917
transform 1 0 2973 0 1 4212
box 0 0 3 6
use FEEDTHRU  F-1918
transform 1 0 2968 0 1 4017
box 0 0 3 6
use FEEDTHRU  F-1919
transform 1 0 2913 0 1 3796
box 0 0 3 6
use FEEDTHRU  F-1920
transform 1 0 2995 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1921
transform 1 0 2920 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1922
transform 1 0 2976 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1923
transform 1 0 2965 0 1 2876
box 0 0 3 6
use FEEDTHRU  F-1924
transform 1 0 2989 0 1 2663
box 0 0 3 6
use FEEDTHRU  F-1925
transform 1 0 2929 0 1 2462
box 0 0 3 6
use FEEDTHRU  F-1926
transform 1 0 2928 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1927
transform 1 0 2921 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1928
transform 1 0 2882 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1929
transform 1 0 2852 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1930
transform 1 0 2872 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1931
transform 1 0 2821 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1932
transform 1 0 2768 0 1 1477
box 0 0 3 6
use FEEDTHRU  F-1933
transform 1 0 3013 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1934
transform 1 0 2932 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1935
transform 1 0 2988 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1936
transform 1 0 2953 0 1 3543
box 0 0 3 6
use FEEDTHRU  F-1937
transform 1 0 2875 0 1 3348
box 0 0 3 6
use FEEDTHRU  F-1938
transform 1 0 2931 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1939
transform 1 0 2883 0 1 2293
box 0 0 3 6
use FEEDTHRU  F-1940
transform 1 0 2876 0 1 2132
box 0 0 3 6
use FEEDTHRU  F-1941
transform 1 0 2834 0 1 1967
box 0 0 3 6
use FEEDTHRU  F-1942
transform 1 0 2807 0 1 1818
box 0 0 3 6
use FEEDTHRU  F-1943
transform 1 0 2827 0 1 1679
box 0 0 3 6
use FEEDTHRU  F-1944
transform 1 0 2779 0 1 1574
box 0 0 3 6
use FEEDTHRU  F-1945
transform 1 0 2872 0 1 4887
box 0 0 3 6
use FEEDTHRU  F-1946
transform 1 0 2887 0 1 5072
box 0 0 3 6
use FEEDTHRU  F-1947
transform 1 0 2872 0 1 5265
box 0 0 3 6
use FEEDTHRU  F-1948
transform 1 0 2822 0 1 5442
box 0 0 3 6
use FEEDTHRU  F-1949
transform 1 0 3078 0 1 3107
box 0 0 3 6
use FEEDTHRU  F-1950
transform 1 0 2865 0 1 1384
box 0 0 3 6
use FEEDTHRU  F-1951
transform 1 0 2780 0 1 1331
box 0 0 3 6
use FEEDTHRU  F-1952
transform 1 0 2914 0 1 5072
box 0 0 3 6
<< metal1 >>
rect 2641 1271 2738 1272
rect 2644 1273 2648 1274
rect 2671 1273 2685 1274
rect 2678 1275 2688 1276
rect 2690 1275 2694 1276
rect 2699 1275 2709 1276
rect 2702 1277 2706 1278
rect 2527 1287 2534 1288
rect 2605 1287 2840 1288
rect 2626 1289 2646 1290
rect 2633 1291 2663 1292
rect 2641 1293 2678 1294
rect 2642 1295 2656 1296
rect 2647 1297 2675 1298
rect 2684 1297 2715 1298
rect 2687 1299 2722 1300
rect 2680 1301 2687 1302
rect 2690 1301 2728 1302
rect 2692 1303 2731 1304
rect 2696 1305 2712 1306
rect 2699 1307 2752 1308
rect 2699 1309 2709 1310
rect 2702 1311 2749 1312
rect 2737 1313 2828 1314
rect 2754 1315 2816 1316
rect 2757 1317 2852 1318
rect 2760 1319 2776 1320
rect 2769 1321 2795 1322
rect 2772 1323 2792 1324
rect 2781 1325 2846 1326
rect 2784 1327 2825 1328
rect 2798 1329 2831 1330
rect 2521 1338 2540 1339
rect 2533 1340 2546 1341
rect 2533 1342 2543 1343
rect 2587 1342 2597 1343
rect 2593 1344 2649 1345
rect 2626 1346 2690 1347
rect 2630 1348 2643 1349
rect 2633 1350 2646 1351
rect 2617 1352 2647 1353
rect 2665 1352 2712 1353
rect 2668 1354 2675 1355
rect 2623 1356 2675 1357
rect 2671 1358 2678 1359
rect 2680 1358 2687 1359
rect 2704 1358 2709 1359
rect 2723 1358 2799 1359
rect 2741 1360 2752 1361
rect 2744 1362 2755 1363
rect 2750 1364 2758 1365
rect 2753 1366 2761 1367
rect 2756 1368 2773 1369
rect 2769 1370 2772 1371
rect 2768 1372 2795 1373
rect 2781 1374 2867 1375
rect 2792 1376 2806 1377
rect 2808 1376 2864 1377
rect 2815 1378 2837 1379
rect 2827 1380 2834 1381
rect 2827 1382 2840 1383
rect 2875 1382 2896 1383
rect 2539 1391 2621 1392
rect 2542 1393 2562 1394
rect 2533 1395 2544 1396
rect 2549 1395 2559 1396
rect 2564 1395 2862 1396
rect 2593 1397 2612 1398
rect 2608 1399 2662 1400
rect 2614 1401 2722 1402
rect 2617 1403 2683 1404
rect 2623 1405 2644 1406
rect 2623 1407 2716 1408
rect 2626 1409 2710 1410
rect 2629 1411 2707 1412
rect 2630 1413 2740 1414
rect 2633 1415 2698 1416
rect 2637 1417 2737 1418
rect 2652 1419 2665 1420
rect 2668 1419 2704 1420
rect 2671 1421 2686 1422
rect 2700 1421 2767 1422
rect 2711 1423 2783 1424
rect 2646 1425 2713 1426
rect 2545 1427 2647 1428
rect 2723 1427 2801 1428
rect 2726 1429 2804 1430
rect 2741 1431 2858 1432
rect 2747 1433 2869 1434
rect 2750 1435 2807 1436
rect 2753 1437 2810 1438
rect 2754 1439 2761 1440
rect 2756 1441 2840 1442
rect 2757 1443 2837 1444
rect 2763 1445 2769 1446
rect 2769 1447 2910 1448
rect 2771 1449 2819 1450
rect 2680 1451 2773 1452
rect 2679 1453 2878 1454
rect 2778 1455 2822 1456
rect 2792 1457 2849 1458
rect 2824 1459 2917 1460
rect 2744 1461 2825 1462
rect 2827 1461 2905 1462
rect 2830 1463 2887 1464
rect 2833 1465 2890 1466
rect 2798 1467 2834 1468
rect 2851 1467 2908 1468
rect 2863 1469 2940 1470
rect 2866 1471 2946 1472
rect 2875 1473 2957 1474
rect 2815 1475 2875 1476
rect 2910 1475 2914 1476
rect 2551 1484 2559 1485
rect 2611 1484 2637 1485
rect 2617 1486 2781 1487
rect 2620 1488 2660 1489
rect 2623 1490 2713 1491
rect 2626 1492 2678 1493
rect 2630 1494 2716 1495
rect 2649 1496 2707 1497
rect 2661 1498 2784 1499
rect 2643 1500 2663 1501
rect 2674 1500 2763 1501
rect 2679 1502 2969 1503
rect 2685 1504 2712 1505
rect 2689 1506 2966 1507
rect 2693 1508 2755 1509
rect 2697 1510 2730 1511
rect 2696 1512 2799 1513
rect 2703 1514 2718 1515
rect 2709 1516 2748 1517
rect 2739 1518 2790 1519
rect 2800 1518 2847 1519
rect 2671 1520 2802 1521
rect 2803 1520 2841 1521
rect 2806 1522 2832 1523
rect 2818 1524 2865 1525
rect 2809 1526 2820 1527
rect 2766 1528 2811 1529
rect 2682 1530 2766 1531
rect 2824 1530 2859 1531
rect 2772 1532 2826 1533
rect 2848 1532 2901 1533
rect 2785 1534 2850 1535
rect 2736 1536 2787 1537
rect 2735 1538 2779 1539
rect 2868 1538 2893 1539
rect 2646 1540 2892 1541
rect 2646 1542 2653 1543
rect 2874 1542 2988 1543
rect 2833 1544 2874 1545
rect 2775 1546 2835 1547
rect 2757 1548 2775 1549
rect 2686 1550 2757 1551
rect 2877 1550 2898 1551
rect 2721 1552 2877 1553
rect 2664 1554 2721 1555
rect 2886 1554 2954 1555
rect 2821 1556 2886 1557
rect 2769 1558 2823 1559
rect 2904 1558 2945 1559
rect 2851 1560 2904 1561
rect 2913 1560 2960 1561
rect 2916 1562 2963 1563
rect 2939 1564 3005 1565
rect 2956 1566 3008 1567
rect 2889 1568 2957 1569
rect 2760 1570 2889 1571
rect 2971 1570 2981 1571
rect 2974 1572 2978 1573
rect 2560 1581 2652 1582
rect 2563 1583 2655 1584
rect 2605 1585 3105 1586
rect 2656 1587 2763 1588
rect 2659 1589 2714 1590
rect 2662 1591 2686 1592
rect 2667 1593 2766 1594
rect 2693 1595 2792 1596
rect 2711 1597 2759 1598
rect 2717 1599 2765 1600
rect 2677 1601 2717 1602
rect 2636 1603 2677 1604
rect 2720 1603 2795 1604
rect 2722 1605 2865 1606
rect 2729 1607 2807 1608
rect 2747 1609 2804 1610
rect 2746 1611 2757 1612
rect 2768 1611 2862 1612
rect 2780 1613 2829 1614
rect 2631 1615 2780 1616
rect 2783 1615 2832 1616
rect 2626 1617 2783 1618
rect 2798 1617 2856 1618
rect 2789 1619 2798 1620
rect 2810 1619 2813 1620
rect 2837 1619 2868 1620
rect 2638 1621 2838 1622
rect 2846 1621 2892 1622
rect 2708 1623 2847 1624
rect 2623 1625 2708 1626
rect 2849 1625 2895 1626
rect 2774 1627 2850 1628
rect 2634 1629 2774 1630
rect 2873 1629 2914 1630
rect 2819 1631 2913 1632
rect 2819 1633 2841 1634
rect 2822 1635 2874 1636
rect 2876 1635 2949 1636
rect 2825 1637 2877 1638
rect 2649 1639 2826 1640
rect 2885 1639 2928 1640
rect 2834 1641 2886 1642
rect 2786 1643 2835 1644
rect 2888 1643 2931 1644
rect 2771 1645 2889 1646
rect 2735 1647 2771 1648
rect 2612 1649 2735 1650
rect 2897 1649 2952 1650
rect 2916 1651 2981 1652
rect 2858 1653 2916 1654
rect 2801 1655 2859 1656
rect 2953 1655 3021 1656
rect 2909 1657 2955 1658
rect 2956 1657 3024 1658
rect 2959 1659 3015 1660
rect 2900 1661 2961 1662
rect 2962 1661 3003 1662
rect 2903 1663 2964 1664
rect 2965 1663 3027 1664
rect 2968 1665 3030 1666
rect 2971 1667 2999 1668
rect 2944 1669 3000 1670
rect 2921 1671 2946 1672
rect 2974 1671 2985 1672
rect 3004 1671 3064 1672
rect 3007 1673 3067 1674
rect 3044 1675 3056 1676
rect 3047 1677 3053 1678
rect 2533 1686 2655 1687
rect 2551 1688 2594 1689
rect 2575 1690 2664 1691
rect 2590 1692 2626 1693
rect 2605 1694 2735 1695
rect 2605 1696 2905 1697
rect 2619 1698 2774 1699
rect 2619 1700 2804 1701
rect 2612 1702 2803 1703
rect 2628 1704 2668 1705
rect 2634 1706 2680 1707
rect 2643 1708 2765 1709
rect 2660 1710 2677 1711
rect 2696 1710 2714 1711
rect 2699 1712 2708 1713
rect 2705 1714 2717 1715
rect 2730 1714 3019 1715
rect 2748 1716 2759 1717
rect 2766 1716 2780 1717
rect 2772 1718 2838 1719
rect 2770 1720 2839 1721
rect 2769 1722 2783 1723
rect 2778 1724 2792 1725
rect 2781 1726 2795 1727
rect 2784 1728 2798 1729
rect 2746 1730 2797 1731
rect 2790 1732 2807 1733
rect 2685 1734 2806 1735
rect 2684 1736 2889 1737
rect 2808 1738 2829 1739
rect 2669 1740 2830 1741
rect 2812 1742 2920 1743
rect 2811 1744 2832 1745
rect 2820 1746 2826 1747
rect 2638 1748 2827 1749
rect 2637 1750 2652 1751
rect 2622 1752 2651 1753
rect 2823 1752 2835 1753
rect 2631 1754 2836 1755
rect 2853 1754 2874 1755
rect 2855 1756 2866 1757
rect 2856 1758 2877 1759
rect 2861 1760 2902 1761
rect 2867 1762 2878 1763
rect 2858 1764 2869 1765
rect 2849 1766 2860 1767
rect 2733 1768 2851 1769
rect 2883 1768 2886 1769
rect 2894 1768 2926 1769
rect 2907 1770 2931 1771
rect 2909 1772 2968 1773
rect 2921 1774 3013 1775
rect 2931 1776 2949 1777
rect 2726 1778 2950 1779
rect 2937 1780 2946 1781
rect 2951 1780 3090 1781
rect 2952 1782 2970 1783
rect 2955 1784 2977 1785
rect 2958 1786 2961 1787
rect 2961 1788 2964 1789
rect 2973 1788 3114 1789
rect 2976 1790 3003 1791
rect 2983 1792 2991 1793
rect 2994 1792 3015 1793
rect 2927 1794 3016 1795
rect 2891 1796 2929 1797
rect 3003 1796 3098 1797
rect 3006 1798 3152 1799
rect 3020 1800 3056 1801
rect 3021 1802 3027 1803
rect 2915 1804 3028 1805
rect 3023 1806 3059 1807
rect 3029 1808 3075 1809
rect 3063 1810 3113 1811
rect 2964 1812 3065 1813
rect 3066 1812 3073 1813
rect 2912 1814 3072 1815
rect 3083 1814 3120 1815
rect 3106 1816 3110 1817
rect 2548 1825 2579 1826
rect 2552 1827 2576 1828
rect 2587 1827 2664 1828
rect 2593 1829 2600 1830
rect 2593 1831 2715 1832
rect 2605 1833 2818 1834
rect 2619 1835 2706 1836
rect 2622 1837 2626 1838
rect 2637 1837 2653 1838
rect 2634 1839 2637 1840
rect 2640 1839 2824 1840
rect 2647 1841 2866 1842
rect 2657 1843 2779 1844
rect 2664 1845 2677 1846
rect 2667 1847 2851 1848
rect 2683 1849 2797 1850
rect 2687 1851 2773 1852
rect 2615 1853 2773 1854
rect 2690 1855 2782 1856
rect 2696 1857 2718 1858
rect 2699 1859 2703 1860
rect 2723 1859 2824 1860
rect 2730 1861 2848 1862
rect 2733 1863 2893 1864
rect 2748 1865 2752 1866
rect 2766 1865 2779 1866
rect 2655 1867 2767 1868
rect 2769 1867 2782 1868
rect 2784 1867 2794 1868
rect 2790 1869 2800 1870
rect 2790 1871 2821 1872
rect 2805 1873 2833 1874
rect 2829 1875 2842 1876
rect 2802 1877 2830 1878
rect 2838 1877 2863 1878
rect 2811 1879 2839 1880
rect 2726 1881 2812 1882
rect 2847 1881 3141 1882
rect 2856 1883 2887 1884
rect 2826 1885 2857 1886
rect 2859 1885 2872 1886
rect 2835 1887 2860 1888
rect 2808 1889 2836 1890
rect 2868 1889 2875 1890
rect 2877 1889 2896 1890
rect 2877 1891 2905 1892
rect 2889 1893 2968 1894
rect 2901 1895 2911 1896
rect 2904 1897 2908 1898
rect 2883 1899 2908 1900
rect 2853 1901 2884 1902
rect 2643 1903 2854 1904
rect 2913 1903 2929 1904
rect 2916 1905 2926 1906
rect 2919 1907 2923 1908
rect 2919 1909 2950 1910
rect 2931 1911 2935 1912
rect 2937 1911 2986 1912
rect 2940 1913 2962 1914
rect 2949 1915 3016 1916
rect 2958 1917 2971 1918
rect 2955 1919 2959 1920
rect 2952 1921 2956 1922
rect 2952 1923 3019 1924
rect 2964 1925 2983 1926
rect 2967 1927 3101 1928
rect 2979 1929 3072 1930
rect 2991 1931 3013 1932
rect 2994 1933 3019 1934
rect 2994 1935 3004 1936
rect 3000 1937 3136 1938
rect 2973 1939 3001 1940
rect 3006 1939 3025 1940
rect 2976 1941 3007 1942
rect 3021 1941 3037 1942
rect 3034 1943 3065 1944
rect 3043 1945 3130 1946
rect 3046 1947 3049 1948
rect 3045 1949 3084 1950
rect 3055 1951 3067 1952
rect 3058 1953 3070 1954
rect 3074 1953 3094 1954
rect 3092 1955 3107 1956
rect 3114 1955 3155 1956
rect 3117 1957 3155 1958
rect 3126 1959 3165 1960
rect 3132 1961 3151 1962
rect 3144 1963 3148 1964
rect 3144 1965 3171 1966
rect 2596 1974 2708 1975
rect 2609 1976 2703 1977
rect 2587 1978 2610 1979
rect 2615 1978 2620 1979
rect 2619 1980 2693 1981
rect 2623 1982 2857 1983
rect 2626 1984 2720 1985
rect 2629 1986 2815 1987
rect 2633 1988 2647 1989
rect 2636 1990 2681 1991
rect 2649 1992 2767 1993
rect 2656 1994 2860 1995
rect 2658 1996 2665 1997
rect 2661 1998 2705 1999
rect 2683 2000 2875 2001
rect 2652 2002 2684 2003
rect 2642 2004 2654 2005
rect 2690 2004 2770 2005
rect 2695 2006 3142 2007
rect 2714 2008 2746 2009
rect 2717 2010 2749 2011
rect 2725 2012 2791 2013
rect 2732 2014 2893 2015
rect 2633 2016 2893 2017
rect 2772 2018 2905 2019
rect 2802 2020 2866 2021
rect 2823 2022 2860 2023
rect 2829 2024 2866 2025
rect 2647 2026 2830 2027
rect 2832 2026 2869 2027
rect 2742 2028 2833 2029
rect 2838 2028 2881 2029
rect 2886 2028 2926 2029
rect 2862 2030 2887 2031
rect 2901 2030 3082 2031
rect 2871 2032 2902 2033
rect 2847 2034 2872 2035
rect 2811 2036 2848 2037
rect 2778 2038 2812 2039
rect 2910 2038 2944 2039
rect 2913 2040 2947 2041
rect 2895 2042 2914 2043
rect 2735 2044 2896 2045
rect 2686 2046 2736 2047
rect 2605 2048 2687 2049
rect 2919 2048 2929 2049
rect 2889 2050 2920 2051
rect 2853 2052 2890 2053
rect 2817 2054 2854 2055
rect 2934 2054 2977 2055
rect 2940 2056 3016 2057
rect 2907 2058 2941 2059
rect 2877 2060 2908 2061
rect 2835 2062 2878 2063
rect 2793 2064 2836 2065
rect 2751 2066 2794 2067
rect 2751 2068 2782 2069
rect 2781 2070 2965 2071
rect 2967 2070 3004 2071
rect 2952 2072 2968 2073
rect 2979 2072 3103 2073
rect 2988 2074 3040 2075
rect 2955 2076 2989 2077
rect 2916 2078 2956 2079
rect 3000 2078 3192 2079
rect 3006 2080 3040 2081
rect 3012 2082 3085 2083
rect 3015 2084 3099 2085
rect 2982 2086 3100 2087
rect 2949 2088 2983 2089
rect 3018 2088 3196 2089
rect 2991 2090 3019 2091
rect 2958 2092 2992 2093
rect 2922 2094 2959 2095
rect 2883 2096 2923 2097
rect 2841 2098 2884 2099
rect 2799 2100 2842 2101
rect 2799 2102 2953 2103
rect 3027 2102 3121 2103
rect 3033 2104 3136 2105
rect 3036 2106 3160 2107
rect 3045 2108 3106 2109
rect 3024 2110 3046 2111
rect 3048 2110 3064 2111
rect 3075 2110 3090 2111
rect 3092 2110 3096 2111
rect 3066 2112 3094 2113
rect 3069 2114 3097 2115
rect 3114 2114 3158 2115
rect 3117 2116 3136 2117
rect 3122 2118 3157 2119
rect 3129 2120 3148 2121
rect 3132 2122 3172 2123
rect 3144 2124 3178 2125
rect 3126 2126 3145 2127
rect 3150 2126 3169 2127
rect 2994 2128 3151 2129
rect 2994 2130 3022 2131
rect 3174 2130 3185 2131
rect 3204 2130 3209 2131
rect 2594 2139 2852 2140
rect 2587 2141 2595 2142
rect 2603 2141 2854 2142
rect 2604 2143 2618 2144
rect 2619 2143 2687 2144
rect 2620 2145 2693 2146
rect 2622 2147 2696 2148
rect 2626 2149 2855 2150
rect 2633 2151 2900 2152
rect 2633 2153 2708 2154
rect 2637 2155 2752 2156
rect 2640 2157 2866 2158
rect 2643 2159 2688 2160
rect 2644 2161 2936 2162
rect 2650 2163 2822 2164
rect 2650 2165 2654 2166
rect 2653 2167 2777 2168
rect 2660 2169 2794 2170
rect 2666 2171 2869 2172
rect 2669 2173 2681 2174
rect 2672 2175 2684 2176
rect 2681 2177 2893 2178
rect 2693 2179 2705 2180
rect 2702 2181 2720 2182
rect 2733 2181 2746 2182
rect 2742 2183 2881 2184
rect 2748 2185 2755 2186
rect 2748 2187 2770 2188
rect 2794 2187 2905 2188
rect 2735 2189 2906 2190
rect 2809 2191 2812 2192
rect 2814 2191 2894 2192
rect 2827 2193 2836 2194
rect 2829 2195 2840 2196
rect 2845 2195 2848 2196
rect 2866 2195 2872 2196
rect 2872 2197 2944 2198
rect 2881 2199 2887 2200
rect 2597 2201 2888 2202
rect 2895 2201 2951 2202
rect 2889 2203 2897 2204
rect 2606 2205 2891 2206
rect 2600 2207 2608 2208
rect 2601 2209 2610 2210
rect 2610 2211 2801 2212
rect 2925 2211 2933 2212
rect 2919 2213 2927 2214
rect 2715 2215 2921 2216
rect 2928 2215 2986 2216
rect 2922 2217 2930 2218
rect 2955 2217 2963 2218
rect 2964 2217 2972 2218
rect 2958 2219 2966 2220
rect 2952 2221 2960 2222
rect 2946 2223 2954 2224
rect 2940 2225 2948 2226
rect 2967 2225 2975 2226
rect 2976 2225 3010 2226
rect 2991 2227 2999 2228
rect 3000 2227 3076 2228
rect 2994 2229 3002 2230
rect 2988 2231 2996 2232
rect 3015 2231 3116 2232
rect 3018 2233 3032 2234
rect 3027 2235 3077 2236
rect 3033 2237 3068 2238
rect 3037 2239 3216 2240
rect 3039 2241 3056 2242
rect 3045 2243 3062 2244
rect 3012 2245 3047 2246
rect 3003 2247 3014 2248
rect 3004 2249 3151 2250
rect 3063 2251 3089 2252
rect 3073 2253 3160 2254
rect 3079 2255 3258 2256
rect 3096 2257 3140 2258
rect 3105 2259 3161 2260
rect 3106 2261 3152 2262
rect 3112 2263 3179 2264
rect 3118 2265 3142 2266
rect 3081 2267 3143 2268
rect 3082 2269 3167 2270
rect 3125 2271 3164 2272
rect 3135 2273 3195 2274
rect 3093 2275 3137 2276
rect 3147 2275 3185 2276
rect 3099 2277 3149 2278
rect 3154 2277 3205 2278
rect 3156 2279 3175 2280
rect 3157 2281 3264 2282
rect 3168 2283 3228 2284
rect 3171 2285 3231 2286
rect 2612 2287 3173 2288
rect 3181 2287 3192 2288
rect 3144 2289 3182 2290
rect 3084 2291 3146 2292
rect 3201 2291 3241 2292
rect 3270 2291 3278 2292
rect 2587 2300 2608 2301
rect 2610 2300 2885 2301
rect 2611 2302 2888 2303
rect 2623 2304 2897 2305
rect 2625 2306 2840 2307
rect 2628 2308 2870 2309
rect 2633 2310 2688 2311
rect 2632 2312 2891 2313
rect 2640 2314 2816 2315
rect 2650 2316 2677 2317
rect 2656 2318 2882 2319
rect 2679 2320 2694 2321
rect 2681 2322 2849 2323
rect 2694 2324 2703 2325
rect 2718 2324 2861 2325
rect 2721 2326 2729 2327
rect 2731 2326 2734 2327
rect 2604 2328 2735 2329
rect 2757 2328 2900 2329
rect 2661 2330 2759 2331
rect 2760 2330 2789 2331
rect 2764 2332 2915 2333
rect 2782 2334 2795 2335
rect 2791 2336 3208 2337
rect 2797 2338 2927 2339
rect 2812 2340 2894 2341
rect 2833 2342 2840 2343
rect 2821 2344 2834 2345
rect 2620 2346 2822 2347
rect 2836 2346 2843 2347
rect 2851 2346 2858 2347
rect 2590 2348 2852 2349
rect 2590 2350 2713 2351
rect 2854 2350 2864 2351
rect 2593 2352 2855 2353
rect 2872 2352 2982 2353
rect 2600 2354 2873 2355
rect 2878 2354 2901 2355
rect 2666 2356 2879 2357
rect 2891 2356 2928 2357
rect 2902 2358 2919 2359
rect 2653 2360 2904 2361
rect 2630 2362 2655 2363
rect 2905 2362 2940 2363
rect 2866 2364 2907 2365
rect 2742 2366 2867 2367
rect 2743 2368 2749 2369
rect 2924 2368 3255 2369
rect 2947 2370 3179 2371
rect 2884 2372 2949 2373
rect 2962 2372 2979 2373
rect 2971 2374 3027 2375
rect 2908 2376 2973 2377
rect 2984 2376 3060 2377
rect 2987 2378 3100 2379
rect 2998 2380 3018 2381
rect 3001 2382 3048 2383
rect 3004 2384 3051 2385
rect 2965 2386 3006 2387
rect 2953 2388 2967 2389
rect 2935 2390 2955 2391
rect 2845 2392 2937 2393
rect 2635 2394 2846 2395
rect 3007 2394 3191 2395
rect 2827 2396 3190 2397
rect 2682 2398 2828 2399
rect 3013 2398 3030 2399
rect 3019 2400 3054 2401
rect 3022 2402 3044 2403
rect 2974 2404 3024 2405
rect 2920 2406 2976 2407
rect 3037 2406 3244 2407
rect 3041 2408 3198 2409
rect 3055 2410 3267 2411
rect 2995 2412 3057 2413
rect 3067 2412 3072 2413
rect 3073 2412 3087 2413
rect 3076 2414 3246 2415
rect 3077 2416 3281 2417
rect 3079 2418 3291 2419
rect 3088 2420 3103 2421
rect 2950 2422 3090 2423
rect 2794 2424 2952 2425
rect 3106 2424 3127 2425
rect 3108 2426 3185 2427
rect 3112 2428 3133 2429
rect 3120 2430 3130 2431
rect 3142 2430 3152 2431
rect 3031 2432 3142 2433
rect 3136 2434 3151 2435
rect 3115 2436 3136 2437
rect 3145 2436 3149 2437
rect 3154 2436 3188 2437
rect 3139 2438 3154 2439
rect 3138 2440 3158 2441
rect 2875 2442 3157 2443
rect 2621 2444 2876 2445
rect 3163 2444 3167 2445
rect 3082 2446 3166 2447
rect 3160 2448 3163 2449
rect 3061 2450 3160 2451
rect 3172 2450 3187 2451
rect 3183 2452 3270 2453
rect 3201 2454 3212 2455
rect 3181 2456 3211 2457
rect 3218 2456 3248 2457
rect 3227 2458 3240 2459
rect 3174 2460 3228 2461
rect 3230 2460 3243 2461
rect 2593 2469 2916 2470
rect 2600 2471 2852 2472
rect 2600 2473 2732 2474
rect 2604 2475 2849 2476
rect 2603 2477 2772 2478
rect 2607 2479 2913 2480
rect 2587 2481 2607 2482
rect 2618 2481 2850 2482
rect 2625 2483 2858 2484
rect 2630 2485 2641 2486
rect 2635 2487 2853 2488
rect 2642 2489 2898 2490
rect 2658 2491 2744 2492
rect 2661 2493 2837 2494
rect 2670 2495 2697 2496
rect 2673 2497 2706 2498
rect 2676 2499 2820 2500
rect 2679 2501 2688 2502
rect 2682 2503 2816 2504
rect 2626 2505 2817 2506
rect 2681 2507 2879 2508
rect 2694 2509 2739 2510
rect 2702 2511 2919 2512
rect 2712 2513 2733 2514
rect 2714 2515 2813 2516
rect 2726 2517 2855 2518
rect 2728 2519 3254 2520
rect 2734 2521 2775 2522
rect 2750 2523 2949 2524
rect 2776 2525 2805 2526
rect 2619 2527 2778 2528
rect 2800 2527 2910 2528
rect 2755 2529 2802 2530
rect 2581 2531 2757 2532
rect 2827 2531 2859 2532
rect 2839 2533 2883 2534
rect 2845 2535 2895 2536
rect 2809 2537 2847 2538
rect 2869 2537 2919 2538
rect 2833 2539 2871 2540
rect 2872 2539 2922 2540
rect 2758 2541 2874 2542
rect 2759 2543 2783 2544
rect 2888 2543 2967 2544
rect 2633 2545 2889 2546
rect 2900 2545 2949 2546
rect 2863 2547 2901 2548
rect 2821 2549 2865 2550
rect 2924 2549 2985 2550
rect 2875 2551 2925 2552
rect 2930 2551 2991 2552
rect 2685 2553 2931 2554
rect 2933 2553 2994 2554
rect 2936 2555 2967 2556
rect 2831 2557 2937 2558
rect 2939 2557 2970 2558
rect 2954 2559 2997 2560
rect 2623 2561 2955 2562
rect 2972 2561 3003 2562
rect 2975 2563 3012 2564
rect 2978 2565 3021 2566
rect 2951 2567 2979 2568
rect 2903 2569 2952 2570
rect 2866 2571 2904 2572
rect 2987 2571 3114 2572
rect 2927 2573 2988 2574
rect 2584 2575 2928 2576
rect 3005 2575 3036 2576
rect 2891 2577 3006 2578
rect 3017 2577 3093 2578
rect 2960 2579 3018 2580
rect 2906 2581 2961 2582
rect 2596 2583 2907 2584
rect 3023 2583 3063 2584
rect 3026 2585 3060 2586
rect 3029 2587 3084 2588
rect 3041 2589 3235 2590
rect 3044 2591 3100 2592
rect 3047 2593 3156 2594
rect 3050 2595 3180 2596
rect 2981 2597 3051 2598
rect 2753 2599 2982 2600
rect 3053 2599 3090 2600
rect 2654 2601 3054 2602
rect 3056 2601 3093 2602
rect 3056 2603 3130 2604
rect 3071 2605 3123 2606
rect 3077 2607 3288 2608
rect 3077 2609 3263 2610
rect 3086 2611 3147 2612
rect 3102 2613 3159 2614
rect 3038 2615 3102 2616
rect 3119 2615 3142 2616
rect 3126 2617 3202 2618
rect 3128 2619 3136 2620
rect 3132 2621 3214 2622
rect 3131 2623 3260 2624
rect 3134 2625 3274 2626
rect 3138 2627 3270 2628
rect 3143 2629 3291 2630
rect 3150 2631 3195 2632
rect 3149 2633 3249 2634
rect 3153 2635 3198 2636
rect 2876 2637 3153 2638
rect 3174 2637 3226 2638
rect 3204 2639 3221 2640
rect 3168 2641 3204 2642
rect 3183 2643 3220 2644
rect 3162 2645 3183 2646
rect 3207 2645 3273 2646
rect 3210 2647 3276 2648
rect 3041 2649 3211 2650
rect 3216 2649 3245 2650
rect 3223 2651 3282 2652
rect 3186 2653 3223 2654
rect 3165 2655 3186 2656
rect 3108 2657 3165 2658
rect 3228 2657 3279 2658
rect 3239 2659 3291 2660
rect 3242 2661 3294 2662
rect 3303 2661 3318 2662
rect 2584 2670 2766 2671
rect 2596 2672 2919 2673
rect 2606 2674 2614 2675
rect 2581 2676 2608 2677
rect 2609 2676 2823 2677
rect 2616 2678 2922 2679
rect 2619 2680 2715 2681
rect 2603 2682 2620 2683
rect 2623 2682 2901 2683
rect 2633 2684 2678 2685
rect 2637 2686 3117 2687
rect 2647 2688 2859 2689
rect 2654 2690 2946 2691
rect 2658 2692 2901 2693
rect 2672 2694 2967 2695
rect 2683 2696 2688 2697
rect 2681 2698 2687 2699
rect 2693 2698 2871 2699
rect 2692 2700 2697 2701
rect 2702 2700 2853 2701
rect 2705 2702 2715 2703
rect 2723 2702 2727 2703
rect 2729 2702 2733 2703
rect 2738 2702 2742 2703
rect 2747 2702 2955 2703
rect 2669 2704 2955 2705
rect 2668 2706 2973 2707
rect 2756 2708 2763 2709
rect 2768 2708 2778 2709
rect 2771 2710 2781 2711
rect 2774 2712 3297 2713
rect 2786 2714 3015 2715
rect 2789 2716 2874 2717
rect 2792 2718 2952 2719
rect 2798 2720 2802 2721
rect 2801 2722 2904 2723
rect 2600 2724 2904 2725
rect 2831 2726 2931 2727
rect 2840 2728 2847 2729
rect 2849 2728 2922 2729
rect 2849 2730 3003 2731
rect 2661 2732 3003 2733
rect 2852 2734 2865 2735
rect 2870 2734 2883 2735
rect 2876 2736 2895 2737
rect 2654 2738 2895 2739
rect 2879 2740 3006 2741
rect 2882 2742 2907 2743
rect 2885 2744 2910 2745
rect 2888 2746 2931 2747
rect 2888 2748 2913 2749
rect 2637 2750 2913 2751
rect 2891 2752 2916 2753
rect 2906 2754 2925 2755
rect 2909 2756 2928 2757
rect 2942 2756 2949 2757
rect 2951 2756 3192 2757
rect 2960 2758 3009 2759
rect 2960 2760 2985 2761
rect 2834 2762 2985 2763
rect 2966 2764 2991 2765
rect 2837 2766 2991 2767
rect 2981 2768 3048 2769
rect 2981 2770 3060 2771
rect 2993 2772 3216 2773
rect 3011 2774 3075 2775
rect 3020 2776 3174 2777
rect 3020 2778 3039 2779
rect 2996 2780 3039 2781
rect 2996 2782 3018 2783
rect 2969 2784 3018 2785
rect 2699 2786 2970 2787
rect 2698 2788 2979 2789
rect 2978 2790 2988 2791
rect 3035 2790 3108 2791
rect 3044 2792 3069 2793
rect 2750 2794 3045 2795
rect 3056 2794 3266 2795
rect 3041 2796 3057 2797
rect 3059 2796 3105 2797
rect 3083 2798 3111 2799
rect 3104 2800 3177 2801
rect 2936 2802 3177 2803
rect 3125 2804 3156 2805
rect 3119 2806 3156 2807
rect 3128 2808 3263 2809
rect 3134 2810 3331 2811
rect 3137 2812 3207 2813
rect 3143 2814 3171 2815
rect 3131 2816 3144 2817
rect 3149 2816 3189 2817
rect 3089 2818 3150 2819
rect 3158 2818 3235 2819
rect 3182 2820 3241 2821
rect 3194 2822 3318 2823
rect 3053 2824 3195 2825
rect 2759 2826 3054 2827
rect 2644 2828 2760 2829
rect 2644 2830 2919 2831
rect 3197 2830 3315 2831
rect 3164 2832 3198 2833
rect 3122 2834 3165 2835
rect 3203 2834 3235 2835
rect 3225 2836 3279 2837
rect 3228 2838 3282 2839
rect 3231 2840 3269 2841
rect 3238 2842 3247 2843
rect 3152 2844 3238 2845
rect 3092 2846 3153 2847
rect 3092 2848 3325 2849
rect 3244 2850 3382 2851
rect 3185 2852 3244 2853
rect 3146 2854 3186 2855
rect 3077 2856 3147 2857
rect 3253 2856 3309 2857
rect 3252 2858 3340 2859
rect 3272 2860 3334 2861
rect 3210 2862 3273 2863
rect 3275 2862 3337 2863
rect 3290 2864 3359 2865
rect 3219 2866 3291 2867
rect 3293 2866 3362 2867
rect 3222 2868 3294 2869
rect 3113 2870 3223 2871
rect 3050 2872 3114 2873
rect 2846 2874 3051 2875
rect 3299 2874 3304 2875
rect 3388 2874 3396 2875
rect 2539 2883 2547 2884
rect 2588 2883 2766 2884
rect 2591 2885 2889 2886
rect 2590 2887 2763 2888
rect 2598 2889 2933 2890
rect 2602 2891 2762 2892
rect 2605 2893 2608 2894
rect 2608 2895 2614 2896
rect 2611 2897 2720 2898
rect 2623 2899 2892 2900
rect 2630 2901 2910 2902
rect 2640 2903 2738 2904
rect 2644 2905 2913 2906
rect 2644 2907 2760 2908
rect 2651 2909 2867 2910
rect 2647 2911 2652 2912
rect 2647 2913 2873 2914
rect 2654 2915 2877 2916
rect 2658 2917 2853 2918
rect 2658 2919 2975 2920
rect 2661 2921 2915 2922
rect 2661 2923 2742 2924
rect 2665 2925 2898 2926
rect 2673 2927 2895 2928
rect 2677 2929 2912 2930
rect 2683 2931 2689 2932
rect 2682 2933 2687 2934
rect 2692 2933 2695 2934
rect 2575 2935 2692 2936
rect 2698 2935 2936 2936
rect 2700 2937 2927 2938
rect 2702 2939 2970 2940
rect 2710 2941 2715 2942
rect 2723 2941 2735 2942
rect 2729 2943 2732 2944
rect 2747 2943 2979 2944
rect 2750 2945 2802 2946
rect 2768 2947 2786 2948
rect 2767 2949 2904 2950
rect 2773 2951 2781 2952
rect 2792 2951 2801 2952
rect 2791 2953 2799 2954
rect 2804 2953 2837 2954
rect 2806 2955 2817 2956
rect 2812 2957 2823 2958
rect 2819 2959 2822 2960
rect 2752 2961 2819 2962
rect 2830 2961 2841 2962
rect 2834 2963 3003 2964
rect 2870 2965 2876 2966
rect 2878 2965 2931 2966
rect 2882 2967 2891 2968
rect 2885 2969 2894 2970
rect 2884 2971 2919 2972
rect 2887 2973 2922 2974
rect 2900 2975 2903 2976
rect 2906 2975 2909 2976
rect 2616 2977 2906 2978
rect 2920 2977 2943 2978
rect 2923 2979 2946 2980
rect 2941 2981 3009 2982
rect 2947 2983 3015 2984
rect 2951 2985 3008 2986
rect 2966 2987 2978 2988
rect 2960 2989 2966 2990
rect 2954 2991 2960 2992
rect 2984 2991 3269 2992
rect 2848 2993 2984 2994
rect 2992 2993 3018 2994
rect 2996 2995 3014 2996
rect 2990 2997 2996 2998
rect 2749 2999 2990 3000
rect 3020 2999 3032 3000
rect 3019 3001 3045 3002
rect 3022 3003 3048 3004
rect 3025 3005 3051 3006
rect 3028 3007 3054 3008
rect 3038 3009 3095 3010
rect 3037 3011 3117 3012
rect 3043 3013 3266 3014
rect 3056 3015 3065 3016
rect 3055 3017 3365 3018
rect 3059 3019 3226 3020
rect 3061 3021 3216 3022
rect 3074 3023 3077 3024
rect 3079 3023 3368 3024
rect 3085 3025 3108 3026
rect 3104 3027 3122 3028
rect 3092 3029 3104 3030
rect 3091 3031 3174 3032
rect 3125 3033 3340 3034
rect 3124 3035 3209 3036
rect 3133 3037 3150 3038
rect 3137 3039 3140 3040
rect 3136 3041 3153 3042
rect 3146 3043 3325 3044
rect 3143 3045 3146 3046
rect 3148 3045 3322 3046
rect 3155 3047 3343 3048
rect 3164 3049 3167 3050
rect 3163 3051 3331 3052
rect 3170 3053 3408 3054
rect 3172 3055 3195 3056
rect 3176 3057 3207 3058
rect 3113 3059 3176 3060
rect 3202 3059 3244 3060
rect 3218 3061 3223 3062
rect 3157 3063 3223 3064
rect 3232 3063 3284 3064
rect 3234 3065 3262 3066
rect 3235 3067 3318 3068
rect 3237 3069 3259 3070
rect 3110 3071 3239 3072
rect 3252 3071 3299 3072
rect 3259 3073 3320 3074
rect 3265 3075 3332 3076
rect 3286 3077 3315 3078
rect 3290 3079 3314 3080
rect 3278 3081 3290 3082
rect 3272 3083 3278 3084
rect 3293 3083 3303 3084
rect 3292 3085 3356 3086
rect 3295 3087 3337 3088
rect 3305 3089 3317 3090
rect 3308 3091 3326 3092
rect 3281 3093 3308 3094
rect 3240 3095 3281 3096
rect 3327 3095 3371 3096
rect 3333 3097 3386 3098
rect 3358 3099 3365 3100
rect 3361 3101 3368 3102
rect 3374 3101 3385 3102
rect 3381 3103 3395 3104
rect 3391 3105 3399 3106
rect 2578 3114 2600 3115
rect 2582 3116 2692 3117
rect 2587 3118 2666 3119
rect 2589 3120 2778 3121
rect 2596 3122 2894 3123
rect 2602 3124 2612 3125
rect 2605 3126 2669 3127
rect 2608 3128 2617 3129
rect 2610 3130 2856 3131
rect 2613 3132 2885 3133
rect 2623 3134 2813 3135
rect 2603 3136 2814 3137
rect 2626 3138 2826 3139
rect 2631 3140 2768 3141
rect 2640 3142 2888 3143
rect 2645 3144 2952 3145
rect 2662 3146 2886 3147
rect 2677 3148 2906 3149
rect 2686 3150 2883 3151
rect 2688 3152 2705 3153
rect 2700 3154 2915 3155
rect 2694 3156 2702 3157
rect 2682 3158 2696 3159
rect 2683 3160 3032 3161
rect 2707 3162 2784 3163
rect 2707 3164 2879 3165
rect 2710 3166 2727 3167
rect 2714 3168 3012 3169
rect 2719 3170 2742 3171
rect 2737 3172 2841 3173
rect 2734 3174 2739 3175
rect 2731 3176 2736 3177
rect 2752 3176 3023 3177
rect 2761 3178 2769 3179
rect 2765 3180 2792 3181
rect 2773 3182 2796 3183
rect 2527 3184 2775 3185
rect 2785 3184 2790 3185
rect 2786 3186 2924 3187
rect 2800 3188 2907 3189
rect 2804 3190 2964 3191
rect 2818 3192 2847 3193
rect 2647 3194 2820 3195
rect 2633 3196 2649 3197
rect 2821 3196 2889 3197
rect 2641 3198 2823 3199
rect 2828 3198 2912 3199
rect 2836 3200 2865 3201
rect 2830 3202 2838 3203
rect 2806 3204 2832 3205
rect 2843 3204 2891 3205
rect 2848 3206 2948 3207
rect 2852 3208 2903 3209
rect 2866 3210 2871 3211
rect 2872 3210 2880 3211
rect 2897 3210 3008 3211
rect 2903 3212 2921 3213
rect 2908 3214 3371 3215
rect 2909 3216 2960 3217
rect 2915 3218 2966 3219
rect 2921 3220 2978 3221
rect 2930 3222 2981 3223
rect 2658 3224 2982 3225
rect 2652 3226 2660 3227
rect 2935 3226 3042 3227
rect 2939 3228 2972 3229
rect 2941 3230 2979 3231
rect 2954 3232 2975 3233
rect 2957 3234 3014 3235
rect 2975 3236 2993 3237
rect 2983 3238 2988 3239
rect 2993 3238 3020 3239
rect 2999 3240 3044 3241
rect 3023 3242 3026 3243
rect 3028 3242 3051 3243
rect 3029 3244 3038 3245
rect 3035 3246 3068 3247
rect 3047 3248 3156 3249
rect 3055 3250 3311 3251
rect 3059 3252 3062 3253
rect 3064 3252 3216 3253
rect 3073 3254 3194 3255
rect 3077 3256 3134 3257
rect 3079 3258 3353 3259
rect 3080 3260 3137 3261
rect 3083 3262 3233 3263
rect 3094 3264 3108 3265
rect 3095 3266 3226 3267
rect 3098 3268 3158 3269
rect 3103 3270 3272 3271
rect 3091 3272 3105 3273
rect 3092 3274 3146 3275
rect 3121 3276 3209 3277
rect 3122 3278 3185 3279
rect 3128 3280 3173 3281
rect 3131 3282 3176 3283
rect 3134 3284 3197 3285
rect 3146 3286 3196 3287
rect 3148 3288 3349 3289
rect 3124 3290 3150 3291
rect 3125 3292 3188 3293
rect 3152 3294 3260 3295
rect 3163 3296 3374 3297
rect 3085 3298 3163 3299
rect 3086 3300 3140 3301
rect 3140 3302 3203 3303
rect 3168 3304 3239 3305
rect 3177 3306 3385 3307
rect 3186 3308 3248 3309
rect 3190 3310 3257 3311
rect 3216 3312 3278 3313
rect 3219 3314 3281 3315
rect 3229 3316 3308 3317
rect 3238 3318 3299 3319
rect 3241 3320 3290 3321
rect 3253 3322 3260 3323
rect 3262 3322 3314 3323
rect 3265 3324 3323 3325
rect 3265 3326 3326 3327
rect 2875 3328 3325 3329
rect 2876 3330 2933 3331
rect 2933 3332 2990 3333
rect 3304 3332 3365 3333
rect 3307 3334 3368 3335
rect 3310 3336 3332 3337
rect 3316 3338 3381 3339
rect 3166 3340 3318 3341
rect 3165 3342 3236 3343
rect 3235 3344 3296 3345
rect 3244 3346 3296 3347
rect 2588 3355 2750 3356
rect 2602 3357 2628 3358
rect 2609 3359 2877 3360
rect 2631 3361 2826 3362
rect 2634 3363 2949 3364
rect 2616 3365 2634 3366
rect 2638 3365 2699 3366
rect 2648 3367 2792 3368
rect 2652 3369 2880 3370
rect 2659 3371 2907 3372
rect 2658 3373 2790 3374
rect 2662 3375 2925 3376
rect 2665 3377 2681 3378
rect 2668 3379 2684 3380
rect 2674 3381 2723 3382
rect 2677 3383 2693 3384
rect 2686 3385 2910 3386
rect 2701 3387 2717 3388
rect 2710 3389 2919 3390
rect 2695 3391 2711 3392
rect 2719 3391 2732 3392
rect 2735 3391 2747 3392
rect 2734 3393 3027 3394
rect 2765 3395 2810 3396
rect 2770 3397 2829 3398
rect 2777 3399 2798 3400
rect 2779 3401 2876 3402
rect 2783 3403 2928 3404
rect 2782 3405 2858 3406
rect 2786 3407 3018 3408
rect 2768 3409 2786 3410
rect 2741 3411 2768 3412
rect 2738 3413 2741 3414
rect 2737 3415 2760 3416
rect 2726 3417 2759 3418
rect 2795 3417 2828 3418
rect 2704 3419 2795 3420
rect 2803 3419 2994 3420
rect 2815 3421 2976 3422
rect 2831 3423 2834 3424
rect 2840 3423 2873 3424
rect 2839 3425 2847 3426
rect 2813 3427 2846 3428
rect 2852 3427 2913 3428
rect 2819 3429 2852 3430
rect 2774 3431 2819 3432
rect 2885 3431 2937 3432
rect 2897 3433 3021 3434
rect 2900 3435 2988 3436
rect 2843 3437 2901 3438
rect 2903 3437 2961 3438
rect 2595 3439 2904 3440
rect 2915 3439 2991 3440
rect 2855 3441 2916 3442
rect 2822 3443 2855 3444
rect 2933 3443 3015 3444
rect 2882 3445 2934 3446
rect 2942 3445 2952 3446
rect 2954 3445 2994 3446
rect 2613 3447 2955 3448
rect 2957 3447 3033 3448
rect 2585 3449 2958 3450
rect 2963 3449 3060 3450
rect 2864 3451 2964 3452
rect 2966 3451 3063 3452
rect 2978 3453 2985 3454
rect 2939 3455 2979 3456
rect 2888 3457 2940 3458
rect 2999 3457 3196 3458
rect 2930 3459 3000 3460
rect 2870 3461 2931 3462
rect 2837 3463 2870 3464
rect 3008 3463 3024 3464
rect 2996 3465 3024 3466
rect 2921 3467 2997 3468
rect 3011 3467 3063 3468
rect 3029 3469 3156 3470
rect 3041 3471 3072 3472
rect 3047 3473 3069 3474
rect 3050 3475 3233 3476
rect 2981 3477 3051 3478
rect 3083 3477 3117 3478
rect 3086 3479 3180 3480
rect 3086 3481 3163 3482
rect 3095 3483 3156 3484
rect 3098 3485 3120 3486
rect 3125 3485 3332 3486
rect 3092 3487 3126 3488
rect 3134 3487 3270 3488
rect 3140 3489 3171 3490
rect 3146 3491 3183 3492
rect 3104 3493 3147 3494
rect 3077 3495 3105 3496
rect 3152 3495 3328 3496
rect 3165 3497 3207 3498
rect 3128 3499 3165 3500
rect 3128 3501 3346 3502
rect 3168 3503 3210 3504
rect 3131 3505 3168 3506
rect 3177 3505 3225 3506
rect 3122 3507 3177 3508
rect 3188 3507 3193 3508
rect 3044 3509 3192 3510
rect 3216 3509 3273 3510
rect 3238 3511 3335 3512
rect 3241 3513 3279 3514
rect 3244 3515 3282 3516
rect 3253 3517 3292 3518
rect 3259 3519 3313 3520
rect 3256 3521 3261 3522
rect 3257 3523 3275 3524
rect 3219 3525 3276 3526
rect 3186 3527 3219 3528
rect 3149 3529 3186 3530
rect 3107 3531 3150 3532
rect 3080 3533 3108 3534
rect 3035 3535 3081 3536
rect 3263 3535 3371 3536
rect 3265 3537 3319 3538
rect 3235 3539 3267 3540
rect 3304 3539 3358 3540
rect 3239 3541 3306 3542
rect 3307 3541 3361 3542
rect 3373 3541 3378 3542
rect 2530 3550 2762 3551
rect 2541 3552 2678 3553
rect 2561 3554 2643 3555
rect 2564 3556 2576 3557
rect 2581 3556 2681 3557
rect 2584 3558 2687 3559
rect 2588 3560 2684 3561
rect 2595 3562 3171 3563
rect 2594 3564 2901 3565
rect 2605 3566 2916 3567
rect 2604 3568 2837 3569
rect 2609 3570 2699 3571
rect 2608 3572 2864 3573
rect 2612 3574 2955 3575
rect 2615 3576 2637 3577
rect 2639 3576 2768 3577
rect 2633 3578 2640 3579
rect 2648 3578 2843 3579
rect 2651 3580 2852 3581
rect 2652 3582 2888 3583
rect 2667 3584 2934 3585
rect 2667 3586 2891 3587
rect 2670 3588 2726 3589
rect 2671 3590 2925 3591
rect 2674 3592 2741 3593
rect 2674 3594 2931 3595
rect 2692 3596 2699 3597
rect 2695 3598 2717 3599
rect 2658 3600 2717 3601
rect 2710 3602 2723 3603
rect 2719 3604 2732 3605
rect 2734 3604 2949 3605
rect 2734 3606 2771 3607
rect 2737 3608 2768 3609
rect 2740 3610 2747 3611
rect 2743 3612 2750 3613
rect 2758 3612 2765 3613
rect 2758 3614 2810 3615
rect 2773 3616 2819 3617
rect 2655 3618 2819 3619
rect 2776 3620 2792 3621
rect 2779 3622 2795 3623
rect 2782 3624 3000 3625
rect 2782 3626 2786 3627
rect 2788 3626 2798 3627
rect 2797 3628 3240 3629
rect 2806 3630 2979 3631
rect 2806 3632 2828 3633
rect 2812 3634 3015 3635
rect 2636 3636 2813 3637
rect 2824 3636 2846 3637
rect 2833 3638 2909 3639
rect 2845 3640 2855 3641
rect 2854 3642 2913 3643
rect 2857 3644 3005 3645
rect 2627 3646 2858 3647
rect 2860 3646 2958 3647
rect 2866 3648 2870 3649
rect 2869 3650 2873 3651
rect 2875 3650 3002 3651
rect 2875 3652 3018 3653
rect 2878 3654 2937 3655
rect 2884 3656 3285 3657
rect 2894 3658 3027 3659
rect 2897 3660 3213 3661
rect 2839 3662 2897 3663
rect 2839 3664 2904 3665
rect 2902 3666 2961 3667
rect 2911 3668 2940 3669
rect 2914 3670 2997 3671
rect 2918 3672 3189 3673
rect 2920 3674 2991 3675
rect 2932 3676 2967 3677
rect 2938 3678 3024 3679
rect 2815 3680 3023 3681
rect 2942 3682 2948 3683
rect 2941 3684 3033 3685
rect 2953 3686 2985 3687
rect 2959 3688 3045 3689
rect 2963 3690 2996 3691
rect 2971 3692 3051 3693
rect 2983 3694 3063 3695
rect 2993 3696 3026 3697
rect 2872 3698 2993 3699
rect 2998 3698 3172 3699
rect 3008 3700 3060 3701
rect 3020 3702 3035 3703
rect 3044 3702 3186 3703
rect 3047 3704 3210 3705
rect 3053 3706 3129 3707
rect 3071 3708 3111 3709
rect 3071 3710 3120 3711
rect 3077 3712 3156 3713
rect 3086 3714 3156 3715
rect 3095 3716 3150 3717
rect 3095 3718 3153 3719
rect 3098 3720 3284 3721
rect 3101 3722 3105 3723
rect 3080 3724 3105 3725
rect 3107 3724 3231 3725
rect 3068 3726 3108 3727
rect 3116 3726 3288 3727
rect 3119 3728 3177 3729
rect 2989 3730 3176 3731
rect 3125 3732 3325 3733
rect 3137 3734 3328 3735
rect 3140 3736 3147 3737
rect 3146 3738 3165 3739
rect 3143 3740 3165 3741
rect 3149 3742 3168 3743
rect 3007 3744 3169 3745
rect 3152 3746 3183 3747
rect 3158 3748 3225 3749
rect 3179 3750 3349 3751
rect 3178 3752 3292 3753
rect 3182 3754 3279 3755
rect 3188 3756 3276 3757
rect 3194 3758 3282 3759
rect 3083 3760 3281 3761
rect 3197 3762 3273 3763
rect 3206 3764 3378 3765
rect 3209 3766 3335 3767
rect 3212 3768 3267 3769
rect 3218 3770 3364 3771
rect 3218 3772 3253 3773
rect 3221 3774 3270 3775
rect 3050 3776 3270 3777
rect 3234 3778 3319 3779
rect 3246 3780 3298 3781
rect 3249 3782 3295 3783
rect 3257 3784 3309 3785
rect 3260 3786 3306 3787
rect 3215 3788 3260 3789
rect 3263 3788 3330 3789
rect 3306 3790 3358 3791
rect 3309 3792 3361 3793
rect 3319 3794 3367 3795
rect 2527 3803 3093 3804
rect 2534 3805 2762 3806
rect 2545 3807 2635 3808
rect 2551 3809 2678 3810
rect 2554 3811 2643 3812
rect 2578 3813 2588 3814
rect 2581 3815 2610 3816
rect 2591 3817 2691 3818
rect 2602 3819 2858 3820
rect 2604 3821 2855 3822
rect 2615 3823 2632 3824
rect 2621 3825 2679 3826
rect 2628 3827 2813 3828
rect 2637 3829 2825 3830
rect 2639 3831 2651 3832
rect 2648 3833 2819 3834
rect 2652 3835 2937 3836
rect 2653 3837 2656 3838
rect 2664 3837 2897 3838
rect 2667 3839 2909 3840
rect 2594 3841 2910 3842
rect 2671 3843 2976 3844
rect 2686 3845 2703 3846
rect 2695 3847 2712 3848
rect 2705 3849 2717 3850
rect 2708 3851 2720 3852
rect 2722 3851 2739 3852
rect 2734 3853 3012 3854
rect 2740 3855 2751 3856
rect 2725 3857 2742 3858
rect 2743 3857 2754 3858
rect 2758 3857 2814 3858
rect 2759 3859 2921 3860
rect 2720 3861 2922 3862
rect 2762 3863 2765 3864
rect 2773 3863 2829 3864
rect 2779 3865 2799 3866
rect 2788 3867 2802 3868
rect 2782 3869 2790 3870
rect 2783 3871 2999 3872
rect 2794 3873 2933 3874
rect 2776 3875 2796 3876
rect 2806 3875 2832 3876
rect 2816 3877 2988 3878
rect 2839 3879 2895 3880
rect 2842 3881 2856 3882
rect 2843 3883 2996 3884
rect 2845 3885 2859 3886
rect 2863 3885 2919 3886
rect 2866 3887 2898 3888
rect 2867 3889 3002 3890
rect 2869 3891 2901 3892
rect 2875 3893 2990 3894
rect 2878 3895 2928 3896
rect 2756 3897 2880 3898
rect 2884 3897 2934 3898
rect 2885 3899 3114 3900
rect 2902 3901 2952 3902
rect 2723 3903 2904 3904
rect 2911 3903 2931 3904
rect 2698 3905 2913 3906
rect 2914 3905 2970 3906
rect 2860 3907 2916 3908
rect 2861 3909 2888 3910
rect 2941 3909 3000 3910
rect 2945 3911 3035 3912
rect 2947 3913 2958 3914
rect 2953 3915 2982 3916
rect 2954 3917 3162 3918
rect 2959 3919 3126 3920
rect 2971 3921 3018 3922
rect 2972 3923 3005 3924
rect 2978 3925 3026 3926
rect 3005 3927 3045 3928
rect 3029 3929 3108 3930
rect 3032 3931 3111 3932
rect 3041 3933 3060 3934
rect 3041 3935 3144 3936
rect 2770 3937 3144 3938
rect 2771 3939 3310 3940
rect 3050 3941 3087 3942
rect 3062 3943 3242 3944
rect 3071 3945 3114 3946
rect 3074 3947 3141 3948
rect 3077 3949 3141 3950
rect 3044 3951 3078 3952
rect 3080 3951 3102 3952
rect 3095 3953 3281 3954
rect 3098 3955 3281 3956
rect 3098 3957 3147 3958
rect 3047 3959 3147 3960
rect 3122 3961 3156 3962
rect 3137 3963 3263 3964
rect 3083 3965 3138 3966
rect 3083 3967 3105 3968
rect 3149 3967 3165 3968
rect 3155 3969 3260 3970
rect 3068 3971 3260 3972
rect 3164 3973 3263 3974
rect 3168 3975 3257 3976
rect 3191 3977 3198 3978
rect 3194 3979 3225 3980
rect 3188 3981 3195 3982
rect 3197 3981 3316 3982
rect 3206 3983 3219 3984
rect 3212 3985 3219 3986
rect 3209 3987 3213 3988
rect 3158 3989 3210 3990
rect 2938 3991 3159 3992
rect 2939 3993 3023 3994
rect 2983 3995 3024 3996
rect 2984 3997 2993 3998
rect 3215 3997 3253 3998
rect 3215 3999 3267 4000
rect 3221 4001 3288 4002
rect 3119 4003 3288 4004
rect 3119 4005 3153 4006
rect 3234 4005 3303 4006
rect 3246 4007 3254 4008
rect 3249 4009 3320 4010
rect 3293 4011 3307 4012
rect 3053 4013 3307 4014
rect 3007 4015 3054 4016
rect 3296 4015 3323 4016
rect 2555 4024 2571 4025
rect 2567 4026 2635 4027
rect 2576 4028 2852 4029
rect 2579 4030 2587 4031
rect 2588 4030 2596 4031
rect 2589 4032 2691 4033
rect 2593 4034 2892 4035
rect 2581 4036 2891 4037
rect 2603 4038 2802 4039
rect 2612 4040 2673 4041
rect 2619 4042 2945 4043
rect 2622 4044 2832 4045
rect 2624 4046 2742 4047
rect 2626 4048 2735 4049
rect 2640 4050 2913 4051
rect 2636 4052 2912 4053
rect 2644 4054 2985 4055
rect 2653 4056 2709 4057
rect 2678 4058 2831 4059
rect 2688 4060 2792 4061
rect 2697 4062 2706 4063
rect 2700 4064 2712 4065
rect 2720 4064 2960 4065
rect 2722 4066 3008 4067
rect 2728 4068 2739 4069
rect 2740 4068 2751 4069
rect 2743 4070 2754 4071
rect 2746 4072 2763 4073
rect 2749 4074 2868 4075
rect 2759 4076 3294 4077
rect 2767 4078 2955 4079
rect 2771 4080 2982 4081
rect 2773 4082 2784 4083
rect 2785 4082 2796 4083
rect 2806 4082 2817 4083
rect 2818 4082 2829 4083
rect 2605 4084 2828 4085
rect 2839 4084 2856 4085
rect 2843 4086 3185 4087
rect 2842 4088 2859 4089
rect 2845 4090 2862 4091
rect 2854 4092 2940 4093
rect 2860 4094 2919 4095
rect 2789 4096 2918 4097
rect 2788 4098 2799 4099
rect 2797 4100 2814 4101
rect 2812 4102 2838 4103
rect 2866 4102 2880 4103
rect 2596 4104 2879 4105
rect 2872 4106 2886 4107
rect 2584 4108 2885 4109
rect 2881 4110 2895 4111
rect 2702 4112 2894 4113
rect 2921 4112 2939 4113
rect 2678 4114 2921 4115
rect 2965 4114 2993 4115
rect 2975 4116 2981 4117
rect 2969 4118 2975 4119
rect 2957 4120 2969 4121
rect 2951 4122 2957 4123
rect 2978 4122 2984 4123
rect 2972 4124 2978 4125
rect 2987 4124 3033 4125
rect 2948 4126 2987 4127
rect 2936 4128 2948 4129
rect 2990 4128 3030 4129
rect 2999 4130 3002 4131
rect 3005 4130 3041 4131
rect 3017 4132 3020 4133
rect 3023 4132 3059 4133
rect 3025 4134 3182 4135
rect 3037 4136 3126 4137
rect 3049 4138 3099 4139
rect 3053 4140 3131 4141
rect 3052 4142 3158 4143
rect 3055 4144 3120 4145
rect 3074 4146 3333 4147
rect 3068 4148 3074 4149
rect 3062 4150 3068 4151
rect 3061 4152 3084 4153
rect 3080 4154 3104 4155
rect 3086 4156 3110 4157
rect 3092 4158 3228 4159
rect 3106 4160 3168 4161
rect 3113 4162 3204 4163
rect 3115 4164 3153 4165
rect 3118 4166 3189 4167
rect 3122 4168 3242 4169
rect 3137 4170 3303 4171
rect 3146 4172 3167 4173
rect 3155 4174 3261 4175
rect 3164 4176 3321 4177
rect 3143 4178 3164 4179
rect 3169 4178 3286 4179
rect 3194 4180 3201 4181
rect 3194 4182 3277 4183
rect 3209 4184 3237 4185
rect 2715 4186 3210 4187
rect 3212 4186 3249 4187
rect 3212 4188 3216 4189
rect 3218 4188 3252 4189
rect 3221 4190 3270 4191
rect 3127 4192 3222 4193
rect 3224 4192 3231 4193
rect 3197 4194 3225 4195
rect 3140 4196 3198 4197
rect 3077 4198 3140 4199
rect 3233 4198 3310 4199
rect 3244 4200 3254 4201
rect 3254 4202 3317 4203
rect 3245 4204 3317 4205
rect 3256 4206 3307 4207
rect 3191 4208 3258 4209
rect 3290 4208 3314 4209
rect 3296 4210 3300 4211
rect 2557 4219 2571 4220
rect 2560 4221 2565 4222
rect 2567 4221 2577 4222
rect 2582 4221 2731 4222
rect 2586 4223 2707 4224
rect 2594 4225 2882 4226
rect 2600 4227 2918 4228
rect 2612 4229 2683 4230
rect 2619 4231 2891 4232
rect 2622 4233 2852 4234
rect 2622 4235 2861 4236
rect 2626 4237 2716 4238
rect 2633 4239 2921 4240
rect 2632 4241 2948 4242
rect 2636 4243 2735 4244
rect 2636 4245 2741 4246
rect 2639 4247 3014 4248
rect 2643 4249 2972 4250
rect 2646 4251 2822 4252
rect 2648 4253 2846 4254
rect 2651 4255 2668 4256
rect 2672 4255 2689 4256
rect 2673 4257 2719 4258
rect 2694 4259 2852 4260
rect 2697 4261 2849 4262
rect 2709 4263 2744 4264
rect 2728 4265 2765 4266
rect 2746 4267 2801 4268
rect 2746 4269 3119 4270
rect 2749 4271 2996 4272
rect 2700 4273 2750 4274
rect 2752 4273 2993 4274
rect 2603 4275 2993 4276
rect 2604 4277 2609 4278
rect 2767 4277 2777 4278
rect 2797 4277 2858 4278
rect 2803 4279 2807 4280
rect 2812 4279 2861 4280
rect 2812 4281 2906 4282
rect 2815 4283 2855 4284
rect 2830 4285 2870 4286
rect 2788 4287 2831 4288
rect 2773 4289 2789 4290
rect 2845 4289 2966 4290
rect 2743 4291 2966 4292
rect 2872 4293 3017 4294
rect 2818 4295 2873 4296
rect 2887 4295 2903 4296
rect 2893 4297 2963 4298
rect 2839 4299 2894 4300
rect 2791 4301 2840 4302
rect 2899 4301 2918 4302
rect 2899 4303 2939 4304
rect 2908 4305 2948 4306
rect 2866 4307 2909 4308
rect 2827 4309 2867 4310
rect 2785 4311 2828 4312
rect 2914 4311 2990 4312
rect 2896 4313 2915 4314
rect 2926 4313 2954 4314
rect 2941 4315 2969 4316
rect 2950 4317 2999 4318
rect 2911 4319 2951 4320
rect 2956 4319 3301 4320
rect 2929 4321 2957 4322
rect 2794 4323 2930 4324
rect 2959 4323 2987 4324
rect 2884 4325 2960 4326
rect 2980 4325 3032 4326
rect 2983 4327 3035 4328
rect 2727 4329 2984 4330
rect 3001 4329 3077 4330
rect 2944 4331 3002 4332
rect 3010 4331 3023 4332
rect 3019 4333 3083 4334
rect 3007 4335 3020 4336
rect 3025 4335 3089 4336
rect 3037 4337 3080 4338
rect 3040 4339 3140 4340
rect 3043 4341 3158 4342
rect 3055 4343 3092 4344
rect 3052 4345 3056 4346
rect 2977 4347 3053 4348
rect 2932 4349 2978 4350
rect 2878 4351 2933 4352
rect 3058 4351 3185 4352
rect 3049 4353 3059 4354
rect 2974 4355 3050 4356
rect 2842 4357 2975 4358
rect 3061 4357 3095 4358
rect 3067 4359 3140 4360
rect 3064 4361 3068 4362
rect 3073 4361 3279 4362
rect 3073 4363 3116 4364
rect 3103 4365 3122 4366
rect 3106 4367 3125 4368
rect 3106 4369 3207 4370
rect 3109 4371 3158 4372
rect 3118 4373 3258 4374
rect 3127 4375 3185 4376
rect 3127 4377 3268 4378
rect 3133 4379 3282 4380
rect 3166 4381 3206 4382
rect 3169 4383 3327 4384
rect 3181 4385 3222 4386
rect 3212 4387 3219 4388
rect 2809 4389 3218 4390
rect 3224 4389 3261 4390
rect 3227 4391 3264 4392
rect 3200 4393 3227 4394
rect 3230 4393 3267 4394
rect 3203 4395 3230 4396
rect 3163 4397 3203 4398
rect 3233 4397 3270 4398
rect 3194 4399 3233 4400
rect 3193 4401 3371 4402
rect 3236 4403 3292 4404
rect 3197 4405 3236 4406
rect 3248 4405 3316 4406
rect 3112 4407 3249 4408
rect 3254 4407 3307 4408
rect 3191 4409 3255 4410
rect 3294 4409 3330 4410
rect 3302 4411 3320 4412
rect 3251 4413 3304 4414
rect 3245 4415 3252 4416
rect 3130 4417 3246 4418
rect 3309 4417 3348 4418
rect 3309 4419 3344 4420
rect 3356 4419 3368 4420
rect 2539 4428 2750 4429
rect 2588 4430 2900 4431
rect 2590 4432 2960 4433
rect 2602 4434 2779 4435
rect 2611 4436 2616 4437
rect 2612 4438 2948 4439
rect 2622 4440 2683 4441
rect 2632 4442 2909 4443
rect 2594 4444 2908 4445
rect 2595 4446 2707 4447
rect 2636 4448 2926 4449
rect 2638 4450 2954 4451
rect 2643 4452 2861 4453
rect 2649 4454 3053 4455
rect 2656 4456 2836 4457
rect 2659 4458 2849 4459
rect 2662 4460 2668 4461
rect 2665 4462 2710 4463
rect 2680 4464 2984 4465
rect 2686 4466 2951 4467
rect 2697 4468 2822 4469
rect 2707 4470 2731 4471
rect 2710 4472 2963 4473
rect 2728 4474 2736 4475
rect 2739 4474 2942 4475
rect 2739 4476 2999 4477
rect 2757 4478 2801 4479
rect 2766 4480 2777 4481
rect 2784 4480 2828 4481
rect 2788 4482 2791 4483
rect 2787 4484 2831 4485
rect 2794 4486 2806 4487
rect 2796 4488 2858 4489
rect 2799 4490 2993 4491
rect 2812 4492 2890 4493
rect 2803 4494 2812 4495
rect 2817 4494 2873 4495
rect 2820 4496 2840 4497
rect 2823 4498 2957 4499
rect 2618 4500 2956 4501
rect 2619 4502 2765 4503
rect 2826 4502 2867 4503
rect 2832 4504 2846 4505
rect 2815 4506 2845 4507
rect 2838 4508 2852 4509
rect 2850 4510 2894 4511
rect 2609 4512 2893 4513
rect 2862 4514 2888 4515
rect 2869 4516 2896 4517
rect 2629 4518 2869 4519
rect 2628 4520 2689 4521
rect 2689 4522 2915 4523
rect 2871 4524 2918 4525
rect 2874 4526 2933 4527
rect 2886 4528 2906 4529
rect 2598 4530 2905 4531
rect 2910 4530 2978 4531
rect 2916 4532 2972 4533
rect 2919 4534 2975 4535
rect 2922 4536 2990 4537
rect 2646 4538 2989 4539
rect 2645 4540 2935 4541
rect 2929 4542 3130 4543
rect 2940 4544 2996 4545
rect 2943 4546 3002 4547
rect 2949 4548 3014 4549
rect 2958 4550 3017 4551
rect 2961 4552 2966 4553
rect 2964 4554 2987 4555
rect 2979 4556 3032 4557
rect 2982 4558 3035 4559
rect 2985 4560 3050 4561
rect 2991 4562 3020 4563
rect 2994 4564 3023 4565
rect 3015 4566 3077 4567
rect 3021 4568 3068 4569
rect 3024 4570 3080 4571
rect 3027 4572 3056 4573
rect 3030 4574 3044 4575
rect 3033 4576 3083 4577
rect 3039 4578 3089 4579
rect 3042 4580 3092 4581
rect 3048 4582 3122 4583
rect 3058 4584 3242 4585
rect 3073 4586 3142 4587
rect 3081 4588 3215 4589
rect 3087 4590 3125 4591
rect 3090 4592 3095 4593
rect 3099 4592 3128 4593
rect 3106 4594 3246 4595
rect 3112 4596 3151 4597
rect 3111 4598 3283 4599
rect 3114 4600 3245 4601
rect 3118 4602 3121 4603
rect 3117 4604 3255 4605
rect 3123 4606 3264 4607
rect 3133 4608 3257 4609
rect 3139 4610 3272 4611
rect 3147 4612 3182 4613
rect 3157 4614 3242 4615
rect 3177 4616 3236 4617
rect 3051 4618 3236 4619
rect 3184 4620 3188 4621
rect 3193 4620 3364 4621
rect 3144 4622 3193 4623
rect 3195 4622 3203 4623
rect 3198 4624 3206 4625
rect 3204 4626 3239 4627
rect 3207 4628 3270 4629
rect 3093 4630 3269 4631
rect 3210 4632 3227 4633
rect 3213 4634 3230 4635
rect 3216 4636 3233 4637
rect 3219 4638 3322 4639
rect 3222 4640 3330 4641
rect 3238 4642 3313 4643
rect 3251 4644 3316 4645
rect 3260 4646 3263 4647
rect 3259 4648 3341 4649
rect 3266 4650 3315 4651
rect 3265 4652 3292 4653
rect 3274 4654 3304 4655
rect 3277 4656 3348 4657
rect 3279 4658 3284 4659
rect 3280 4660 3310 4661
rect 3286 4662 3307 4663
rect 3294 4664 3338 4665
rect 2575 4673 2785 4674
rect 2581 4675 2708 4676
rect 2582 4677 2779 4678
rect 2588 4679 2875 4680
rect 2599 4681 2751 4682
rect 2605 4683 2926 4684
rect 2609 4685 2800 4686
rect 2613 4687 2687 4688
rect 2635 4689 2874 4690
rect 2628 4691 2636 4692
rect 2642 4691 2869 4692
rect 2645 4693 2784 4694
rect 2649 4695 2821 4696
rect 2652 4697 2950 4698
rect 2655 4699 2663 4700
rect 2667 4699 2896 4700
rect 2680 4701 2962 4702
rect 2679 4703 2684 4704
rect 2686 4703 2699 4704
rect 2692 4705 2986 4706
rect 2692 4707 2711 4708
rect 2707 4709 2788 4710
rect 2710 4711 2758 4712
rect 2713 4713 2983 4714
rect 2723 4715 2941 4716
rect 2725 4717 2980 4718
rect 2616 4719 2727 4720
rect 2617 4721 2893 4722
rect 2735 4723 3126 4724
rect 2739 4725 2899 4726
rect 2747 4727 2818 4728
rect 2766 4729 2769 4730
rect 2774 4729 2791 4730
rect 2780 4731 2827 4732
rect 2792 4733 2833 4734
rect 2798 4735 2839 4736
rect 2805 4737 2820 4738
rect 2804 4739 2851 4740
rect 2816 4741 2845 4742
rect 2649 4743 2844 4744
rect 2823 4745 3311 4746
rect 2828 4747 2905 4748
rect 2661 4749 2904 4750
rect 2831 4751 2908 4752
rect 2837 4753 2965 4754
rect 2840 4755 2923 4756
rect 2849 4757 2917 4758
rect 2732 4759 2916 4760
rect 2732 4761 2797 4762
rect 2795 4763 2836 4764
rect 2834 4765 2863 4766
rect 2852 4767 2920 4768
rect 2855 4769 2911 4770
rect 2861 4771 2935 4772
rect 2867 4773 2944 4774
rect 2871 4775 2877 4776
rect 2879 4775 2956 4776
rect 2882 4777 2959 4778
rect 2886 4779 2892 4780
rect 2889 4781 2919 4782
rect 2897 4783 2952 4784
rect 2901 4785 2967 4786
rect 2909 4787 2989 4788
rect 2912 4789 3069 4790
rect 2927 4791 2995 4792
rect 2930 4793 2992 4794
rect 2933 4795 3016 4796
rect 2939 4797 3022 4798
rect 2957 4799 3034 4800
rect 2728 4801 3033 4802
rect 2963 4803 3025 4804
rect 2969 4805 3040 4806
rect 2975 4807 3121 4808
rect 2978 4809 3046 4810
rect 2990 4811 3028 4812
rect 2996 4813 3082 4814
rect 3002 4815 3166 4816
rect 3014 4817 3100 4818
rect 3030 4819 3036 4820
rect 3038 4819 3112 4820
rect 3042 4821 3081 4822
rect 3041 4823 3124 4824
rect 3047 4825 3052 4826
rect 3065 4825 3088 4826
rect 3083 4827 3132 4828
rect 3098 4829 3148 4830
rect 3101 4831 3151 4832
rect 3104 4833 3196 4834
rect 3090 4835 3195 4836
rect 3107 4837 3199 4838
rect 3110 4839 3193 4840
rect 3114 4841 3254 4842
rect 3113 4843 3145 4844
rect 3020 4845 3144 4846
rect 3117 4847 3236 4848
rect 3000 4849 3117 4850
rect 3122 4849 3208 4850
rect 3129 4851 3157 4852
rect 3128 4853 3217 4854
rect 3137 4855 3223 4856
rect 3141 4857 3190 4858
rect 3134 4859 3141 4860
rect 3153 4859 3211 4860
rect 3165 4861 3202 4862
rect 3093 4863 3201 4864
rect 3177 4865 3294 4866
rect 3182 4867 3214 4868
rect 3185 4869 3260 4870
rect 3188 4871 3263 4872
rect 3197 4873 3275 4874
rect 3206 4875 3281 4876
rect 3209 4877 3284 4878
rect 3219 4879 3297 4880
rect 3238 4881 3257 4882
rect 3265 4881 3335 4882
rect 3277 4883 3329 4884
rect 3289 4885 3301 4886
rect 3343 4885 3351 4886
rect 2570 4894 2704 4895
rect 2582 4896 2832 4897
rect 2589 4898 2805 4899
rect 2593 4900 2847 4901
rect 2596 4902 2665 4903
rect 2597 4904 2621 4905
rect 2600 4906 2841 4907
rect 2603 4908 2668 4909
rect 2611 4910 2781 4911
rect 2617 4912 2784 4913
rect 2623 4914 2865 4915
rect 2635 4916 2643 4917
rect 2638 4918 2659 4919
rect 2606 4920 2639 4921
rect 2641 4920 2656 4921
rect 2647 4922 2880 4923
rect 2661 4924 2862 4925
rect 2654 4926 2862 4927
rect 2663 4928 2895 4929
rect 2666 4930 2790 4931
rect 2675 4932 2693 4933
rect 2681 4934 2799 4935
rect 2707 4936 2736 4937
rect 2719 4938 2733 4939
rect 2575 4940 2733 4941
rect 2576 4942 2584 4943
rect 2738 4942 2748 4943
rect 2604 4944 2748 4945
rect 2741 4946 2751 4947
rect 2744 4948 2916 4949
rect 2689 4950 2916 4951
rect 2688 4952 2913 4953
rect 2723 4954 2913 4955
rect 2753 4956 2877 4957
rect 2765 4958 2769 4959
rect 2771 4958 2775 4959
rect 2777 4958 2793 4959
rect 2795 4958 2898 4959
rect 2795 4960 2811 4961
rect 2807 4962 2817 4963
rect 2810 4964 2820 4965
rect 2679 4966 2820 4967
rect 2813 4968 2835 4969
rect 2825 4970 2844 4971
rect 2828 4972 2844 4973
rect 2831 4974 2856 4975
rect 2651 4976 2856 4977
rect 2852 4978 2859 4979
rect 2870 4978 2892 4979
rect 2607 4980 2892 4981
rect 2873 4982 2889 4983
rect 2882 4984 2886 4985
rect 2867 4986 2883 4987
rect 2613 4988 2868 4989
rect 2614 4990 2727 4991
rect 2900 4990 2904 4991
rect 2903 4992 2910 4993
rect 2921 4992 2928 4993
rect 2726 4994 2928 4995
rect 2939 4994 2946 4995
rect 2939 4996 2967 4997
rect 2969 4996 2982 4997
rect 2957 4998 2970 4999
rect 2951 5000 2958 5001
rect 2933 5002 2952 5003
rect 2975 5002 2994 5003
rect 2930 5004 2976 5005
rect 2918 5006 2931 5007
rect 2837 5008 2919 5009
rect 2987 5008 3117 5009
rect 2990 5010 3027 5011
rect 2996 5012 3009 5013
rect 2978 5014 2997 5015
rect 2933 5016 2979 5017
rect 3020 5016 3072 5017
rect 3020 5018 3195 5019
rect 2710 5020 3196 5021
rect 3023 5022 3033 5023
rect 3035 5022 3141 5023
rect 3035 5024 3126 5025
rect 3038 5026 3178 5027
rect 3041 5028 3184 5029
rect 3047 5030 3057 5031
rect 3047 5032 3066 5033
rect 3068 5032 3108 5033
rect 3071 5034 3204 5035
rect 3080 5036 3090 5037
rect 2963 5038 3081 5039
rect 2695 5040 2964 5041
rect 3083 5040 3093 5041
rect 3095 5040 3099 5041
rect 3098 5042 3102 5043
rect 3104 5042 3215 5043
rect 3107 5044 3111 5045
rect 3110 5046 3114 5047
rect 3122 5046 3135 5047
rect 3128 5048 3213 5049
rect 3131 5050 3234 5051
rect 3119 5052 3233 5053
rect 3143 5054 3240 5055
rect 3153 5056 3162 5057
rect 3137 5058 3153 5059
rect 3077 5060 3138 5061
rect 3156 5060 3165 5061
rect 2936 5062 3156 5063
rect 3180 5062 3186 5063
rect 3188 5062 3257 5063
rect 3192 5064 3198 5065
rect 3209 5064 3254 5065
rect 3206 5066 3209 5067
rect 3014 5068 3206 5069
rect 3002 5070 3015 5071
rect 2563 5079 2775 5080
rect 2586 5081 2591 5082
rect 2593 5081 2742 5082
rect 2593 5083 2952 5084
rect 2596 5085 2868 5086
rect 2604 5087 2853 5088
rect 2603 5089 2844 5090
rect 2607 5091 2639 5092
rect 2617 5093 2621 5094
rect 2623 5093 2916 5094
rect 2629 5095 2642 5096
rect 2638 5097 2892 5098
rect 2642 5099 2883 5100
rect 2645 5101 2648 5102
rect 2651 5101 2898 5102
rect 2661 5103 2676 5104
rect 2664 5105 2895 5106
rect 2666 5107 2838 5108
rect 2671 5109 2772 5110
rect 2678 5111 2820 5112
rect 2632 5113 2820 5114
rect 2632 5115 2847 5116
rect 2678 5117 2715 5118
rect 2681 5119 2871 5120
rect 2681 5121 2901 5122
rect 2697 5123 2704 5124
rect 2707 5123 2727 5124
rect 2717 5125 2892 5126
rect 2720 5127 2733 5128
rect 2723 5129 2736 5130
rect 2729 5131 2931 5132
rect 2732 5133 2739 5134
rect 2735 5135 2754 5136
rect 2674 5137 2754 5138
rect 2747 5139 2877 5140
rect 2747 5141 2766 5142
rect 2765 5143 2796 5144
rect 2771 5145 2778 5146
rect 2777 5147 2790 5148
rect 2783 5149 2808 5150
rect 2786 5151 2811 5152
rect 2801 5153 2826 5154
rect 2807 5155 2832 5156
rect 2810 5157 2886 5158
rect 2816 5159 2919 5160
rect 2825 5161 3078 5162
rect 2831 5163 2850 5164
rect 2849 5165 2865 5166
rect 2864 5167 3081 5168
rect 2870 5169 2904 5170
rect 2873 5171 2889 5172
rect 2897 5171 2934 5172
rect 2900 5173 2937 5174
rect 2903 5175 2985 5176
rect 2909 5177 2928 5178
rect 2912 5179 2916 5180
rect 2703 5181 2913 5182
rect 2918 5181 2940 5182
rect 2921 5183 2979 5184
rect 2924 5185 2958 5186
rect 2930 5187 2946 5188
rect 2933 5189 3117 5190
rect 2936 5191 2988 5192
rect 2942 5193 2970 5194
rect 2948 5195 2982 5196
rect 2960 5197 3024 5198
rect 2963 5199 3138 5200
rect 2963 5201 2997 5202
rect 2966 5203 3178 5204
rect 2987 5205 3057 5206
rect 2999 5207 3093 5208
rect 3002 5209 3015 5210
rect 3008 5211 3015 5212
rect 3011 5213 3165 5214
rect 3017 5215 3069 5216
rect 3020 5217 3206 5218
rect 3026 5219 3159 5220
rect 3032 5221 3108 5222
rect 3035 5223 3068 5224
rect 3035 5225 3072 5226
rect 3038 5227 3096 5228
rect 3047 5229 3175 5230
rect 2993 5231 3049 5232
rect 3064 5231 3120 5232
rect 3070 5233 3087 5234
rect 3073 5235 3084 5236
rect 3089 5235 3147 5236
rect 3095 5237 3162 5238
rect 3098 5239 3203 5240
rect 3105 5241 3263 5242
rect 3108 5243 3181 5244
rect 3110 5245 3171 5246
rect 3089 5247 3171 5248
rect 3111 5249 3184 5250
rect 3120 5251 3193 5252
rect 3123 5253 3153 5254
rect 3131 5255 3236 5256
rect 3134 5257 3233 5258
rect 3140 5259 3247 5260
rect 3143 5261 3254 5262
rect 3164 5263 3209 5264
rect 2576 5272 2721 5273
rect 2573 5274 2577 5275
rect 2605 5274 2630 5275
rect 2610 5276 2850 5277
rect 2617 5278 2621 5279
rect 2623 5278 2665 5279
rect 2626 5280 2832 5281
rect 2632 5282 2636 5283
rect 2632 5284 2877 5285
rect 2638 5286 2811 5287
rect 2625 5288 2812 5289
rect 2649 5290 2754 5291
rect 2655 5292 3121 5293
rect 2661 5294 2689 5295
rect 2569 5296 2690 5297
rect 2570 5298 2775 5299
rect 2671 5300 2748 5301
rect 2641 5302 2749 5303
rect 2671 5304 2693 5305
rect 2674 5306 2817 5307
rect 2677 5308 2724 5309
rect 2681 5310 2871 5311
rect 2683 5312 2766 5313
rect 2686 5314 2698 5315
rect 2695 5316 2733 5317
rect 2704 5318 2736 5319
rect 2717 5320 2901 5321
rect 2680 5322 2718 5323
rect 2720 5322 2836 5323
rect 2724 5324 2872 5325
rect 2736 5326 2784 5327
rect 2739 5328 2787 5329
rect 2751 5330 2772 5331
rect 2760 5332 2778 5333
rect 2766 5334 2869 5335
rect 2769 5336 2919 5337
rect 2784 5338 2808 5339
rect 2787 5340 2802 5341
rect 2790 5342 2820 5343
rect 2796 5344 2838 5345
rect 2802 5346 2856 5347
rect 2808 5348 2853 5349
rect 2813 5350 2818 5351
rect 2814 5352 2859 5353
rect 2820 5354 2862 5355
rect 2823 5356 2874 5357
rect 2700 5358 2875 5359
rect 2825 5360 2985 5361
rect 2629 5362 2827 5363
rect 2841 5362 2892 5363
rect 2847 5364 2916 5365
rect 2850 5366 2904 5367
rect 2856 5368 2898 5369
rect 2862 5370 2910 5371
rect 2864 5372 2982 5373
rect 2710 5374 2866 5375
rect 2877 5374 3010 5375
rect 2880 5376 2931 5377
rect 2883 5378 2934 5379
rect 2886 5380 2925 5381
rect 2892 5382 2943 5383
rect 2898 5384 2937 5385
rect 2910 5386 2961 5387
rect 2922 5388 3000 5389
rect 2912 5390 3000 5391
rect 2913 5392 2964 5393
rect 2925 5394 3003 5395
rect 2934 5396 2988 5397
rect 2940 5398 3036 5399
rect 2946 5400 3038 5401
rect 2948 5402 3003 5403
rect 2955 5404 3068 5405
rect 2958 5406 3012 5407
rect 2961 5408 3015 5409
rect 2964 5410 3018 5411
rect 2966 5412 3049 5413
rect 2979 5414 3033 5415
rect 2982 5416 3046 5417
rect 3026 5418 3155 5419
rect 3040 5420 3148 5421
rect 3043 5422 3090 5423
rect 3052 5424 3109 5425
rect 3055 5426 3077 5427
rect 3055 5428 3112 5429
rect 3061 5430 3144 5431
rect 3064 5432 3141 5433
rect 3070 5434 3103 5435
rect 3073 5436 3080 5437
rect 3085 5436 3124 5437
rect 3088 5438 3171 5439
rect 3105 5440 3168 5441
rect 2563 5449 2577 5450
rect 2563 5451 2567 5452
rect 2566 5453 2606 5454
rect 2570 5455 2687 5456
rect 2573 5457 2690 5458
rect 2575 5459 2583 5460
rect 2596 5459 2636 5460
rect 2611 5461 2639 5462
rect 2615 5463 2824 5464
rect 2618 5465 2703 5466
rect 2622 5467 2803 5468
rect 2625 5469 2797 5470
rect 2632 5471 2651 5472
rect 2644 5473 2678 5474
rect 2648 5475 2821 5476
rect 2653 5477 2696 5478
rect 2662 5479 2772 5480
rect 2667 5481 2693 5482
rect 2674 5483 2711 5484
rect 2679 5485 2737 5486
rect 2683 5487 2740 5488
rect 2686 5489 2796 5490
rect 2693 5491 2884 5492
rect 2704 5493 2721 5494
rect 2705 5495 2749 5496
rect 2612 5497 2748 5498
rect 2708 5499 2752 5500
rect 2711 5501 2866 5502
rect 2714 5503 2761 5504
rect 2738 5505 2809 5506
rect 2741 5507 2785 5508
rect 2744 5509 2788 5510
rect 2750 5511 2812 5512
rect 2753 5513 2815 5514
rect 2756 5515 2791 5516
rect 2759 5517 2827 5518
rect 2762 5519 2863 5520
rect 2766 5521 2848 5522
rect 2765 5523 2881 5524
rect 2769 5525 2857 5526
rect 2768 5527 2818 5528
rect 2780 5529 2836 5530
rect 2786 5531 2842 5532
rect 2792 5533 2851 5534
rect 2801 5535 2911 5536
rect 2804 5537 2869 5538
rect 2807 5539 2872 5540
rect 2822 5541 2968 5542
rect 2825 5543 2887 5544
rect 2828 5545 2993 5546
rect 2834 5547 2926 5548
rect 2837 5549 2923 5550
rect 2840 5551 2893 5552
rect 2843 5553 2914 5554
rect 2846 5555 2920 5556
rect 2852 5557 2892 5558
rect 2864 5559 2935 5560
rect 2882 5561 2983 5562
rect 2885 5563 2941 5564
rect 2888 5565 2965 5566
rect 2898 5567 2996 5568
rect 2849 5569 2899 5570
rect 2901 5569 2986 5570
rect 2910 5571 2924 5572
rect 2913 5573 2934 5574
rect 2930 5575 2962 5576
rect 2937 5577 2947 5578
rect 2947 5579 3041 5580
rect 2955 5581 2961 5582
rect 2958 5583 3014 5584
rect 2957 5585 3059 5586
rect 2969 5587 3095 5588
rect 2972 5589 3053 5590
rect 2975 5591 3056 5592
rect 2979 5593 3003 5594
rect 3014 5593 3019 5594
rect 3027 5593 3086 5594
rect 3043 5595 3109 5596
rect 3088 5597 3099 5598
rect 2563 5606 2579 5607
rect 2581 5606 2654 5607
rect 2599 5608 2703 5609
rect 2602 5610 2769 5611
rect 2606 5612 2685 5613
rect 2612 5614 2760 5615
rect 2566 5616 2761 5617
rect 2615 5618 2757 5619
rect 2619 5620 2715 5621
rect 2619 5622 2645 5623
rect 2626 5624 2742 5625
rect 2629 5626 2745 5627
rect 2642 5628 2706 5629
rect 2645 5630 2709 5631
rect 2650 5632 2718 5633
rect 2662 5634 2706 5635
rect 2665 5636 2715 5637
rect 2681 5638 2739 5639
rect 2687 5640 2793 5641
rect 2690 5642 2796 5643
rect 2693 5644 2838 5645
rect 2693 5646 2748 5647
rect 2696 5648 2751 5649
rect 2711 5650 2799 5651
rect 2711 5652 2772 5653
rect 2739 5654 2781 5655
rect 2745 5656 2787 5657
rect 2751 5658 2805 5659
rect 2763 5660 2826 5661
rect 2769 5662 2841 5663
rect 2772 5664 2829 5665
rect 2775 5666 2853 5667
rect 2782 5668 2883 5669
rect 2801 5670 2823 5671
rect 2766 5672 2801 5673
rect 2803 5672 2850 5673
rect 2815 5674 2847 5675
rect 2830 5676 2889 5677
rect 2834 5678 2917 5679
rect 2812 5680 2834 5681
rect 2836 5680 2914 5681
rect 2840 5682 2938 5683
rect 2843 5684 2948 5685
rect 2864 5686 2892 5687
rect 2865 5688 2958 5689
rect 2868 5690 2961 5691
rect 2877 5692 2973 5693
rect 2880 5694 2976 5695
rect 2885 5696 2895 5697
rect 2753 5698 2894 5699
rect 2754 5700 2808 5701
rect 2806 5702 2819 5703
rect 2910 5702 2920 5703
rect 2969 5702 3022 5703
rect 3001 5704 3009 5705
rect 2575 5713 2620 5714
rect 2599 5715 2607 5716
rect 2602 5717 2685 5718
rect 2613 5719 2694 5720
rect 2635 5721 2697 5722
rect 2642 5723 2676 5724
rect 2652 5725 2715 5726
rect 2581 5727 2714 5728
rect 2656 5729 2682 5730
rect 2648 5731 2656 5732
rect 2658 5731 2686 5732
rect 2661 5733 2712 5734
rect 2664 5735 2718 5736
rect 2666 5737 2706 5738
rect 2678 5739 2695 5740
rect 2641 5741 2680 5742
rect 2682 5741 2698 5742
rect 2690 5743 2755 5744
rect 2687 5745 2692 5746
rect 2707 5745 2740 5746
rect 2719 5747 2735 5748
rect 2723 5749 2746 5750
rect 2728 5751 2773 5752
rect 2730 5753 2752 5754
rect 2731 5755 2776 5756
rect 2737 5757 2756 5758
rect 2740 5759 2801 5760
rect 2746 5761 2816 5762
rect 2761 5763 2807 5764
rect 2763 5765 2770 5766
rect 2764 5767 2848 5768
rect 2773 5769 2831 5770
rect 2779 5771 2813 5772
rect 2789 5773 2878 5774
rect 2803 5775 2834 5776
rect 2836 5775 2844 5776
rect 2862 5775 2866 5776
rect 2868 5775 2875 5776
rect 2880 5775 2884 5776
rect 2617 5784 2762 5785
rect 2644 5786 2665 5787
rect 2648 5788 2790 5789
rect 2651 5790 2662 5791
rect 2665 5792 2686 5793
rect 2674 5794 2692 5795
rect 2677 5796 2698 5797
rect 2694 5798 2704 5799
rect 2707 5798 2729 5799
rect 2710 5800 2732 5801
rect 2713 5802 2720 5803
rect 2737 5802 2774 5803
rect 2740 5804 2768 5805
rect 2746 5806 2787 5807
rect 2764 5808 2771 5809
rect 2623 5817 2738 5818
rect 2653 5819 2678 5820
rect 2656 5821 2669 5822
rect 2665 5823 2675 5824
rect 2707 5823 2717 5824
rect 2710 5825 2714 5826
<< metal2 >>
rect 2641 1271 2642 1281
rect 2737 1271 2738 1281
rect 2644 1273 2645 1281
rect 2647 1273 2648 1281
rect 2671 1273 2672 1281
rect 2684 1273 2685 1281
rect 2678 1275 2679 1281
rect 2687 1275 2688 1281
rect 2690 1275 2691 1281
rect 2693 1275 2694 1281
rect 2699 1275 2700 1281
rect 2708 1275 2709 1281
rect 2702 1277 2703 1281
rect 2705 1277 2706 1281
rect 2527 1287 2528 1332
rect 2533 1287 2534 1332
rect 2605 1287 2606 1332
rect 2839 1287 2840 1332
rect 2626 1289 2627 1332
rect 2645 1289 2646 1332
rect 2633 1291 2634 1332
rect 2662 1291 2663 1332
rect 2641 1285 2642 1294
rect 2677 1293 2678 1332
rect 2642 1295 2643 1332
rect 2655 1295 2656 1332
rect 2647 1285 2648 1298
rect 2674 1297 2675 1332
rect 2684 1285 2685 1298
rect 2714 1297 2715 1332
rect 2687 1285 2688 1300
rect 2721 1299 2722 1332
rect 2680 1301 2681 1332
rect 2686 1301 2687 1332
rect 2690 1285 2691 1302
rect 2727 1301 2728 1332
rect 2692 1303 2693 1332
rect 2730 1303 2731 1332
rect 2696 1305 2697 1332
rect 2711 1305 2712 1332
rect 2699 1285 2700 1308
rect 2751 1307 2752 1332
rect 2699 1309 2700 1332
rect 2708 1309 2709 1332
rect 2702 1285 2703 1312
rect 2748 1311 2749 1332
rect 2737 1285 2738 1314
rect 2827 1313 2828 1332
rect 2754 1315 2755 1332
rect 2815 1315 2816 1332
rect 2757 1317 2758 1332
rect 2851 1317 2852 1332
rect 2760 1319 2761 1332
rect 2775 1319 2776 1332
rect 2769 1321 2770 1332
rect 2794 1321 2795 1332
rect 2772 1323 2773 1332
rect 2791 1323 2792 1332
rect 2781 1325 2782 1332
rect 2845 1325 2846 1332
rect 2784 1327 2785 1332
rect 2824 1327 2825 1332
rect 2798 1329 2799 1332
rect 2830 1329 2831 1332
rect 2521 1338 2522 1385
rect 2539 1338 2540 1385
rect 2533 1336 2534 1341
rect 2545 1340 2546 1385
rect 2533 1342 2534 1385
rect 2542 1342 2543 1385
rect 2587 1342 2588 1385
rect 2596 1342 2597 1385
rect 2593 1344 2594 1385
rect 2648 1336 2649 1345
rect 2626 1346 2627 1385
rect 2689 1336 2690 1347
rect 2630 1336 2631 1349
rect 2642 1336 2643 1349
rect 2633 1336 2634 1351
rect 2645 1336 2646 1351
rect 2617 1352 2618 1385
rect 2646 1352 2647 1385
rect 2665 1336 2666 1353
rect 2711 1336 2712 1353
rect 2668 1354 2669 1385
rect 2674 1336 2675 1355
rect 2623 1356 2624 1385
rect 2674 1356 2675 1385
rect 2671 1358 2672 1385
rect 2677 1336 2678 1359
rect 2680 1358 2681 1385
rect 2686 1336 2687 1359
rect 2704 1358 2705 1385
rect 2708 1336 2709 1359
rect 2723 1358 2724 1385
rect 2798 1358 2799 1385
rect 2726 1360 2727 1385
rect 2727 1336 2728 1361
rect 2741 1360 2742 1385
rect 2751 1336 2752 1361
rect 2744 1362 2745 1385
rect 2754 1336 2755 1363
rect 2747 1364 2748 1385
rect 2748 1336 2749 1365
rect 2750 1364 2751 1385
rect 2757 1336 2758 1365
rect 2753 1366 2754 1385
rect 2760 1336 2761 1367
rect 2756 1368 2757 1385
rect 2772 1336 2773 1369
rect 2769 1336 2770 1371
rect 2771 1370 2772 1385
rect 2768 1372 2769 1385
rect 2794 1336 2795 1373
rect 2781 1336 2782 1375
rect 2866 1374 2867 1385
rect 2792 1376 2793 1385
rect 2805 1336 2806 1377
rect 2808 1336 2809 1377
rect 2863 1376 2864 1385
rect 2815 1378 2816 1385
rect 2836 1336 2837 1379
rect 2827 1336 2828 1381
rect 2833 1380 2834 1385
rect 2827 1382 2828 1385
rect 2839 1336 2840 1383
rect 2875 1382 2876 1385
rect 2895 1382 2896 1385
rect 2539 1389 2540 1392
rect 2620 1391 2621 1478
rect 2542 1389 2543 1394
rect 2561 1393 2562 1478
rect 2533 1395 2534 1478
rect 2543 1395 2544 1478
rect 2549 1395 2550 1478
rect 2558 1395 2559 1478
rect 2564 1395 2565 1478
rect 2861 1395 2862 1478
rect 2593 1389 2594 1398
rect 2611 1397 2612 1478
rect 2608 1399 2609 1478
rect 2661 1399 2662 1478
rect 2614 1401 2615 1478
rect 2721 1401 2722 1478
rect 2617 1403 2618 1478
rect 2682 1403 2683 1478
rect 2623 1389 2624 1406
rect 2643 1405 2644 1478
rect 2623 1407 2624 1478
rect 2715 1407 2716 1478
rect 2626 1389 2627 1410
rect 2709 1409 2710 1478
rect 2629 1389 2630 1412
rect 2706 1411 2707 1478
rect 2630 1413 2631 1478
rect 2739 1413 2740 1478
rect 2633 1415 2634 1478
rect 2697 1415 2698 1478
rect 2637 1417 2638 1478
rect 2736 1417 2737 1478
rect 2652 1419 2653 1478
rect 2664 1419 2665 1478
rect 2668 1389 2669 1420
rect 2703 1419 2704 1478
rect 2671 1389 2672 1422
rect 2685 1421 2686 1478
rect 2700 1389 2701 1422
rect 2766 1421 2767 1478
rect 2711 1389 2712 1424
rect 2782 1423 2783 1478
rect 2646 1389 2647 1426
rect 2712 1425 2713 1478
rect 2545 1389 2546 1428
rect 2646 1427 2647 1478
rect 2723 1389 2724 1428
rect 2800 1427 2801 1478
rect 2726 1389 2727 1430
rect 2803 1429 2804 1478
rect 2741 1389 2742 1432
rect 2857 1431 2858 1478
rect 2747 1389 2748 1434
rect 2868 1433 2869 1478
rect 2750 1389 2751 1436
rect 2806 1435 2807 1478
rect 2753 1389 2754 1438
rect 2809 1437 2810 1478
rect 2754 1439 2755 1478
rect 2760 1439 2761 1478
rect 2756 1389 2757 1442
rect 2839 1441 2840 1478
rect 2757 1443 2758 1478
rect 2836 1443 2837 1478
rect 2763 1445 2764 1478
rect 2768 1389 2769 1446
rect 2769 1447 2770 1478
rect 2909 1389 2910 1448
rect 2771 1389 2772 1450
rect 2818 1449 2819 1478
rect 2680 1389 2681 1452
rect 2772 1451 2773 1478
rect 2679 1453 2680 1478
rect 2877 1453 2878 1478
rect 2778 1455 2779 1478
rect 2821 1455 2822 1478
rect 2792 1389 2793 1458
rect 2848 1457 2849 1478
rect 2824 1389 2825 1460
rect 2916 1459 2917 1478
rect 2744 1389 2745 1462
rect 2824 1461 2825 1478
rect 2827 1389 2828 1462
rect 2904 1461 2905 1478
rect 2830 1389 2831 1464
rect 2886 1463 2887 1478
rect 2833 1389 2834 1466
rect 2889 1465 2890 1478
rect 2798 1389 2799 1468
rect 2833 1467 2834 1478
rect 2851 1467 2852 1478
rect 2907 1467 2908 1478
rect 2863 1389 2864 1470
rect 2939 1469 2940 1478
rect 2866 1389 2867 1472
rect 2945 1471 2946 1478
rect 2875 1389 2876 1474
rect 2956 1473 2957 1478
rect 2815 1389 2816 1476
rect 2874 1475 2875 1478
rect 2910 1475 2911 1478
rect 2913 1475 2914 1478
rect 2551 1484 2552 1575
rect 2558 1482 2559 1485
rect 2560 1484 2561 1575
rect 2561 1482 2562 1485
rect 2563 1484 2564 1575
rect 2564 1482 2565 1485
rect 2611 1482 2612 1485
rect 2636 1484 2637 1575
rect 2617 1482 2618 1487
rect 2780 1486 2781 1575
rect 2620 1482 2621 1489
rect 2659 1488 2660 1575
rect 2623 1482 2624 1491
rect 2712 1482 2713 1491
rect 2626 1492 2627 1575
rect 2677 1492 2678 1575
rect 2630 1494 2631 1575
rect 2715 1482 2716 1495
rect 2649 1482 2650 1497
rect 2706 1482 2707 1497
rect 2661 1482 2662 1499
rect 2783 1498 2784 1575
rect 2643 1482 2644 1501
rect 2662 1500 2663 1575
rect 2674 1500 2675 1575
rect 2762 1500 2763 1575
rect 2679 1482 2680 1503
rect 2968 1502 2969 1575
rect 2685 1482 2686 1505
rect 2711 1504 2712 1575
rect 2689 1506 2690 1575
rect 2965 1506 2966 1575
rect 2693 1508 2694 1575
rect 2754 1482 2755 1509
rect 2697 1482 2698 1511
rect 2729 1510 2730 1575
rect 2696 1512 2697 1575
rect 2798 1512 2799 1575
rect 2703 1482 2704 1515
rect 2717 1514 2718 1575
rect 2709 1482 2710 1517
rect 2747 1516 2748 1575
rect 2739 1482 2740 1519
rect 2789 1518 2790 1575
rect 2800 1482 2801 1519
rect 2846 1518 2847 1575
rect 2671 1520 2672 1575
rect 2801 1520 2802 1575
rect 2803 1482 2804 1521
rect 2840 1520 2841 1575
rect 2806 1482 2807 1523
rect 2831 1522 2832 1575
rect 2818 1482 2819 1525
rect 2864 1524 2865 1575
rect 2809 1482 2810 1527
rect 2819 1526 2820 1575
rect 2766 1482 2767 1529
rect 2810 1528 2811 1575
rect 2682 1482 2683 1531
rect 2765 1530 2766 1575
rect 2824 1482 2825 1531
rect 2858 1530 2859 1575
rect 2772 1482 2773 1533
rect 2825 1532 2826 1575
rect 2836 1482 2837 1533
rect 2837 1532 2838 1575
rect 2848 1482 2849 1533
rect 2900 1532 2901 1575
rect 2785 1482 2786 1535
rect 2849 1534 2850 1575
rect 2736 1482 2737 1537
rect 2786 1536 2787 1575
rect 2735 1538 2736 1575
rect 2778 1482 2779 1539
rect 2868 1482 2869 1539
rect 2892 1482 2893 1539
rect 2646 1482 2647 1541
rect 2891 1540 2892 1575
rect 2646 1542 2647 1575
rect 2652 1482 2653 1543
rect 2874 1482 2875 1543
rect 2987 1542 2988 1575
rect 2833 1482 2834 1545
rect 2873 1544 2874 1575
rect 2775 1482 2776 1547
rect 2834 1546 2835 1575
rect 2757 1482 2758 1549
rect 2774 1548 2775 1575
rect 2686 1550 2687 1575
rect 2756 1550 2757 1575
rect 2877 1482 2878 1551
rect 2897 1550 2898 1575
rect 2721 1482 2722 1553
rect 2876 1552 2877 1575
rect 2664 1482 2665 1555
rect 2720 1554 2721 1575
rect 2886 1482 2887 1555
rect 2953 1554 2954 1575
rect 2821 1482 2822 1557
rect 2885 1556 2886 1575
rect 2769 1482 2770 1559
rect 2822 1558 2823 1575
rect 2904 1482 2905 1559
rect 2944 1558 2945 1575
rect 2851 1482 2852 1561
rect 2903 1560 2904 1575
rect 2913 1482 2914 1561
rect 2959 1560 2960 1575
rect 2916 1482 2917 1563
rect 2962 1562 2963 1575
rect 2939 1482 2940 1565
rect 3004 1564 3005 1575
rect 2956 1482 2957 1567
rect 3007 1566 3008 1575
rect 2889 1482 2890 1569
rect 2956 1568 2957 1575
rect 2760 1482 2761 1571
rect 2888 1570 2889 1575
rect 2971 1570 2972 1575
rect 2980 1570 2981 1575
rect 2974 1572 2975 1575
rect 2977 1572 2978 1575
rect 2551 1581 2552 1680
rect 2551 1579 2552 1582
rect 2560 1579 2561 1582
rect 2651 1581 2652 1680
rect 2563 1579 2564 1584
rect 2654 1583 2655 1680
rect 2605 1585 2606 1680
rect 3104 1585 3105 1680
rect 2656 1579 2657 1588
rect 2762 1579 2763 1588
rect 2659 1579 2660 1590
rect 2713 1589 2714 1680
rect 2662 1579 2663 1592
rect 2685 1591 2686 1680
rect 2667 1593 2668 1680
rect 2765 1579 2766 1594
rect 2693 1579 2694 1596
rect 2791 1595 2792 1680
rect 2711 1579 2712 1598
rect 2758 1597 2759 1680
rect 2717 1579 2718 1600
rect 2764 1599 2765 1680
rect 2677 1579 2678 1602
rect 2716 1601 2717 1680
rect 2636 1579 2637 1604
rect 2676 1603 2677 1680
rect 2720 1579 2721 1604
rect 2794 1603 2795 1680
rect 2722 1605 2723 1680
rect 2864 1579 2865 1606
rect 2729 1579 2730 1608
rect 2806 1607 2807 1680
rect 2747 1579 2748 1610
rect 2803 1609 2804 1680
rect 2746 1611 2747 1680
rect 2756 1579 2757 1612
rect 2768 1579 2769 1612
rect 2861 1611 2862 1680
rect 2780 1579 2781 1614
rect 2828 1613 2829 1680
rect 2631 1615 2632 1680
rect 2779 1615 2780 1680
rect 2783 1579 2784 1616
rect 2831 1615 2832 1680
rect 2626 1579 2627 1618
rect 2782 1617 2783 1680
rect 2798 1579 2799 1618
rect 2855 1617 2856 1680
rect 2789 1579 2790 1620
rect 2797 1619 2798 1680
rect 2810 1579 2811 1620
rect 2812 1619 2813 1680
rect 2837 1579 2838 1620
rect 2867 1619 2868 1680
rect 2638 1621 2639 1680
rect 2837 1621 2838 1680
rect 2846 1579 2847 1622
rect 2891 1621 2892 1680
rect 2708 1579 2709 1624
rect 2846 1623 2847 1680
rect 2623 1579 2624 1626
rect 2707 1625 2708 1680
rect 2849 1579 2850 1626
rect 2894 1625 2895 1680
rect 2774 1579 2775 1628
rect 2849 1627 2850 1680
rect 2634 1629 2635 1680
rect 2773 1629 2774 1680
rect 2873 1579 2874 1630
rect 2913 1579 2914 1630
rect 2819 1579 2820 1632
rect 2912 1631 2913 1680
rect 2819 1633 2820 1680
rect 2840 1579 2841 1634
rect 2822 1579 2823 1636
rect 2873 1635 2874 1680
rect 2876 1579 2877 1636
rect 2948 1635 2949 1680
rect 2825 1579 2826 1638
rect 2876 1637 2877 1680
rect 2649 1579 2650 1640
rect 2825 1639 2826 1680
rect 2885 1579 2886 1640
rect 2927 1639 2928 1680
rect 2834 1579 2835 1642
rect 2885 1641 2886 1680
rect 2786 1579 2787 1644
rect 2834 1643 2835 1680
rect 2888 1579 2889 1644
rect 2930 1643 2931 1680
rect 2771 1579 2772 1646
rect 2888 1645 2889 1680
rect 2735 1579 2736 1648
rect 2770 1647 2771 1680
rect 2612 1649 2613 1680
rect 2734 1649 2735 1680
rect 2897 1579 2898 1650
rect 2951 1649 2952 1680
rect 2916 1579 2917 1652
rect 2980 1651 2981 1680
rect 2858 1579 2859 1654
rect 2915 1653 2916 1680
rect 2801 1579 2802 1656
rect 2858 1655 2859 1680
rect 2953 1579 2954 1656
rect 3020 1655 3021 1680
rect 2909 1657 2910 1680
rect 2954 1657 2955 1680
rect 2956 1579 2957 1658
rect 3023 1657 3024 1680
rect 2959 1579 2960 1660
rect 3014 1659 3015 1680
rect 2900 1579 2901 1662
rect 2960 1661 2961 1680
rect 2962 1579 2963 1662
rect 3002 1661 3003 1680
rect 2903 1579 2904 1664
rect 2963 1663 2964 1680
rect 2965 1579 2966 1664
rect 3026 1663 3027 1680
rect 2968 1579 2969 1666
rect 3029 1665 3030 1680
rect 2971 1579 2972 1668
rect 2998 1579 2999 1668
rect 2944 1579 2945 1670
rect 2999 1669 3000 1680
rect 2921 1671 2922 1680
rect 2945 1671 2946 1680
rect 2974 1579 2975 1672
rect 2984 1579 2985 1672
rect 3004 1579 3005 1672
rect 3063 1671 3064 1680
rect 3007 1579 3008 1674
rect 3066 1673 3067 1680
rect 3044 1675 3045 1680
rect 3055 1579 3056 1676
rect 3047 1677 3048 1680
rect 3052 1579 3053 1678
rect 2533 1686 2534 1819
rect 2654 1684 2655 1687
rect 2551 1684 2552 1689
rect 2593 1688 2594 1819
rect 2575 1690 2576 1819
rect 2663 1690 2664 1819
rect 2590 1692 2591 1819
rect 2625 1692 2626 1819
rect 2605 1684 2606 1695
rect 2734 1684 2735 1695
rect 2605 1696 2606 1819
rect 2904 1696 2905 1819
rect 2619 1684 2620 1699
rect 2773 1684 2774 1699
rect 2619 1700 2620 1819
rect 2803 1684 2804 1701
rect 2612 1684 2613 1703
rect 2802 1702 2803 1819
rect 2628 1704 2629 1819
rect 2667 1684 2668 1705
rect 2634 1706 2635 1819
rect 2679 1684 2680 1707
rect 2643 1708 2644 1819
rect 2764 1684 2765 1709
rect 2660 1710 2661 1819
rect 2676 1684 2677 1711
rect 2696 1710 2697 1819
rect 2713 1684 2714 1711
rect 2699 1712 2700 1819
rect 2707 1684 2708 1713
rect 2705 1714 2706 1819
rect 2716 1684 2717 1715
rect 2730 1714 2731 1819
rect 3018 1714 3019 1819
rect 2748 1716 2749 1819
rect 2758 1684 2759 1717
rect 2766 1716 2767 1819
rect 2779 1684 2780 1717
rect 2772 1718 2773 1819
rect 2837 1684 2838 1719
rect 2770 1684 2771 1721
rect 2838 1720 2839 1819
rect 2769 1722 2770 1819
rect 2782 1684 2783 1723
rect 2778 1724 2779 1819
rect 2791 1684 2792 1725
rect 2781 1726 2782 1819
rect 2794 1684 2795 1727
rect 2784 1728 2785 1819
rect 2797 1684 2798 1729
rect 2746 1684 2747 1731
rect 2796 1730 2797 1819
rect 2790 1732 2791 1819
rect 2806 1684 2807 1733
rect 2685 1684 2686 1735
rect 2805 1734 2806 1819
rect 2684 1736 2685 1819
rect 2888 1684 2889 1737
rect 2808 1738 2809 1819
rect 2828 1684 2829 1739
rect 2669 1740 2670 1819
rect 2829 1740 2830 1819
rect 2812 1684 2813 1743
rect 2919 1742 2920 1819
rect 2811 1744 2812 1819
rect 2831 1684 2832 1745
rect 2820 1746 2821 1819
rect 2825 1684 2826 1747
rect 2638 1684 2639 1749
rect 2826 1748 2827 1819
rect 2637 1750 2638 1819
rect 2651 1684 2652 1751
rect 2622 1684 2623 1753
rect 2650 1752 2651 1819
rect 2823 1752 2824 1819
rect 2834 1684 2835 1753
rect 2631 1754 2632 1819
rect 2835 1754 2836 1819
rect 2846 1684 2847 1755
rect 2847 1754 2848 1819
rect 2853 1754 2854 1819
rect 2873 1684 2874 1755
rect 2855 1684 2856 1757
rect 2865 1756 2866 1819
rect 2856 1758 2857 1819
rect 2876 1684 2877 1759
rect 2861 1684 2862 1761
rect 2901 1760 2902 1819
rect 2867 1684 2868 1763
rect 2877 1762 2878 1819
rect 2858 1684 2859 1765
rect 2868 1764 2869 1819
rect 2849 1684 2850 1767
rect 2859 1766 2860 1819
rect 2733 1768 2734 1819
rect 2850 1768 2851 1819
rect 2883 1768 2884 1819
rect 2885 1684 2886 1769
rect 2894 1684 2895 1769
rect 2925 1768 2926 1819
rect 2907 1770 2908 1819
rect 2930 1684 2931 1771
rect 2909 1684 2910 1773
rect 2967 1772 2968 1819
rect 2921 1684 2922 1775
rect 3012 1774 3013 1819
rect 2931 1776 2932 1819
rect 2948 1684 2949 1777
rect 2726 1778 2727 1819
rect 2949 1778 2950 1819
rect 2937 1780 2938 1819
rect 2945 1684 2946 1781
rect 2951 1684 2952 1781
rect 3089 1780 3090 1819
rect 2952 1782 2953 1819
rect 2969 1684 2970 1783
rect 2955 1784 2956 1819
rect 2976 1684 2977 1785
rect 2958 1786 2959 1819
rect 2960 1684 2961 1787
rect 2961 1788 2962 1819
rect 2963 1684 2964 1789
rect 2973 1788 2974 1819
rect 3113 1684 3114 1789
rect 2976 1790 2977 1819
rect 3002 1684 3003 1791
rect 2983 1684 2984 1793
rect 2990 1684 2991 1793
rect 2994 1792 2995 1819
rect 3014 1684 3015 1793
rect 2927 1684 2928 1795
rect 3015 1794 3016 1819
rect 2891 1684 2892 1797
rect 2928 1796 2929 1819
rect 2999 1684 3000 1797
rect 3000 1796 3001 1819
rect 3003 1796 3004 1819
rect 3097 1684 3098 1797
rect 3006 1798 3007 1819
rect 3151 1798 3152 1819
rect 3020 1684 3021 1801
rect 3055 1800 3056 1819
rect 3021 1802 3022 1819
rect 3026 1684 3027 1803
rect 2915 1684 2916 1805
rect 3027 1804 3028 1819
rect 3023 1684 3024 1807
rect 3058 1806 3059 1819
rect 3029 1684 3030 1809
rect 3074 1808 3075 1819
rect 3043 1810 3044 1819
rect 3044 1684 3045 1811
rect 3046 1810 3047 1819
rect 3047 1684 3048 1811
rect 3063 1684 3064 1811
rect 3112 1810 3113 1819
rect 2964 1812 2965 1819
rect 3064 1812 3065 1819
rect 3066 1684 3067 1813
rect 3072 1684 3073 1813
rect 2912 1684 2913 1815
rect 3071 1814 3072 1819
rect 3083 1814 3084 1819
rect 3119 1814 3120 1819
rect 3106 1816 3107 1819
rect 3109 1816 3110 1819
rect 2548 1823 2549 1826
rect 2578 1823 2579 1826
rect 2552 1823 2553 1828
rect 2575 1823 2576 1828
rect 2587 1823 2588 1828
rect 2663 1823 2664 1828
rect 2593 1823 2594 1830
rect 2599 1829 2600 1968
rect 2593 1831 2594 1968
rect 2714 1831 2715 1968
rect 2605 1823 2606 1834
rect 2817 1833 2818 1968
rect 2619 1835 2620 1968
rect 2705 1823 2706 1836
rect 2622 1823 2623 1838
rect 2625 1823 2626 1838
rect 2637 1823 2638 1838
rect 2652 1837 2653 1968
rect 2634 1823 2635 1840
rect 2636 1839 2637 1968
rect 2640 1823 2641 1840
rect 2823 1823 2824 1840
rect 2647 1823 2648 1842
rect 2865 1823 2866 1842
rect 2657 1823 2658 1844
rect 2778 1823 2779 1844
rect 2660 1823 2661 1846
rect 2661 1845 2662 1968
rect 2664 1845 2665 1968
rect 2676 1845 2677 1968
rect 2667 1847 2668 1968
rect 2850 1823 2851 1848
rect 2683 1849 2684 1968
rect 2796 1823 2797 1850
rect 2687 1823 2688 1852
rect 2772 1823 2773 1852
rect 2615 1823 2616 1854
rect 2772 1853 2773 1968
rect 2690 1855 2691 1968
rect 2781 1823 2782 1856
rect 2696 1823 2697 1858
rect 2717 1857 2718 1968
rect 2699 1823 2700 1860
rect 2702 1859 2703 1968
rect 2723 1823 2724 1860
rect 2823 1859 2824 1968
rect 2730 1823 2731 1862
rect 2847 1823 2848 1862
rect 2733 1823 2734 1864
rect 2892 1863 2893 1968
rect 2748 1823 2749 1866
rect 2751 1865 2752 1968
rect 2766 1823 2767 1866
rect 2778 1865 2779 1968
rect 2655 1867 2656 1968
rect 2766 1867 2767 1968
rect 2769 1823 2770 1868
rect 2781 1867 2782 1968
rect 2784 1823 2785 1868
rect 2793 1867 2794 1968
rect 2790 1823 2791 1870
rect 2799 1869 2800 1968
rect 2790 1871 2791 1968
rect 2820 1823 2821 1872
rect 2805 1823 2806 1874
rect 2832 1873 2833 1968
rect 2829 1823 2830 1876
rect 2841 1875 2842 1968
rect 2802 1823 2803 1878
rect 2829 1877 2830 1968
rect 2838 1823 2839 1878
rect 2862 1877 2863 1968
rect 2811 1823 2812 1880
rect 2838 1879 2839 1968
rect 2726 1823 2727 1882
rect 2811 1881 2812 1968
rect 2847 1881 2848 1968
rect 3140 1823 3141 1882
rect 2856 1823 2857 1884
rect 2886 1883 2887 1968
rect 2826 1823 2827 1886
rect 2856 1885 2857 1968
rect 2859 1823 2860 1886
rect 2871 1885 2872 1968
rect 2835 1823 2836 1888
rect 2859 1887 2860 1968
rect 2808 1823 2809 1890
rect 2835 1889 2836 1968
rect 2868 1823 2869 1890
rect 2874 1889 2875 1968
rect 2877 1823 2878 1890
rect 2895 1889 2896 1968
rect 2877 1891 2878 1968
rect 2904 1823 2905 1892
rect 2889 1893 2890 1968
rect 2967 1823 2968 1894
rect 2901 1823 2902 1896
rect 2910 1895 2911 1968
rect 2904 1897 2905 1968
rect 2907 1823 2908 1898
rect 2883 1823 2884 1900
rect 2907 1899 2908 1968
rect 2853 1823 2854 1902
rect 2883 1901 2884 1968
rect 2643 1823 2644 1904
rect 2853 1903 2854 1968
rect 2913 1903 2914 1968
rect 2928 1823 2929 1904
rect 2916 1905 2917 1968
rect 2925 1823 2926 1906
rect 2919 1823 2920 1908
rect 2922 1907 2923 1968
rect 2919 1909 2920 1968
rect 2949 1823 2950 1910
rect 2931 1823 2932 1912
rect 2934 1911 2935 1968
rect 2937 1823 2938 1912
rect 2985 1911 2986 1968
rect 2940 1913 2941 1968
rect 2961 1823 2962 1914
rect 2949 1915 2950 1968
rect 3015 1823 3016 1916
rect 2958 1823 2959 1918
rect 2970 1823 2971 1918
rect 2955 1823 2956 1920
rect 2958 1919 2959 1968
rect 2952 1823 2953 1922
rect 2955 1921 2956 1968
rect 2952 1923 2953 1968
rect 3018 1823 3019 1924
rect 2964 1823 2965 1926
rect 2982 1925 2983 1968
rect 2967 1927 2968 1968
rect 3100 1823 3101 1928
rect 2979 1929 2980 1968
rect 3071 1823 3072 1930
rect 2991 1931 2992 1968
rect 3012 1823 3013 1932
rect 2994 1823 2995 1934
rect 3018 1933 3019 1968
rect 2994 1935 2995 1968
rect 3003 1823 3004 1936
rect 3000 1823 3001 1938
rect 3135 1937 3136 1968
rect 2973 1823 2974 1940
rect 3000 1939 3001 1968
rect 3006 1823 3007 1940
rect 3024 1939 3025 1968
rect 2976 1823 2977 1942
rect 3006 1941 3007 1968
rect 3021 1823 3022 1942
rect 3036 1941 3037 1968
rect 3034 1823 3035 1944
rect 3064 1823 3065 1944
rect 3043 1823 3044 1946
rect 3129 1945 3130 1968
rect 3046 1823 3047 1948
rect 3048 1947 3049 1968
rect 3045 1949 3046 1968
rect 3083 1823 3084 1950
rect 3055 1823 3056 1952
rect 3066 1951 3067 1968
rect 3058 1823 3059 1954
rect 3069 1953 3070 1968
rect 3074 1823 3075 1954
rect 3093 1823 3094 1954
rect 3092 1955 3093 1968
rect 3106 1823 3107 1956
rect 3114 1955 3115 1968
rect 3154 1823 3155 1956
rect 3117 1957 3118 1968
rect 3154 1957 3155 1968
rect 3126 1959 3127 1968
rect 3164 1959 3165 1968
rect 3132 1961 3133 1968
rect 3150 1961 3151 1968
rect 3144 1823 3145 1964
rect 3147 1963 3148 1968
rect 3144 1965 3145 1968
rect 3170 1965 3171 1968
rect 2596 1972 2597 1975
rect 2707 1974 2708 2133
rect 2599 1972 2600 1977
rect 2600 1976 2601 2133
rect 2609 1972 2610 1977
rect 2702 1972 2703 1977
rect 2587 1978 2588 2133
rect 2609 1978 2610 2133
rect 2615 1978 2616 2133
rect 2619 1972 2620 1979
rect 2619 1980 2620 2133
rect 2692 1980 2693 2133
rect 2623 1972 2624 1983
rect 2856 1972 2857 1983
rect 2626 1984 2627 2133
rect 2719 1984 2720 2133
rect 2629 1986 2630 2133
rect 2814 1986 2815 2133
rect 2633 1972 2634 1989
rect 2646 1972 2647 1989
rect 2636 1972 2637 1991
rect 2680 1990 2681 2133
rect 2649 1972 2650 1993
rect 2766 1972 2767 1993
rect 2656 1994 2657 2133
rect 2859 1972 2860 1995
rect 2658 1972 2659 1997
rect 2664 1972 2665 1997
rect 2661 1972 2662 1999
rect 2704 1998 2705 2133
rect 2683 1972 2684 2001
rect 2874 1972 2875 2001
rect 2652 1972 2653 2003
rect 2683 2002 2684 2133
rect 2642 1972 2643 2005
rect 2653 2004 2654 2133
rect 2690 1972 2691 2005
rect 2769 2004 2770 2133
rect 2695 2006 2696 2133
rect 3141 1972 3142 2007
rect 2714 1972 2715 2009
rect 2745 2008 2746 2133
rect 2717 1972 2718 2011
rect 2748 2010 2749 2133
rect 2725 2012 2726 2133
rect 2790 1972 2791 2013
rect 2732 1972 2733 2015
rect 2892 1972 2893 2015
rect 2633 2016 2634 2133
rect 2892 2016 2893 2133
rect 2772 1972 2773 2019
rect 2904 2018 2905 2133
rect 2802 2020 2803 2133
rect 2865 1972 2866 2021
rect 2823 1972 2824 2023
rect 2859 2022 2860 2133
rect 2829 1972 2830 2025
rect 2865 2024 2866 2133
rect 2647 2026 2648 2133
rect 2829 2026 2830 2133
rect 2832 1972 2833 2027
rect 2868 2026 2869 2133
rect 2742 2028 2743 2133
rect 2832 2028 2833 2133
rect 2838 1972 2839 2029
rect 2880 2028 2881 2133
rect 2886 1972 2887 2029
rect 2925 2028 2926 2133
rect 2862 1972 2863 2031
rect 2886 2030 2887 2133
rect 2901 1972 2902 2031
rect 3081 2030 3082 2133
rect 2871 1972 2872 2033
rect 2901 2032 2902 2133
rect 2847 1972 2848 2035
rect 2871 2034 2872 2133
rect 2811 1972 2812 2037
rect 2847 2036 2848 2133
rect 2778 1972 2779 2039
rect 2811 2038 2812 2133
rect 2910 1972 2911 2039
rect 2943 2038 2944 2133
rect 2913 1972 2914 2041
rect 2946 2040 2947 2133
rect 2895 1972 2896 2043
rect 2913 2042 2914 2133
rect 2735 1972 2736 2045
rect 2895 2044 2896 2133
rect 2686 1972 2687 2047
rect 2735 2046 2736 2133
rect 2605 1972 2606 2049
rect 2686 2048 2687 2133
rect 2919 1972 2920 2049
rect 2928 2048 2929 2133
rect 2889 1972 2890 2051
rect 2919 2050 2920 2133
rect 2853 1972 2854 2053
rect 2889 2052 2890 2133
rect 2817 1972 2818 2055
rect 2853 2054 2854 2133
rect 2934 1972 2935 2055
rect 2976 2054 2977 2133
rect 2940 1972 2941 2057
rect 3015 1972 3016 2057
rect 2907 1972 2908 2059
rect 2940 2058 2941 2133
rect 2877 1972 2878 2061
rect 2907 2060 2908 2133
rect 2835 1972 2836 2063
rect 2877 2062 2878 2133
rect 2793 1972 2794 2065
rect 2835 2064 2836 2133
rect 2751 1972 2752 2067
rect 2793 2066 2794 2133
rect 2751 2068 2752 2133
rect 2781 1972 2782 2069
rect 2781 2070 2782 2133
rect 2964 2070 2965 2133
rect 2967 1972 2968 2071
rect 3003 2070 3004 2133
rect 2952 1972 2953 2073
rect 2967 2072 2968 2133
rect 2979 1972 2980 2073
rect 3102 2072 3103 2133
rect 2988 1972 2989 2075
rect 3039 1972 3040 2075
rect 2955 1972 2956 2077
rect 2988 2076 2989 2133
rect 2916 1972 2917 2079
rect 2955 2078 2956 2133
rect 3000 1972 3001 2079
rect 3191 2078 3192 2133
rect 3006 1972 3007 2081
rect 3039 2080 3040 2133
rect 3012 1972 3013 2083
rect 3084 2082 3085 2133
rect 3015 2084 3016 2133
rect 3098 1972 3099 2085
rect 2982 1972 2983 2087
rect 3099 2086 3100 2133
rect 2949 1972 2950 2089
rect 2982 2088 2983 2133
rect 3018 1972 3019 2089
rect 3195 2088 3196 2133
rect 2991 1972 2992 2091
rect 3018 2090 3019 2133
rect 2958 1972 2959 2093
rect 2991 2092 2992 2133
rect 2922 1972 2923 2095
rect 2958 2094 2959 2133
rect 2883 1972 2884 2097
rect 2922 2096 2923 2133
rect 2841 1972 2842 2099
rect 2883 2098 2884 2133
rect 2799 1972 2800 2101
rect 2841 2100 2842 2133
rect 2799 2102 2800 2133
rect 2952 2102 2953 2133
rect 3027 2102 3028 2133
rect 3120 1972 3121 2103
rect 3033 2104 3034 2133
rect 3135 1972 3136 2105
rect 3036 1972 3037 2107
rect 3159 2106 3160 2133
rect 3045 1972 3046 2109
rect 3105 2108 3106 2133
rect 3024 1972 3025 2111
rect 3045 2110 3046 2133
rect 3048 1972 3049 2111
rect 3063 2110 3064 2133
rect 3075 2110 3076 2133
rect 3089 1972 3090 2111
rect 3092 1972 3093 2111
rect 3095 1972 3096 2111
rect 3066 1972 3067 2113
rect 3093 2112 3094 2133
rect 3069 1972 3070 2115
rect 3096 2114 3097 2133
rect 3114 1972 3115 2115
rect 3157 1972 3158 2115
rect 3117 1972 3118 2117
rect 3135 2116 3136 2133
rect 3122 2118 3123 2133
rect 3156 2118 3157 2133
rect 3129 1972 3130 2121
rect 3147 2120 3148 2133
rect 3132 1972 3133 2123
rect 3171 2122 3172 2133
rect 3144 1972 3145 2125
rect 3177 1972 3178 2125
rect 3126 1972 3127 2127
rect 3144 2126 3145 2133
rect 3150 1972 3151 2127
rect 3168 2126 3169 2133
rect 2994 1972 2995 2129
rect 3150 2128 3151 2133
rect 2994 2130 2995 2133
rect 3021 2130 3022 2133
rect 3174 2130 3175 2133
rect 3184 2130 3185 2133
rect 3204 2130 3205 2133
rect 3208 2130 3209 2133
rect 2594 2137 2595 2140
rect 2851 2139 2852 2294
rect 2587 2137 2588 2142
rect 2594 2141 2595 2294
rect 2603 2137 2604 2142
rect 2853 2137 2854 2142
rect 2604 2143 2605 2294
rect 2617 2143 2618 2294
rect 2619 2137 2620 2144
rect 2686 2137 2687 2144
rect 2620 2145 2621 2294
rect 2692 2137 2693 2146
rect 2622 2137 2623 2148
rect 2695 2137 2696 2148
rect 2626 2149 2627 2294
rect 2854 2149 2855 2294
rect 2633 2137 2634 2152
rect 2899 2151 2900 2294
rect 2633 2153 2634 2294
rect 2707 2137 2708 2154
rect 2637 2155 2638 2294
rect 2751 2137 2752 2156
rect 2640 2157 2641 2294
rect 2865 2137 2866 2158
rect 2643 2137 2644 2160
rect 2687 2159 2688 2294
rect 2644 2161 2645 2294
rect 2935 2161 2936 2294
rect 2650 2137 2651 2164
rect 2821 2163 2822 2294
rect 2650 2165 2651 2294
rect 2653 2137 2654 2166
rect 2653 2167 2654 2294
rect 2776 2167 2777 2294
rect 2660 2169 2661 2294
rect 2793 2137 2794 2170
rect 2666 2171 2667 2294
rect 2868 2137 2869 2172
rect 2669 2173 2670 2294
rect 2680 2137 2681 2174
rect 2672 2175 2673 2294
rect 2683 2137 2684 2176
rect 2681 2177 2682 2294
rect 2892 2137 2893 2178
rect 2693 2179 2694 2294
rect 2704 2137 2705 2180
rect 2702 2181 2703 2294
rect 2719 2137 2720 2182
rect 2733 2181 2734 2294
rect 2745 2137 2746 2182
rect 2742 2183 2743 2294
rect 2880 2137 2881 2184
rect 2748 2137 2749 2186
rect 2754 2185 2755 2294
rect 2748 2187 2749 2294
rect 2769 2137 2770 2188
rect 2794 2187 2795 2294
rect 2904 2137 2905 2188
rect 2735 2137 2736 2190
rect 2905 2189 2906 2294
rect 2809 2191 2810 2294
rect 2811 2137 2812 2192
rect 2814 2137 2815 2192
rect 2893 2191 2894 2294
rect 2827 2193 2828 2294
rect 2835 2137 2836 2194
rect 2829 2137 2830 2196
rect 2839 2195 2840 2294
rect 2845 2195 2846 2294
rect 2847 2137 2848 2196
rect 2859 2137 2860 2196
rect 2860 2195 2861 2294
rect 2866 2195 2867 2294
rect 2871 2137 2872 2196
rect 2872 2197 2873 2294
rect 2943 2137 2944 2198
rect 2881 2199 2882 2294
rect 2886 2137 2887 2200
rect 2597 2201 2598 2294
rect 2887 2201 2888 2294
rect 2895 2137 2896 2202
rect 2950 2201 2951 2294
rect 2889 2137 2890 2204
rect 2896 2203 2897 2294
rect 2606 2137 2607 2206
rect 2890 2205 2891 2294
rect 2600 2137 2601 2208
rect 2607 2207 2608 2294
rect 2601 2209 2602 2294
rect 2609 2137 2610 2210
rect 2610 2211 2611 2294
rect 2800 2211 2801 2294
rect 2901 2137 2902 2212
rect 2902 2211 2903 2294
rect 2907 2137 2908 2212
rect 2908 2211 2909 2294
rect 2913 2137 2914 2212
rect 2914 2211 2915 2294
rect 2925 2137 2926 2212
rect 2932 2211 2933 2294
rect 2919 2137 2920 2214
rect 2926 2213 2927 2294
rect 2715 2215 2716 2294
rect 2920 2215 2921 2294
rect 2928 2137 2929 2216
rect 2985 2137 2986 2216
rect 2922 2137 2923 2218
rect 2929 2217 2930 2294
rect 2955 2137 2956 2218
rect 2962 2217 2963 2294
rect 2964 2137 2965 2218
rect 2971 2217 2972 2294
rect 2958 2137 2959 2220
rect 2965 2219 2966 2294
rect 2952 2137 2953 2222
rect 2959 2221 2960 2294
rect 2946 2137 2947 2224
rect 2953 2223 2954 2294
rect 2940 2137 2941 2226
rect 2947 2225 2948 2294
rect 2967 2137 2968 2226
rect 2974 2225 2975 2294
rect 2976 2137 2977 2226
rect 3009 2137 3010 2226
rect 2991 2137 2992 2228
rect 2998 2227 2999 2294
rect 3000 2137 3001 2228
rect 3075 2137 3076 2228
rect 2994 2137 2995 2230
rect 3001 2229 3002 2294
rect 2988 2137 2989 2232
rect 2995 2231 2996 2294
rect 3015 2137 3016 2232
rect 3115 2231 3116 2294
rect 3018 2137 3019 2234
rect 3031 2233 3032 2294
rect 3027 2137 3028 2236
rect 3076 2235 3077 2294
rect 3033 2137 3034 2238
rect 3067 2237 3068 2294
rect 3037 2239 3038 2294
rect 3215 2239 3216 2294
rect 3039 2137 3040 2242
rect 3055 2241 3056 2294
rect 3045 2137 3046 2244
rect 3061 2243 3062 2294
rect 3012 2137 3013 2246
rect 3046 2245 3047 2294
rect 3003 2137 3004 2248
rect 3013 2247 3014 2294
rect 3004 2249 3005 2294
rect 3150 2137 3151 2250
rect 3063 2137 3064 2252
rect 3088 2251 3089 2294
rect 3073 2253 3074 2294
rect 3159 2137 3160 2254
rect 3079 2255 3080 2294
rect 3257 2255 3258 2294
rect 3096 2137 3097 2258
rect 3139 2257 3140 2294
rect 3105 2137 3106 2260
rect 3160 2259 3161 2294
rect 3106 2261 3107 2294
rect 3151 2261 3152 2294
rect 3112 2263 3113 2294
rect 3178 2263 3179 2294
rect 3118 2137 3119 2266
rect 3141 2137 3142 2266
rect 3081 2137 3082 2268
rect 3142 2267 3143 2294
rect 3082 2269 3083 2294
rect 3166 2269 3167 2294
rect 3125 2137 3126 2272
rect 3163 2271 3164 2294
rect 3135 2137 3136 2274
rect 3194 2273 3195 2294
rect 3093 2137 3094 2276
rect 3136 2275 3137 2294
rect 3147 2137 3148 2276
rect 3184 2275 3185 2294
rect 3099 2137 3100 2278
rect 3148 2277 3149 2294
rect 3154 2277 3155 2294
rect 3204 2277 3205 2294
rect 3156 2137 3157 2280
rect 3174 2137 3175 2280
rect 3157 2281 3158 2294
rect 3263 2281 3264 2294
rect 3168 2137 3169 2284
rect 3227 2283 3228 2294
rect 3171 2137 3172 2286
rect 3230 2285 3231 2294
rect 2612 2137 2613 2288
rect 3172 2287 3173 2294
rect 3181 2137 3182 2288
rect 3191 2137 3192 2288
rect 3144 2137 3145 2290
rect 3181 2289 3182 2294
rect 3084 2137 3085 2292
rect 3145 2291 3146 2294
rect 3201 2291 3202 2294
rect 3240 2291 3241 2294
rect 3270 2291 3271 2294
rect 3277 2291 3278 2294
rect 2587 2300 2588 2463
rect 2607 2298 2608 2301
rect 2610 2298 2611 2301
rect 2884 2298 2885 2301
rect 2611 2302 2612 2463
rect 2887 2298 2888 2303
rect 2623 2298 2624 2305
rect 2896 2298 2897 2305
rect 2625 2306 2626 2463
rect 2839 2298 2840 2307
rect 2628 2308 2629 2463
rect 2869 2308 2870 2463
rect 2633 2298 2634 2311
rect 2687 2298 2688 2311
rect 2632 2312 2633 2463
rect 2890 2298 2891 2313
rect 2640 2298 2641 2315
rect 2815 2314 2816 2463
rect 2650 2298 2651 2317
rect 2676 2316 2677 2463
rect 2656 2298 2657 2319
rect 2881 2298 2882 2319
rect 2669 2298 2670 2321
rect 2670 2320 2671 2463
rect 2672 2298 2673 2321
rect 2673 2320 2674 2463
rect 2679 2320 2680 2463
rect 2693 2298 2694 2321
rect 2681 2298 2682 2323
rect 2848 2322 2849 2463
rect 2694 2324 2695 2463
rect 2702 2298 2703 2325
rect 2718 2298 2719 2325
rect 2860 2298 2861 2325
rect 2721 2326 2722 2463
rect 2728 2326 2729 2463
rect 2731 2326 2732 2463
rect 2733 2298 2734 2327
rect 2604 2298 2605 2329
rect 2734 2328 2735 2463
rect 2754 2298 2755 2329
rect 2755 2328 2756 2463
rect 2757 2298 2758 2329
rect 2899 2298 2900 2329
rect 2661 2330 2662 2463
rect 2758 2330 2759 2463
rect 2760 2298 2761 2331
rect 2788 2298 2789 2331
rect 2764 2298 2765 2333
rect 2914 2298 2915 2333
rect 2776 2332 2777 2463
rect 2776 2298 2777 2333
rect 2782 2334 2783 2463
rect 2794 2298 2795 2335
rect 2791 2298 2792 2337
rect 3207 2336 3208 2463
rect 2797 2338 2798 2463
rect 2926 2298 2927 2339
rect 2800 2338 2801 2463
rect 2800 2298 2801 2339
rect 2809 2338 2810 2463
rect 2809 2298 2810 2339
rect 2812 2340 2813 2463
rect 2893 2298 2894 2341
rect 2833 2298 2834 2343
rect 2839 2342 2840 2463
rect 2821 2298 2822 2345
rect 2833 2344 2834 2463
rect 2620 2298 2621 2347
rect 2821 2346 2822 2463
rect 2836 2346 2837 2463
rect 2842 2298 2843 2347
rect 2851 2298 2852 2347
rect 2857 2346 2858 2463
rect 2590 2298 2591 2349
rect 2851 2348 2852 2463
rect 2590 2350 2591 2463
rect 2712 2350 2713 2463
rect 2854 2298 2855 2351
rect 2863 2350 2864 2463
rect 2593 2352 2594 2463
rect 2854 2352 2855 2463
rect 2872 2298 2873 2353
rect 2981 2352 2982 2463
rect 2600 2354 2601 2463
rect 2872 2354 2873 2463
rect 2878 2298 2879 2355
rect 2900 2354 2901 2463
rect 2666 2298 2667 2357
rect 2878 2356 2879 2463
rect 2891 2356 2892 2463
rect 2927 2356 2928 2463
rect 2902 2298 2903 2359
rect 2918 2358 2919 2463
rect 2653 2298 2654 2361
rect 2903 2360 2904 2463
rect 2630 2298 2631 2363
rect 2654 2362 2655 2463
rect 2905 2298 2906 2363
rect 2939 2362 2940 2463
rect 2866 2298 2867 2365
rect 2906 2364 2907 2463
rect 2742 2298 2743 2367
rect 2866 2366 2867 2463
rect 2743 2368 2744 2463
rect 2748 2298 2749 2369
rect 2924 2368 2925 2463
rect 3254 2298 3255 2369
rect 2929 2298 2930 2371
rect 2930 2370 2931 2463
rect 2932 2298 2933 2371
rect 2933 2370 2934 2463
rect 2947 2298 2948 2371
rect 3178 2298 3179 2371
rect 2884 2372 2885 2463
rect 2948 2372 2949 2463
rect 2959 2298 2960 2373
rect 2960 2372 2961 2463
rect 2962 2298 2963 2373
rect 2978 2372 2979 2463
rect 2971 2298 2972 2375
rect 3026 2374 3027 2463
rect 2908 2298 2909 2377
rect 2972 2376 2973 2463
rect 2984 2376 2985 2463
rect 3059 2376 3060 2463
rect 2987 2378 2988 2463
rect 3099 2378 3100 2463
rect 2998 2298 2999 2381
rect 3017 2380 3018 2463
rect 3001 2298 3002 2383
rect 3047 2382 3048 2463
rect 3004 2298 3005 2385
rect 3050 2384 3051 2463
rect 2965 2298 2966 2387
rect 3005 2386 3006 2463
rect 2953 2298 2954 2389
rect 2966 2388 2967 2463
rect 2935 2298 2936 2391
rect 2954 2390 2955 2463
rect 2845 2298 2846 2393
rect 2936 2392 2937 2463
rect 2635 2394 2636 2463
rect 2845 2394 2846 2463
rect 3007 2298 3008 2395
rect 3190 2298 3191 2395
rect 2827 2298 2828 2397
rect 3189 2396 3190 2463
rect 2682 2398 2683 2463
rect 2827 2398 2828 2463
rect 3013 2298 3014 2399
rect 3029 2398 3030 2463
rect 3019 2298 3020 2401
rect 3053 2400 3054 2463
rect 3022 2298 3023 2403
rect 3043 2298 3044 2403
rect 2974 2298 2975 2405
rect 3023 2404 3024 2463
rect 2920 2298 2921 2407
rect 2975 2406 2976 2463
rect 3037 2298 3038 2407
rect 3243 2298 3244 2407
rect 3041 2408 3042 2463
rect 3197 2298 3198 2409
rect 3055 2298 3056 2411
rect 3266 2410 3267 2463
rect 2995 2298 2996 2413
rect 3056 2412 3057 2463
rect 3067 2298 3068 2413
rect 3071 2412 3072 2463
rect 3073 2298 3074 2413
rect 3086 2412 3087 2463
rect 3076 2298 3077 2415
rect 3245 2414 3246 2463
rect 3077 2416 3078 2463
rect 3280 2416 3281 2463
rect 3079 2298 3080 2419
rect 3290 2418 3291 2463
rect 3088 2298 3089 2421
rect 3102 2420 3103 2463
rect 2950 2298 2951 2423
rect 3089 2422 3090 2463
rect 2794 2424 2795 2463
rect 2951 2424 2952 2463
rect 3106 2298 3107 2425
rect 3126 2424 3127 2463
rect 3108 2426 3109 2463
rect 3184 2298 3185 2427
rect 3112 2298 3113 2429
rect 3132 2428 3133 2463
rect 3120 2430 3121 2463
rect 3129 2430 3130 2463
rect 3142 2298 3143 2431
rect 3151 2298 3152 2431
rect 3031 2298 3032 2433
rect 3141 2432 3142 2463
rect 3136 2298 3137 2435
rect 3150 2434 3151 2463
rect 3115 2298 3116 2437
rect 3135 2436 3136 2463
rect 3145 2298 3146 2437
rect 3148 2298 3149 2437
rect 3154 2298 3155 2437
rect 3187 2298 3188 2437
rect 3139 2298 3140 2439
rect 3153 2438 3154 2463
rect 3138 2440 3139 2463
rect 3157 2298 3158 2441
rect 2875 2298 2876 2443
rect 3156 2442 3157 2463
rect 2621 2444 2622 2463
rect 2875 2444 2876 2463
rect 3163 2298 3164 2445
rect 3166 2298 3167 2445
rect 3082 2298 3083 2447
rect 3165 2446 3166 2463
rect 3160 2298 3161 2449
rect 3162 2448 3163 2463
rect 3061 2298 3062 2451
rect 3159 2450 3160 2463
rect 3172 2298 3173 2451
rect 3186 2450 3187 2463
rect 3183 2452 3184 2463
rect 3269 2452 3270 2463
rect 3201 2298 3202 2455
rect 3211 2298 3212 2455
rect 3181 2298 3182 2457
rect 3210 2456 3211 2463
rect 3218 2298 3219 2457
rect 3247 2298 3248 2457
rect 3227 2298 3228 2459
rect 3239 2458 3240 2463
rect 3174 2460 3175 2463
rect 3227 2460 3228 2463
rect 3230 2298 3231 2461
rect 3242 2460 3243 2463
rect 2593 2467 2594 2470
rect 2915 2469 2916 2664
rect 2600 2467 2601 2472
rect 2851 2467 2852 2472
rect 2600 2473 2601 2664
rect 2731 2467 2732 2474
rect 2604 2467 2605 2476
rect 2848 2467 2849 2476
rect 2603 2477 2604 2664
rect 2771 2477 2772 2664
rect 2607 2467 2608 2480
rect 2912 2479 2913 2664
rect 2587 2467 2588 2482
rect 2606 2481 2607 2664
rect 2618 2467 2619 2482
rect 2849 2481 2850 2664
rect 2625 2467 2626 2484
rect 2857 2467 2858 2484
rect 2630 2485 2631 2664
rect 2640 2485 2641 2664
rect 2635 2467 2636 2488
rect 2852 2487 2853 2664
rect 2642 2467 2643 2490
rect 2897 2489 2898 2664
rect 2658 2467 2659 2492
rect 2743 2467 2744 2492
rect 2661 2467 2662 2494
rect 2836 2467 2837 2494
rect 2670 2467 2671 2496
rect 2696 2495 2697 2664
rect 2673 2467 2674 2498
rect 2705 2497 2706 2664
rect 2676 2467 2677 2500
rect 2819 2499 2820 2664
rect 2679 2467 2680 2502
rect 2687 2501 2688 2664
rect 2682 2467 2683 2504
rect 2815 2467 2816 2504
rect 2626 2505 2627 2664
rect 2816 2505 2817 2664
rect 2681 2507 2682 2664
rect 2878 2467 2879 2508
rect 2694 2467 2695 2510
rect 2738 2509 2739 2664
rect 2702 2511 2703 2664
rect 2918 2467 2919 2512
rect 2712 2467 2713 2514
rect 2732 2513 2733 2664
rect 2714 2515 2715 2664
rect 2812 2467 2813 2516
rect 2726 2517 2727 2664
rect 2854 2467 2855 2518
rect 2728 2467 2729 2520
rect 3253 2519 3254 2664
rect 2734 2467 2735 2522
rect 2774 2521 2775 2664
rect 2750 2523 2751 2664
rect 2948 2467 2949 2524
rect 2776 2467 2777 2526
rect 2804 2525 2805 2664
rect 2619 2527 2620 2664
rect 2777 2527 2778 2664
rect 2800 2467 2801 2528
rect 2909 2527 2910 2664
rect 2755 2467 2756 2530
rect 2801 2529 2802 2664
rect 2581 2467 2582 2532
rect 2756 2531 2757 2664
rect 2827 2467 2828 2532
rect 2858 2531 2859 2664
rect 2839 2467 2840 2534
rect 2882 2533 2883 2664
rect 2845 2467 2846 2536
rect 2894 2535 2895 2664
rect 2809 2467 2810 2538
rect 2846 2537 2847 2664
rect 2869 2467 2870 2538
rect 2918 2537 2919 2664
rect 2833 2467 2834 2540
rect 2870 2539 2871 2664
rect 2872 2467 2873 2540
rect 2921 2539 2922 2664
rect 2758 2467 2759 2542
rect 2873 2541 2874 2664
rect 2759 2543 2760 2664
rect 2782 2467 2783 2544
rect 2888 2467 2889 2544
rect 2966 2467 2967 2544
rect 2633 2545 2634 2664
rect 2888 2545 2889 2664
rect 2900 2467 2901 2546
rect 2948 2545 2949 2664
rect 2863 2467 2864 2548
rect 2900 2547 2901 2664
rect 2821 2467 2822 2550
rect 2864 2549 2865 2664
rect 2924 2467 2925 2550
rect 2984 2549 2985 2664
rect 2875 2467 2876 2552
rect 2924 2551 2925 2664
rect 2930 2467 2931 2552
rect 2990 2551 2991 2664
rect 2685 2467 2686 2554
rect 2930 2553 2931 2664
rect 2933 2467 2934 2554
rect 2993 2553 2994 2664
rect 2936 2467 2937 2556
rect 2966 2555 2967 2664
rect 2831 2557 2832 2664
rect 2936 2557 2937 2664
rect 2939 2467 2940 2558
rect 2969 2557 2970 2664
rect 2954 2467 2955 2560
rect 2996 2559 2997 2664
rect 2623 2561 2624 2664
rect 2954 2561 2955 2664
rect 2972 2467 2973 2562
rect 3002 2561 3003 2664
rect 2975 2467 2976 2564
rect 3011 2563 3012 2664
rect 2978 2467 2979 2566
rect 3020 2565 3021 2664
rect 2951 2467 2952 2568
rect 2978 2567 2979 2664
rect 2903 2467 2904 2570
rect 2951 2569 2952 2664
rect 2866 2467 2867 2572
rect 2903 2571 2904 2664
rect 2987 2467 2988 2572
rect 3113 2571 3114 2664
rect 2927 2467 2928 2574
rect 2987 2573 2988 2664
rect 2584 2467 2585 2576
rect 2927 2575 2928 2664
rect 3005 2467 3006 2576
rect 3035 2575 3036 2664
rect 2891 2467 2892 2578
rect 3005 2577 3006 2664
rect 3017 2467 3018 2578
rect 3092 2467 3093 2578
rect 2960 2467 2961 2580
rect 3017 2579 3018 2664
rect 2906 2467 2907 2582
rect 2960 2581 2961 2664
rect 2596 2583 2597 2664
rect 2906 2583 2907 2664
rect 3023 2467 3024 2584
rect 3062 2467 3063 2584
rect 3026 2467 3027 2586
rect 3059 2467 3060 2586
rect 3029 2467 3030 2588
rect 3083 2587 3084 2664
rect 3041 2467 3042 2590
rect 3234 2589 3235 2664
rect 3044 2591 3045 2664
rect 3099 2467 3100 2592
rect 3047 2467 3048 2594
rect 3155 2593 3156 2664
rect 3050 2467 3051 2596
rect 3179 2595 3180 2664
rect 2981 2467 2982 2598
rect 3050 2597 3051 2664
rect 2753 2599 2754 2664
rect 2981 2599 2982 2664
rect 3053 2467 3054 2600
rect 3089 2599 3090 2664
rect 2654 2467 2655 2602
rect 3053 2601 3054 2664
rect 3056 2467 3057 2602
rect 3092 2601 3093 2664
rect 3056 2603 3057 2664
rect 3129 2467 3130 2604
rect 3071 2467 3072 2606
rect 3122 2605 3123 2664
rect 3077 2467 3078 2608
rect 3287 2467 3288 2608
rect 3077 2609 3078 2664
rect 3262 2609 3263 2664
rect 3086 2467 3087 2612
rect 3146 2611 3147 2664
rect 3102 2467 3103 2614
rect 3158 2613 3159 2664
rect 3038 2615 3039 2664
rect 3101 2615 3102 2664
rect 3119 2615 3120 2664
rect 3141 2467 3142 2616
rect 3126 2467 3127 2618
rect 3201 2467 3202 2618
rect 3128 2619 3129 2664
rect 3135 2467 3136 2620
rect 3132 2467 3133 2622
rect 3213 2467 3214 2622
rect 3131 2623 3132 2664
rect 3259 2623 3260 2664
rect 3134 2625 3135 2664
rect 3273 2467 3274 2626
rect 3138 2467 3139 2628
rect 3269 2627 3270 2664
rect 3143 2629 3144 2664
rect 3290 2467 3291 2630
rect 3150 2467 3151 2632
rect 3194 2631 3195 2664
rect 3149 2633 3150 2664
rect 3248 2467 3249 2634
rect 3153 2467 3154 2636
rect 3197 2635 3198 2664
rect 2876 2637 2877 2664
rect 3152 2637 3153 2664
rect 3174 2467 3175 2638
rect 3225 2637 3226 2664
rect 3204 2467 3205 2640
rect 3220 2467 3221 2640
rect 3168 2467 3169 2642
rect 3203 2641 3204 2664
rect 3183 2467 3184 2644
rect 3219 2643 3220 2664
rect 3162 2467 3163 2646
rect 3182 2645 3183 2664
rect 3207 2467 3208 2646
rect 3272 2645 3273 2664
rect 3210 2467 3211 2648
rect 3275 2647 3276 2664
rect 3041 2649 3042 2664
rect 3210 2649 3211 2664
rect 3216 2467 3217 2650
rect 3244 2649 3245 2664
rect 3223 2467 3224 2652
rect 3281 2651 3282 2664
rect 3186 2467 3187 2654
rect 3222 2653 3223 2664
rect 3165 2467 3166 2656
rect 3185 2655 3186 2664
rect 3108 2467 3109 2658
rect 3164 2657 3165 2664
rect 3228 2657 3229 2664
rect 3278 2657 3279 2664
rect 3239 2467 3240 2660
rect 3290 2659 3291 2664
rect 3242 2467 3243 2662
rect 3293 2661 3294 2664
rect 3303 2661 3304 2664
rect 3317 2661 3318 2664
rect 2584 2670 2585 2877
rect 2765 2670 2766 2877
rect 2596 2668 2597 2673
rect 2918 2668 2919 2673
rect 2606 2668 2607 2675
rect 2613 2674 2614 2877
rect 2581 2676 2582 2877
rect 2607 2676 2608 2877
rect 2609 2668 2610 2677
rect 2822 2676 2823 2877
rect 2616 2668 2617 2679
rect 2921 2668 2922 2679
rect 2619 2668 2620 2681
rect 2714 2668 2715 2681
rect 2603 2668 2604 2683
rect 2619 2682 2620 2877
rect 2623 2682 2624 2877
rect 2900 2668 2901 2683
rect 2633 2684 2634 2877
rect 2677 2684 2678 2877
rect 2637 2668 2638 2687
rect 3116 2686 3117 2877
rect 2647 2688 2648 2877
rect 2858 2668 2859 2689
rect 2654 2668 2655 2691
rect 2945 2690 2946 2877
rect 2658 2692 2659 2877
rect 2900 2692 2901 2877
rect 2672 2668 2673 2695
rect 2966 2668 2967 2695
rect 2683 2696 2684 2877
rect 2687 2668 2688 2697
rect 2681 2668 2682 2699
rect 2686 2698 2687 2877
rect 2693 2668 2694 2699
rect 2870 2668 2871 2699
rect 2692 2700 2693 2877
rect 2696 2668 2697 2701
rect 2702 2700 2703 2877
rect 2852 2668 2853 2701
rect 2705 2668 2706 2703
rect 2714 2702 2715 2877
rect 2723 2702 2724 2877
rect 2726 2668 2727 2703
rect 2729 2702 2730 2877
rect 2732 2668 2733 2703
rect 2738 2668 2739 2703
rect 2741 2702 2742 2877
rect 2747 2702 2748 2877
rect 2954 2668 2955 2703
rect 2669 2668 2670 2705
rect 2954 2704 2955 2877
rect 2668 2706 2669 2877
rect 2972 2706 2973 2877
rect 2756 2668 2757 2709
rect 2762 2708 2763 2877
rect 2768 2708 2769 2877
rect 2777 2668 2778 2709
rect 2771 2668 2772 2711
rect 2780 2710 2781 2877
rect 2774 2668 2775 2713
rect 3296 2668 3297 2713
rect 2786 2714 2787 2877
rect 3014 2714 3015 2877
rect 2789 2716 2790 2877
rect 2873 2668 2874 2717
rect 2792 2718 2793 2877
rect 2951 2668 2952 2719
rect 2798 2720 2799 2877
rect 2801 2668 2802 2721
rect 2801 2722 2802 2877
rect 2903 2668 2904 2723
rect 2600 2668 2601 2725
rect 2903 2724 2904 2877
rect 2804 2724 2805 2877
rect 2804 2668 2805 2725
rect 2816 2724 2817 2877
rect 2816 2668 2817 2725
rect 2819 2724 2820 2877
rect 2819 2668 2820 2725
rect 2831 2668 2832 2727
rect 2930 2668 2931 2727
rect 2840 2728 2841 2877
rect 2846 2668 2847 2729
rect 2849 2668 2850 2729
rect 2921 2728 2922 2877
rect 2849 2730 2850 2877
rect 3002 2668 3003 2731
rect 2661 2732 2662 2877
rect 3002 2732 3003 2877
rect 2852 2734 2853 2877
rect 2864 2668 2865 2735
rect 2870 2734 2871 2877
rect 2882 2668 2883 2735
rect 2876 2736 2877 2877
rect 2894 2668 2895 2737
rect 2654 2738 2655 2877
rect 2894 2738 2895 2877
rect 2879 2668 2880 2741
rect 3005 2668 3006 2741
rect 2882 2742 2883 2877
rect 2906 2668 2907 2743
rect 2885 2744 2886 2877
rect 2909 2668 2910 2745
rect 2888 2668 2889 2747
rect 2930 2746 2931 2877
rect 2888 2748 2889 2877
rect 2912 2668 2913 2749
rect 2637 2750 2638 2877
rect 2912 2750 2913 2877
rect 2891 2752 2892 2877
rect 2915 2668 2916 2753
rect 2897 2752 2898 2877
rect 2897 2668 2898 2753
rect 2906 2754 2907 2877
rect 2924 2668 2925 2755
rect 2909 2756 2910 2877
rect 2927 2668 2928 2757
rect 2942 2756 2943 2877
rect 2948 2668 2949 2757
rect 2951 2756 2952 2877
rect 3191 2756 3192 2877
rect 2960 2668 2961 2759
rect 3008 2758 3009 2877
rect 2960 2760 2961 2877
rect 2984 2668 2985 2761
rect 2834 2762 2835 2877
rect 2984 2762 2985 2877
rect 2966 2764 2967 2877
rect 2990 2668 2991 2765
rect 2837 2766 2838 2877
rect 2990 2766 2991 2877
rect 2981 2668 2982 2769
rect 3047 2768 3048 2877
rect 2981 2770 2982 2877
rect 3059 2668 3060 2771
rect 2993 2668 2994 2773
rect 3215 2772 3216 2877
rect 3011 2668 3012 2775
rect 3074 2774 3075 2877
rect 3020 2668 3021 2777
rect 3173 2776 3174 2877
rect 3020 2778 3021 2877
rect 3038 2668 3039 2779
rect 2996 2668 2997 2781
rect 3038 2780 3039 2877
rect 2996 2782 2997 2877
rect 3017 2668 3018 2783
rect 2969 2668 2970 2785
rect 3017 2784 3018 2877
rect 2699 2668 2700 2787
rect 2969 2786 2970 2877
rect 2698 2788 2699 2877
rect 2978 2668 2979 2789
rect 2978 2790 2979 2877
rect 2987 2668 2988 2791
rect 3035 2668 3036 2791
rect 3107 2790 3108 2877
rect 3044 2668 3045 2793
rect 3068 2792 3069 2877
rect 2750 2668 2751 2795
rect 3044 2794 3045 2877
rect 3056 2668 3057 2795
rect 3265 2794 3266 2877
rect 3041 2668 3042 2797
rect 3056 2796 3057 2877
rect 3059 2796 3060 2877
rect 3104 2668 3105 2797
rect 3083 2668 3084 2799
rect 3110 2798 3111 2877
rect 3104 2800 3105 2877
rect 3176 2668 3177 2801
rect 2936 2668 2937 2803
rect 3176 2802 3177 2877
rect 3125 2804 3126 2877
rect 3155 2668 3156 2805
rect 3119 2668 3120 2807
rect 3155 2806 3156 2877
rect 3128 2668 3129 2809
rect 3262 2668 3263 2809
rect 3134 2668 3135 2811
rect 3330 2810 3331 2877
rect 3137 2812 3138 2877
rect 3206 2812 3207 2877
rect 3143 2668 3144 2815
rect 3170 2814 3171 2877
rect 3131 2668 3132 2817
rect 3143 2816 3144 2877
rect 3149 2668 3150 2817
rect 3188 2816 3189 2877
rect 3089 2668 3090 2819
rect 3149 2818 3150 2877
rect 3158 2668 3159 2819
rect 3234 2668 3235 2819
rect 3182 2668 3183 2821
rect 3240 2820 3241 2877
rect 3194 2668 3195 2823
rect 3317 2822 3318 2877
rect 3053 2668 3054 2825
rect 3194 2824 3195 2877
rect 2759 2668 2760 2827
rect 3053 2826 3054 2877
rect 2644 2668 2645 2829
rect 2759 2828 2760 2877
rect 2644 2830 2645 2877
rect 2918 2830 2919 2877
rect 3197 2668 3198 2831
rect 3314 2830 3315 2877
rect 3164 2668 3165 2833
rect 3197 2832 3198 2877
rect 3122 2668 3123 2835
rect 3164 2834 3165 2877
rect 3203 2668 3204 2835
rect 3234 2834 3235 2877
rect 3225 2668 3226 2837
rect 3278 2836 3279 2877
rect 3228 2668 3229 2839
rect 3281 2838 3282 2877
rect 3231 2668 3232 2841
rect 3268 2840 3269 2877
rect 3238 2668 3239 2843
rect 3246 2842 3247 2877
rect 3152 2668 3153 2845
rect 3237 2844 3238 2877
rect 3092 2668 3093 2847
rect 3152 2846 3153 2877
rect 3092 2848 3093 2877
rect 3324 2848 3325 2877
rect 3244 2668 3245 2851
rect 3381 2850 3382 2877
rect 3185 2668 3186 2853
rect 3243 2852 3244 2877
rect 3146 2668 3147 2855
rect 3185 2854 3186 2877
rect 3077 2668 3078 2857
rect 3146 2856 3147 2877
rect 3253 2668 3254 2857
rect 3308 2856 3309 2877
rect 3252 2858 3253 2877
rect 3339 2858 3340 2877
rect 3272 2668 3273 2861
rect 3333 2860 3334 2877
rect 3210 2668 3211 2863
rect 3272 2862 3273 2877
rect 3275 2668 3276 2863
rect 3336 2862 3337 2877
rect 3290 2668 3291 2865
rect 3358 2864 3359 2877
rect 3219 2668 3220 2867
rect 3290 2866 3291 2877
rect 3293 2668 3294 2867
rect 3361 2866 3362 2877
rect 3222 2668 3223 2869
rect 3293 2868 3294 2877
rect 3113 2668 3114 2871
rect 3222 2870 3223 2877
rect 3050 2668 3051 2873
rect 3113 2872 3114 2877
rect 2846 2874 2847 2877
rect 3050 2874 3051 2877
rect 3299 2668 3300 2875
rect 3303 2668 3304 2875
rect 3327 2874 3328 2877
rect 3327 2668 3328 2875
rect 3388 2874 3389 2877
rect 3395 2874 3396 2877
rect 2539 2883 2540 3108
rect 2546 2883 2547 3108
rect 2588 2881 2589 2884
rect 2765 2881 2766 2884
rect 2591 2881 2592 2886
rect 2888 2881 2889 2886
rect 2590 2887 2591 3108
rect 2762 2881 2763 2888
rect 2598 2881 2599 2890
rect 2932 2889 2933 3108
rect 2602 2891 2603 3108
rect 2761 2891 2762 3108
rect 2605 2893 2606 3108
rect 2607 2881 2608 2894
rect 2608 2895 2609 3108
rect 2613 2881 2614 2896
rect 2611 2897 2612 3108
rect 2719 2897 2720 3108
rect 2623 2881 2624 2900
rect 2891 2881 2892 2900
rect 2630 2881 2631 2902
rect 2909 2881 2910 2902
rect 2633 2901 2634 3108
rect 2633 2881 2634 2902
rect 2640 2903 2641 3108
rect 2737 2903 2738 3108
rect 2644 2881 2645 2906
rect 2912 2881 2913 2906
rect 2644 2907 2645 3108
rect 2759 2881 2760 2908
rect 2651 2881 2652 2910
rect 2866 2909 2867 3108
rect 2647 2881 2648 2912
rect 2651 2911 2652 3108
rect 2647 2913 2648 3108
rect 2872 2913 2873 3108
rect 2654 2881 2655 2916
rect 2876 2881 2877 2916
rect 2658 2881 2659 2918
rect 2852 2881 2853 2918
rect 2658 2919 2659 3108
rect 2974 2919 2975 3108
rect 2661 2881 2662 2922
rect 2914 2921 2915 3108
rect 2661 2923 2662 3108
rect 2741 2881 2742 2924
rect 2665 2881 2666 2926
rect 2897 2881 2898 2926
rect 2673 2927 2674 3108
rect 2894 2881 2895 2928
rect 2677 2881 2678 2930
rect 2911 2929 2912 3108
rect 2683 2881 2684 2932
rect 2688 2931 2689 3108
rect 2682 2933 2683 3108
rect 2686 2881 2687 2934
rect 2692 2881 2693 2934
rect 2694 2933 2695 3108
rect 2575 2935 2576 3108
rect 2691 2935 2692 3108
rect 2698 2881 2699 2936
rect 2935 2935 2936 3108
rect 2700 2937 2701 3108
rect 2926 2937 2927 3108
rect 2702 2881 2703 2940
rect 2969 2881 2970 2940
rect 2710 2941 2711 3108
rect 2714 2881 2715 2942
rect 2723 2881 2724 2942
rect 2734 2941 2735 3108
rect 2729 2881 2730 2944
rect 2731 2943 2732 3108
rect 2747 2881 2748 2944
rect 2978 2881 2979 2944
rect 2750 2881 2751 2946
rect 2801 2881 2802 2946
rect 2768 2881 2769 2948
rect 2785 2947 2786 3108
rect 2767 2949 2768 3108
rect 2903 2881 2904 2950
rect 2773 2951 2774 3108
rect 2780 2881 2781 2952
rect 2792 2881 2793 2952
rect 2800 2951 2801 3108
rect 2791 2953 2792 3108
rect 2798 2881 2799 2954
rect 2804 2881 2805 2954
rect 2836 2953 2837 3108
rect 2806 2955 2807 3108
rect 2816 2881 2817 2956
rect 2812 2957 2813 3108
rect 2822 2881 2823 2958
rect 2819 2881 2820 2960
rect 2821 2959 2822 3108
rect 2752 2961 2753 3108
rect 2818 2961 2819 3108
rect 2830 2961 2831 3108
rect 2840 2881 2841 2962
rect 2834 2881 2835 2964
rect 3002 2881 3003 2964
rect 2870 2881 2871 2966
rect 2875 2965 2876 3108
rect 2878 2965 2879 3108
rect 2930 2881 2931 2966
rect 2882 2881 2883 2968
rect 2890 2967 2891 3108
rect 2885 2881 2886 2970
rect 2893 2969 2894 3108
rect 2884 2971 2885 3108
rect 2918 2881 2919 2972
rect 2887 2973 2888 3108
rect 2921 2881 2922 2974
rect 2900 2881 2901 2976
rect 2902 2975 2903 3108
rect 2906 2881 2907 2976
rect 2908 2975 2909 3108
rect 2616 2881 2617 2978
rect 2905 2977 2906 3108
rect 2920 2977 2921 3108
rect 2942 2881 2943 2978
rect 2923 2979 2924 3108
rect 2945 2881 2946 2980
rect 2941 2981 2942 3108
rect 3008 2881 3009 2982
rect 2947 2983 2948 3108
rect 3014 2881 3015 2984
rect 2951 2881 2952 2986
rect 3007 2985 3008 3108
rect 2966 2881 2967 2988
rect 2977 2987 2978 3108
rect 2960 2881 2961 2990
rect 2965 2989 2966 3108
rect 2954 2881 2955 2992
rect 2959 2991 2960 3108
rect 2971 2991 2972 3108
rect 2972 2881 2973 2992
rect 2984 2881 2985 2992
rect 3268 2881 3269 2992
rect 2848 2993 2849 3108
rect 2983 2993 2984 3108
rect 2992 2993 2993 3108
rect 3017 2881 3018 2994
rect 2996 2881 2997 2996
rect 3013 2995 3014 3108
rect 2990 2881 2991 2998
rect 2995 2997 2996 3108
rect 2749 2999 2750 3108
rect 2989 2999 2990 3108
rect 3020 2881 3021 3000
rect 3031 2999 3032 3108
rect 3019 3001 3020 3108
rect 3044 2881 3045 3002
rect 3022 3003 3023 3108
rect 3047 2881 3048 3004
rect 3025 3005 3026 3108
rect 3050 2881 3051 3006
rect 3028 3007 3029 3108
rect 3053 2881 3054 3008
rect 3038 2881 3039 3010
rect 3094 3009 3095 3108
rect 3037 3011 3038 3108
rect 3116 2881 3117 3012
rect 3043 3013 3044 3108
rect 3265 2881 3266 3014
rect 3056 2881 3057 3016
rect 3064 3015 3065 3108
rect 3055 3017 3056 3108
rect 3364 2881 3365 3018
rect 3059 2881 3060 3020
rect 3225 3019 3226 3108
rect 3061 3021 3062 3108
rect 3215 3021 3216 3108
rect 3067 3023 3068 3108
rect 3068 2881 3069 3024
rect 3074 2881 3075 3024
rect 3076 3023 3077 3108
rect 3079 3023 3080 3108
rect 3367 2881 3368 3024
rect 3085 3025 3086 3108
rect 3107 2881 3108 3026
rect 3104 2881 3105 3028
rect 3121 3027 3122 3108
rect 3092 2881 3093 3030
rect 3103 3029 3104 3108
rect 3091 3031 3092 3108
rect 3173 2881 3174 3032
rect 3125 2881 3126 3034
rect 3339 2881 3340 3034
rect 3124 3035 3125 3108
rect 3208 3035 3209 3108
rect 3133 3037 3134 3108
rect 3149 2881 3150 3038
rect 3137 2881 3138 3040
rect 3139 3039 3140 3108
rect 3136 3041 3137 3108
rect 3152 2881 3153 3042
rect 3146 2881 3147 3044
rect 3324 2881 3325 3044
rect 3143 2881 3144 3046
rect 3145 3045 3146 3108
rect 3148 3045 3149 3108
rect 3321 2881 3322 3046
rect 3155 2881 3156 3048
rect 3342 2881 3343 3048
rect 3164 2881 3165 3050
rect 3166 3049 3167 3108
rect 3163 3051 3164 3108
rect 3330 2881 3331 3052
rect 3170 2881 3171 3054
rect 3407 3053 3408 3108
rect 3172 3055 3173 3108
rect 3194 2881 3195 3056
rect 3176 2881 3177 3058
rect 3206 2881 3207 3058
rect 3113 2881 3114 3060
rect 3175 3059 3176 3108
rect 3184 3059 3185 3108
rect 3185 2881 3186 3060
rect 3187 3059 3188 3108
rect 3188 2881 3189 3060
rect 3196 3059 3197 3108
rect 3197 2881 3198 3060
rect 3202 3059 3203 3108
rect 3243 2881 3244 3060
rect 3218 3061 3219 3108
rect 3222 2881 3223 3062
rect 3157 3063 3158 3108
rect 3222 3063 3223 3108
rect 3232 3063 3233 3108
rect 3283 3063 3284 3108
rect 3234 2881 3235 3066
rect 3261 2881 3262 3066
rect 3235 3067 3236 3108
rect 3317 2881 3318 3068
rect 3237 2881 3238 3070
rect 3258 2881 3259 3070
rect 3110 2881 3111 3072
rect 3238 3071 3239 3108
rect 3246 2881 3247 3072
rect 3247 3071 3248 3108
rect 3252 2881 3253 3072
rect 3298 3071 3299 3108
rect 3259 3073 3260 3108
rect 3319 3073 3320 3108
rect 3265 3075 3266 3108
rect 3331 3075 3332 3108
rect 3286 3077 3287 3108
rect 3314 2881 3315 3078
rect 3290 2881 3291 3080
rect 3313 3079 3314 3108
rect 3278 2881 3279 3082
rect 3289 3081 3290 3108
rect 3272 2881 3273 3084
rect 3277 3083 3278 3108
rect 3293 2881 3294 3084
rect 3302 2881 3303 3084
rect 3292 3085 3293 3108
rect 3355 3085 3356 3108
rect 3295 3087 3296 3108
rect 3336 2881 3337 3088
rect 3305 2881 3306 3090
rect 3316 3089 3317 3108
rect 3308 2881 3309 3092
rect 3325 3091 3326 3108
rect 3281 2881 3282 3094
rect 3307 3093 3308 3108
rect 3240 2881 3241 3096
rect 3280 3095 3281 3108
rect 3327 2881 3328 3096
rect 3370 3095 3371 3108
rect 3333 2881 3334 3098
rect 3385 2881 3386 3098
rect 3358 2881 3359 3100
rect 3364 3099 3365 3108
rect 3361 2881 3362 3102
rect 3367 3101 3368 3108
rect 3374 2881 3375 3102
rect 3384 3101 3385 3108
rect 3381 2881 3382 3104
rect 3394 3103 3395 3108
rect 3391 3105 3392 3108
rect 3398 3105 3399 3108
rect 2578 3114 2579 3349
rect 2599 3114 2600 3349
rect 2582 3116 2583 3349
rect 2691 3112 2692 3117
rect 2587 3112 2588 3119
rect 2665 3118 2666 3349
rect 2589 3120 2590 3349
rect 2777 3120 2778 3349
rect 2596 3122 2597 3349
rect 2893 3112 2894 3123
rect 2602 3112 2603 3125
rect 2611 3112 2612 3125
rect 2605 3112 2606 3127
rect 2668 3126 2669 3349
rect 2608 3112 2609 3129
rect 2616 3128 2617 3349
rect 2610 3130 2611 3349
rect 2855 3130 2856 3349
rect 2613 3132 2614 3349
rect 2884 3112 2885 3133
rect 2623 3112 2624 3135
rect 2812 3112 2813 3135
rect 2603 3136 2604 3349
rect 2813 3136 2814 3349
rect 2626 3112 2627 3139
rect 2825 3138 2826 3349
rect 2631 3140 2632 3349
rect 2767 3112 2768 3141
rect 2640 3112 2641 3143
rect 2887 3112 2888 3143
rect 2645 3144 2646 3349
rect 2951 3144 2952 3349
rect 2662 3146 2663 3349
rect 2885 3146 2886 3349
rect 2677 3148 2678 3349
rect 2905 3112 2906 3149
rect 2686 3150 2687 3349
rect 2882 3150 2883 3349
rect 2688 3112 2689 3153
rect 2704 3152 2705 3349
rect 2700 3112 2701 3155
rect 2914 3112 2915 3155
rect 2694 3112 2695 3157
rect 2701 3156 2702 3349
rect 2682 3112 2683 3159
rect 2695 3158 2696 3349
rect 2683 3160 2684 3349
rect 3031 3112 3032 3161
rect 2707 3112 2708 3163
rect 2783 3162 2784 3349
rect 2707 3164 2708 3349
rect 2878 3112 2879 3165
rect 2710 3112 2711 3167
rect 2726 3166 2727 3349
rect 2714 3168 2715 3349
rect 3011 3168 3012 3349
rect 2719 3112 2720 3171
rect 2741 3170 2742 3349
rect 2737 3112 2738 3173
rect 2840 3172 2841 3349
rect 2734 3112 2735 3175
rect 2738 3174 2739 3349
rect 2731 3112 2732 3177
rect 2735 3176 2736 3349
rect 2752 3112 2753 3177
rect 3022 3112 3023 3177
rect 2761 3112 2762 3179
rect 2768 3178 2769 3349
rect 2765 3180 2766 3349
rect 2791 3112 2792 3181
rect 2773 3112 2774 3183
rect 2795 3182 2796 3349
rect 2527 3112 2528 3185
rect 2774 3184 2775 3349
rect 2785 3112 2786 3185
rect 2789 3184 2790 3349
rect 2786 3186 2787 3349
rect 2923 3112 2924 3187
rect 2800 3112 2801 3189
rect 2906 3188 2907 3349
rect 2804 3190 2805 3349
rect 2963 3190 2964 3349
rect 2818 3112 2819 3193
rect 2846 3192 2847 3349
rect 2647 3112 2648 3195
rect 2819 3194 2820 3349
rect 2633 3112 2634 3197
rect 2648 3196 2649 3349
rect 2821 3112 2822 3197
rect 2888 3196 2889 3349
rect 2641 3198 2642 3349
rect 2822 3198 2823 3349
rect 2828 3198 2829 3349
rect 2911 3112 2912 3199
rect 2836 3112 2837 3201
rect 2864 3200 2865 3349
rect 2830 3112 2831 3203
rect 2837 3202 2838 3349
rect 2806 3112 2807 3205
rect 2831 3204 2832 3349
rect 2843 3204 2844 3349
rect 2890 3112 2891 3205
rect 2848 3112 2849 3207
rect 2947 3112 2948 3207
rect 2852 3208 2853 3349
rect 2902 3112 2903 3209
rect 2866 3112 2867 3211
rect 2870 3210 2871 3349
rect 2872 3112 2873 3211
rect 2879 3210 2880 3349
rect 2897 3210 2898 3349
rect 3007 3112 3008 3211
rect 2903 3212 2904 3349
rect 2920 3112 2921 3213
rect 2908 3112 2909 3215
rect 3370 3112 3371 3215
rect 2909 3216 2910 3349
rect 2959 3112 2960 3217
rect 2915 3218 2916 3349
rect 2965 3112 2966 3219
rect 2921 3220 2922 3349
rect 2977 3112 2978 3221
rect 2926 3112 2927 3223
rect 2927 3222 2928 3349
rect 2930 3222 2931 3349
rect 2980 3112 2981 3223
rect 2658 3112 2659 3225
rect 2981 3224 2982 3349
rect 2652 3226 2653 3349
rect 2659 3226 2660 3349
rect 2935 3112 2936 3227
rect 3041 3226 3042 3349
rect 2939 3228 2940 3349
rect 2971 3112 2972 3229
rect 2941 3112 2942 3231
rect 2978 3230 2979 3349
rect 2954 3232 2955 3349
rect 2974 3112 2975 3233
rect 2957 3234 2958 3349
rect 3013 3112 3014 3235
rect 2975 3236 2976 3349
rect 2992 3112 2993 3237
rect 2983 3112 2984 3239
rect 2987 3238 2988 3349
rect 2993 3238 2994 3349
rect 3019 3112 3020 3239
rect 2995 3112 2996 3241
rect 2996 3240 2997 3349
rect 2999 3240 3000 3349
rect 3043 3112 3044 3241
rect 3023 3242 3024 3349
rect 3025 3112 3026 3243
rect 3028 3112 3029 3243
rect 3050 3242 3051 3349
rect 3029 3244 3030 3349
rect 3037 3112 3038 3245
rect 3035 3246 3036 3349
rect 3067 3112 3068 3247
rect 3047 3248 3048 3349
rect 3155 3248 3156 3349
rect 3055 3112 3056 3251
rect 3310 3112 3311 3251
rect 3059 3252 3060 3349
rect 3061 3112 3062 3253
rect 3064 3112 3065 3253
rect 3215 3112 3216 3253
rect 3073 3112 3074 3255
rect 3193 3112 3194 3255
rect 3077 3256 3078 3349
rect 3133 3112 3134 3257
rect 3079 3112 3080 3259
rect 3352 3112 3353 3259
rect 3080 3260 3081 3349
rect 3136 3112 3137 3261
rect 3083 3262 3084 3349
rect 3232 3262 3233 3349
rect 3094 3112 3095 3265
rect 3107 3264 3108 3349
rect 3095 3266 3096 3349
rect 3225 3112 3226 3267
rect 3098 3268 3099 3349
rect 3157 3112 3158 3269
rect 3103 3112 3104 3271
rect 3271 3270 3272 3349
rect 3091 3112 3092 3273
rect 3104 3272 3105 3349
rect 3092 3274 3093 3349
rect 3145 3112 3146 3275
rect 3121 3112 3122 3277
rect 3208 3112 3209 3277
rect 3122 3278 3123 3349
rect 3184 3112 3185 3279
rect 3128 3280 3129 3349
rect 3172 3112 3173 3281
rect 3131 3282 3132 3349
rect 3175 3112 3176 3283
rect 3134 3284 3135 3349
rect 3196 3112 3197 3285
rect 3146 3286 3147 3349
rect 3195 3286 3196 3349
rect 3148 3112 3149 3289
rect 3348 3112 3349 3289
rect 3124 3112 3125 3291
rect 3149 3290 3150 3349
rect 3125 3292 3126 3349
rect 3187 3112 3188 3293
rect 3152 3294 3153 3349
rect 3259 3112 3260 3295
rect 3163 3112 3164 3297
rect 3373 3112 3374 3297
rect 3085 3112 3086 3299
rect 3162 3298 3163 3349
rect 3086 3300 3087 3349
rect 3139 3112 3140 3301
rect 3140 3302 3141 3349
rect 3202 3112 3203 3303
rect 3168 3304 3169 3349
rect 3238 3112 3239 3305
rect 3177 3306 3178 3349
rect 3384 3112 3385 3307
rect 3186 3308 3187 3349
rect 3247 3112 3248 3309
rect 3190 3112 3191 3311
rect 3256 3310 3257 3349
rect 3216 3312 3217 3349
rect 3277 3112 3278 3313
rect 3219 3314 3220 3349
rect 3280 3112 3281 3315
rect 3229 3112 3230 3317
rect 3307 3112 3308 3317
rect 3238 3318 3239 3349
rect 3298 3112 3299 3319
rect 3241 3320 3242 3349
rect 3289 3112 3290 3321
rect 3253 3322 3254 3349
rect 3259 3322 3260 3349
rect 3262 3322 3263 3349
rect 3313 3112 3314 3323
rect 3265 3112 3266 3325
rect 3322 3112 3323 3325
rect 3265 3326 3266 3349
rect 3325 3112 3326 3327
rect 2875 3112 2876 3329
rect 3324 3328 3325 3349
rect 2876 3330 2877 3349
rect 2932 3112 2933 3331
rect 2933 3332 2934 3349
rect 2989 3112 2990 3333
rect 3292 3332 3293 3349
rect 3292 3112 3293 3333
rect 3304 3332 3305 3349
rect 3364 3112 3365 3333
rect 3307 3334 3308 3349
rect 3367 3112 3368 3335
rect 3310 3336 3311 3349
rect 3331 3112 3332 3337
rect 3316 3112 3317 3339
rect 3380 3112 3381 3339
rect 3166 3112 3167 3341
rect 3317 3340 3318 3349
rect 3165 3342 3166 3349
rect 3235 3112 3236 3343
rect 3235 3344 3236 3349
rect 3295 3112 3296 3345
rect 3244 3346 3245 3349
rect 3295 3346 3296 3349
rect 2588 3355 2589 3544
rect 2749 3355 2750 3544
rect 2602 3357 2603 3544
rect 2627 3357 2628 3544
rect 2609 3359 2610 3544
rect 2876 3353 2877 3360
rect 2631 3353 2632 3362
rect 2825 3353 2826 3362
rect 2634 3353 2635 3364
rect 2948 3363 2949 3544
rect 2616 3353 2617 3366
rect 2633 3365 2634 3544
rect 2638 3353 2639 3366
rect 2698 3365 2699 3544
rect 2648 3367 2649 3544
rect 2791 3367 2792 3544
rect 2652 3353 2653 3370
rect 2879 3353 2880 3370
rect 2659 3353 2660 3372
rect 2906 3353 2907 3372
rect 2658 3373 2659 3544
rect 2789 3353 2790 3374
rect 2662 3353 2663 3376
rect 2924 3375 2925 3544
rect 2665 3353 2666 3378
rect 2680 3377 2681 3544
rect 2668 3353 2669 3380
rect 2683 3379 2684 3544
rect 2674 3381 2675 3544
rect 2722 3381 2723 3544
rect 2677 3353 2678 3384
rect 2692 3383 2693 3544
rect 2686 3353 2687 3386
rect 2909 3353 2910 3386
rect 2701 3353 2702 3388
rect 2716 3387 2717 3544
rect 2710 3353 2711 3390
rect 2918 3389 2919 3544
rect 2695 3353 2696 3392
rect 2710 3391 2711 3544
rect 2719 3391 2720 3544
rect 2731 3391 2732 3544
rect 2735 3353 2736 3392
rect 2746 3391 2747 3544
rect 2734 3393 2735 3544
rect 3026 3393 3027 3544
rect 2765 3353 2766 3396
rect 2809 3395 2810 3544
rect 2770 3397 2771 3544
rect 2828 3353 2829 3398
rect 2777 3353 2778 3400
rect 2797 3399 2798 3544
rect 2779 3401 2780 3544
rect 2875 3401 2876 3544
rect 2783 3353 2784 3404
rect 2927 3353 2928 3404
rect 2782 3405 2783 3544
rect 2857 3405 2858 3544
rect 2786 3353 2787 3408
rect 3017 3407 3018 3544
rect 2768 3353 2769 3410
rect 2785 3409 2786 3544
rect 2741 3353 2742 3412
rect 2767 3411 2768 3544
rect 2738 3353 2739 3414
rect 2740 3413 2741 3544
rect 2737 3415 2738 3544
rect 2759 3353 2760 3416
rect 2726 3353 2727 3418
rect 2758 3417 2759 3544
rect 2795 3353 2796 3418
rect 2827 3417 2828 3544
rect 2704 3353 2705 3420
rect 2794 3419 2795 3544
rect 2803 3419 2804 3544
rect 2993 3353 2994 3420
rect 2815 3421 2816 3544
rect 2975 3353 2976 3422
rect 2831 3353 2832 3424
rect 2833 3423 2834 3544
rect 2840 3353 2841 3424
rect 2872 3423 2873 3544
rect 2839 3425 2840 3544
rect 2846 3353 2847 3426
rect 2813 3353 2814 3428
rect 2845 3427 2846 3544
rect 2852 3353 2853 3428
rect 2912 3427 2913 3544
rect 2819 3353 2820 3430
rect 2851 3429 2852 3544
rect 2774 3353 2775 3432
rect 2818 3431 2819 3544
rect 2885 3353 2886 3432
rect 2936 3431 2937 3544
rect 2897 3353 2898 3434
rect 3020 3433 3021 3544
rect 2900 3353 2901 3436
rect 2987 3353 2988 3436
rect 2843 3353 2844 3438
rect 2900 3437 2901 3544
rect 2903 3353 2904 3438
rect 2960 3437 2961 3544
rect 2595 3439 2596 3544
rect 2903 3439 2904 3544
rect 2915 3353 2916 3440
rect 2990 3439 2991 3544
rect 2855 3353 2856 3442
rect 2915 3441 2916 3544
rect 2822 3353 2823 3444
rect 2854 3443 2855 3544
rect 2933 3353 2934 3444
rect 3014 3443 3015 3544
rect 2882 3353 2883 3446
rect 2933 3445 2934 3544
rect 2942 3445 2943 3544
rect 2951 3353 2952 3446
rect 2954 3353 2955 3446
rect 2993 3445 2994 3544
rect 2613 3353 2614 3448
rect 2954 3447 2955 3544
rect 2957 3353 2958 3448
rect 3032 3447 3033 3544
rect 2585 3353 2586 3450
rect 2957 3449 2958 3544
rect 2963 3353 2964 3450
rect 3059 3353 3060 3450
rect 2864 3353 2865 3452
rect 2963 3451 2964 3544
rect 2966 3451 2967 3544
rect 3062 3353 3063 3452
rect 2978 3353 2979 3454
rect 2984 3453 2985 3544
rect 2939 3353 2940 3456
rect 2978 3455 2979 3544
rect 2888 3353 2889 3458
rect 2939 3457 2940 3544
rect 2999 3353 3000 3458
rect 3195 3353 3196 3458
rect 2930 3353 2931 3460
rect 2999 3459 3000 3544
rect 2870 3353 2871 3462
rect 2930 3461 2931 3544
rect 2837 3353 2838 3464
rect 2869 3463 2870 3544
rect 3008 3463 3009 3544
rect 3023 3353 3024 3464
rect 2996 3353 2997 3466
rect 3023 3465 3024 3544
rect 2921 3353 2922 3468
rect 2996 3467 2997 3544
rect 3011 3353 3012 3468
rect 3062 3467 3063 3544
rect 3029 3353 3030 3470
rect 3155 3353 3156 3470
rect 3041 3353 3042 3472
rect 3071 3471 3072 3544
rect 3047 3353 3048 3474
rect 3068 3473 3069 3544
rect 3050 3353 3051 3476
rect 3232 3353 3233 3476
rect 2981 3353 2982 3478
rect 3050 3477 3051 3544
rect 3083 3353 3084 3478
rect 3116 3477 3117 3544
rect 3086 3353 3087 3480
rect 3179 3479 3180 3544
rect 3086 3481 3087 3544
rect 3162 3353 3163 3482
rect 3095 3353 3096 3484
rect 3155 3483 3156 3544
rect 3098 3353 3099 3486
rect 3119 3485 3120 3544
rect 3125 3353 3126 3486
rect 3331 3485 3332 3544
rect 3092 3353 3093 3488
rect 3125 3487 3126 3544
rect 3134 3353 3135 3488
rect 3269 3487 3270 3544
rect 3140 3353 3141 3490
rect 3170 3489 3171 3544
rect 3146 3353 3147 3492
rect 3182 3491 3183 3544
rect 3104 3353 3105 3494
rect 3146 3493 3147 3544
rect 3077 3353 3078 3496
rect 3104 3495 3105 3544
rect 3152 3495 3153 3544
rect 3327 3495 3328 3544
rect 3165 3353 3166 3498
rect 3206 3497 3207 3544
rect 3128 3353 3129 3500
rect 3164 3499 3165 3544
rect 3128 3501 3129 3544
rect 3345 3501 3346 3544
rect 3168 3353 3169 3504
rect 3209 3503 3210 3544
rect 3131 3353 3132 3506
rect 3167 3505 3168 3544
rect 3177 3353 3178 3506
rect 3224 3505 3225 3544
rect 3122 3353 3123 3508
rect 3176 3507 3177 3544
rect 3188 3507 3189 3544
rect 3192 3353 3193 3508
rect 3044 3509 3045 3544
rect 3191 3509 3192 3544
rect 3216 3353 3217 3510
rect 3272 3509 3273 3544
rect 3238 3353 3239 3512
rect 3334 3353 3335 3512
rect 3241 3353 3242 3514
rect 3278 3513 3279 3544
rect 3244 3353 3245 3516
rect 3281 3515 3282 3544
rect 3253 3353 3254 3518
rect 3291 3517 3292 3544
rect 3259 3353 3260 3520
rect 3312 3519 3313 3544
rect 3256 3353 3257 3522
rect 3260 3521 3261 3544
rect 3257 3523 3258 3544
rect 3274 3353 3275 3524
rect 3219 3353 3220 3526
rect 3275 3525 3276 3544
rect 3186 3353 3187 3528
rect 3218 3527 3219 3544
rect 3149 3353 3150 3530
rect 3185 3529 3186 3544
rect 3107 3353 3108 3532
rect 3149 3531 3150 3544
rect 3080 3353 3081 3534
rect 3107 3533 3108 3544
rect 3035 3353 3036 3536
rect 3080 3535 3081 3544
rect 3263 3535 3264 3544
rect 3370 3535 3371 3544
rect 3265 3353 3266 3538
rect 3318 3537 3319 3544
rect 3235 3353 3236 3540
rect 3266 3539 3267 3544
rect 3304 3353 3305 3540
rect 3357 3539 3358 3544
rect 3239 3541 3240 3544
rect 3305 3541 3306 3544
rect 3307 3353 3308 3542
rect 3360 3541 3361 3544
rect 3373 3541 3374 3544
rect 3377 3541 3378 3544
rect 2530 3550 2531 3797
rect 2761 3550 2762 3797
rect 2541 3552 2542 3797
rect 2677 3552 2678 3797
rect 2561 3554 2562 3797
rect 2642 3554 2643 3797
rect 2564 3556 2565 3797
rect 2575 3556 2576 3797
rect 2581 3548 2582 3557
rect 2680 3548 2681 3557
rect 2584 3548 2585 3559
rect 2686 3558 2687 3797
rect 2588 3548 2589 3561
rect 2683 3548 2684 3561
rect 2595 3548 2596 3563
rect 3170 3548 3171 3563
rect 2594 3564 2595 3797
rect 2900 3548 2901 3565
rect 2605 3548 2606 3567
rect 2915 3548 2916 3567
rect 2604 3568 2605 3797
rect 2836 3568 2837 3797
rect 2609 3548 2610 3571
rect 2698 3548 2699 3571
rect 2608 3572 2609 3797
rect 2863 3572 2864 3797
rect 2612 3548 2613 3575
rect 2954 3548 2955 3575
rect 2615 3576 2616 3797
rect 2636 3548 2637 3577
rect 2639 3548 2640 3577
rect 2767 3548 2768 3577
rect 2633 3548 2634 3579
rect 2639 3578 2640 3797
rect 2648 3548 2649 3579
rect 2842 3578 2843 3797
rect 2651 3548 2652 3581
rect 2851 3548 2852 3581
rect 2652 3582 2653 3797
rect 2887 3582 2888 3797
rect 2667 3548 2668 3585
rect 2933 3548 2934 3585
rect 2667 3586 2668 3797
rect 2890 3586 2891 3797
rect 2670 3548 2671 3589
rect 2725 3588 2726 3797
rect 2671 3590 2672 3797
rect 2924 3548 2925 3591
rect 2674 3548 2675 3593
rect 2740 3548 2741 3593
rect 2674 3594 2675 3797
rect 2930 3548 2931 3595
rect 2692 3548 2693 3597
rect 2698 3596 2699 3797
rect 2695 3598 2696 3797
rect 2716 3548 2717 3599
rect 2658 3548 2659 3601
rect 2716 3600 2717 3797
rect 2710 3548 2711 3603
rect 2722 3602 2723 3797
rect 2719 3604 2720 3797
rect 2731 3548 2732 3605
rect 2734 3548 2735 3605
rect 2948 3548 2949 3605
rect 2734 3606 2735 3797
rect 2770 3548 2771 3607
rect 2737 3608 2738 3797
rect 2767 3608 2768 3797
rect 2740 3610 2741 3797
rect 2746 3548 2747 3611
rect 2743 3612 2744 3797
rect 2749 3548 2750 3613
rect 2758 3548 2759 3613
rect 2764 3612 2765 3797
rect 2758 3614 2759 3797
rect 2809 3548 2810 3615
rect 2773 3616 2774 3797
rect 2818 3548 2819 3617
rect 2655 3548 2656 3619
rect 2818 3618 2819 3797
rect 2776 3620 2777 3797
rect 2791 3548 2792 3621
rect 2779 3622 2780 3797
rect 2794 3548 2795 3623
rect 2782 3548 2783 3625
rect 2999 3548 3000 3625
rect 2782 3626 2783 3797
rect 2785 3548 2786 3627
rect 2788 3626 2789 3797
rect 2797 3548 2798 3627
rect 2797 3628 2798 3797
rect 3239 3548 3240 3629
rect 2806 3548 2807 3631
rect 2978 3548 2979 3631
rect 2806 3632 2807 3797
rect 2827 3548 2828 3633
rect 2812 3548 2813 3635
rect 3014 3548 3015 3635
rect 2636 3636 2637 3797
rect 2812 3636 2813 3797
rect 2824 3636 2825 3797
rect 2845 3548 2846 3637
rect 2833 3548 2834 3639
rect 2908 3638 2909 3797
rect 2845 3640 2846 3797
rect 2854 3548 2855 3641
rect 2854 3642 2855 3797
rect 2912 3548 2913 3643
rect 2857 3548 2858 3645
rect 3004 3644 3005 3797
rect 2627 3548 2628 3647
rect 2857 3646 2858 3797
rect 2860 3646 2861 3797
rect 2957 3548 2958 3647
rect 2866 3648 2867 3797
rect 2869 3548 2870 3649
rect 2869 3650 2870 3797
rect 2872 3548 2873 3651
rect 2875 3548 2876 3651
rect 3001 3650 3002 3797
rect 2875 3652 2876 3797
rect 3017 3548 3018 3653
rect 2878 3654 2879 3797
rect 2936 3548 2937 3655
rect 2884 3656 2885 3797
rect 3284 3548 3285 3657
rect 2894 3548 2895 3659
rect 3026 3548 3027 3659
rect 2897 3548 2898 3661
rect 3212 3548 3213 3661
rect 2839 3548 2840 3663
rect 2896 3662 2897 3797
rect 2839 3664 2840 3797
rect 2903 3548 2904 3665
rect 2902 3666 2903 3797
rect 2960 3548 2961 3667
rect 2911 3668 2912 3797
rect 2939 3548 2940 3669
rect 2914 3670 2915 3797
rect 2996 3548 2997 3671
rect 2918 3548 2919 3673
rect 3188 3548 3189 3673
rect 2920 3674 2921 3797
rect 2990 3548 2991 3675
rect 2932 3676 2933 3797
rect 2966 3548 2967 3677
rect 2938 3678 2939 3797
rect 3023 3548 3024 3679
rect 2815 3548 2816 3681
rect 3022 3680 3023 3797
rect 2942 3548 2943 3683
rect 2947 3682 2948 3797
rect 2941 3684 2942 3797
rect 3032 3548 3033 3685
rect 2953 3686 2954 3797
rect 2984 3548 2985 3687
rect 2959 3688 2960 3797
rect 3044 3548 3045 3689
rect 2963 3548 2964 3691
rect 2995 3690 2996 3797
rect 2971 3692 2972 3797
rect 3050 3548 3051 3693
rect 2983 3694 2984 3797
rect 3062 3548 3063 3695
rect 2993 3548 2994 3697
rect 3025 3696 3026 3797
rect 2872 3698 2873 3797
rect 2992 3698 2993 3797
rect 2998 3698 2999 3797
rect 3171 3698 3172 3797
rect 3008 3548 3009 3701
rect 3059 3700 3060 3797
rect 3020 3548 3021 3703
rect 3034 3702 3035 3797
rect 3044 3702 3045 3797
rect 3185 3548 3186 3703
rect 3047 3704 3048 3797
rect 3209 3548 3210 3705
rect 3053 3706 3054 3797
rect 3128 3548 3129 3707
rect 3071 3548 3072 3709
rect 3110 3708 3111 3797
rect 3071 3710 3072 3797
rect 3119 3548 3120 3711
rect 3077 3712 3078 3797
rect 3155 3548 3156 3713
rect 3086 3548 3087 3715
rect 3155 3714 3156 3797
rect 3095 3548 3096 3717
rect 3149 3548 3150 3717
rect 3095 3718 3096 3797
rect 3152 3548 3153 3719
rect 3098 3720 3099 3797
rect 3283 3720 3284 3797
rect 3101 3722 3102 3797
rect 3104 3548 3105 3723
rect 3080 3548 3081 3725
rect 3104 3724 3105 3797
rect 3107 3548 3108 3725
rect 3230 3548 3231 3725
rect 3068 3548 3069 3727
rect 3107 3726 3108 3797
rect 3116 3548 3117 3727
rect 3287 3548 3288 3727
rect 3119 3728 3120 3797
rect 3176 3548 3177 3729
rect 2989 3730 2990 3797
rect 3175 3730 3176 3797
rect 3125 3548 3126 3733
rect 3324 3548 3325 3733
rect 3137 3734 3138 3797
rect 3327 3548 3328 3735
rect 3140 3736 3141 3797
rect 3146 3548 3147 3737
rect 3146 3738 3147 3797
rect 3164 3548 3165 3739
rect 3143 3740 3144 3797
rect 3164 3740 3165 3797
rect 3149 3742 3150 3797
rect 3167 3548 3168 3743
rect 3007 3744 3008 3797
rect 3168 3744 3169 3797
rect 3152 3746 3153 3797
rect 3182 3548 3183 3747
rect 3158 3748 3159 3797
rect 3224 3548 3225 3749
rect 3179 3548 3180 3751
rect 3348 3548 3349 3751
rect 3178 3752 3179 3797
rect 3291 3548 3292 3753
rect 3182 3754 3183 3797
rect 3278 3548 3279 3755
rect 3188 3756 3189 3797
rect 3275 3548 3276 3757
rect 3194 3758 3195 3797
rect 3281 3548 3282 3759
rect 3083 3760 3084 3797
rect 3280 3760 3281 3797
rect 3197 3762 3198 3797
rect 3272 3548 3273 3763
rect 3206 3548 3207 3765
rect 3377 3548 3378 3765
rect 3209 3766 3210 3797
rect 3334 3548 3335 3767
rect 3212 3768 3213 3797
rect 3266 3548 3267 3769
rect 3218 3548 3219 3771
rect 3363 3548 3364 3771
rect 3218 3772 3219 3797
rect 3252 3772 3253 3797
rect 3221 3774 3222 3797
rect 3269 3548 3270 3775
rect 3050 3776 3051 3797
rect 3269 3776 3270 3797
rect 3234 3778 3235 3797
rect 3318 3548 3319 3779
rect 3246 3780 3247 3797
rect 3297 3780 3298 3797
rect 3249 3782 3250 3797
rect 3294 3782 3295 3797
rect 3257 3548 3258 3785
rect 3308 3548 3309 3785
rect 3260 3548 3261 3787
rect 3305 3548 3306 3787
rect 3215 3788 3216 3797
rect 3259 3788 3260 3797
rect 3263 3548 3264 3789
rect 3329 3788 3330 3797
rect 3306 3790 3307 3797
rect 3357 3548 3358 3791
rect 3309 3792 3310 3797
rect 3360 3548 3361 3793
rect 3319 3794 3320 3797
rect 3366 3548 3367 3795
rect 2527 3801 2528 3804
rect 3092 3803 3093 4018
rect 2534 3801 2535 3806
rect 2761 3801 2762 3806
rect 2545 3807 2546 4018
rect 2634 3807 2635 4018
rect 2551 3801 2552 3810
rect 2677 3801 2678 3810
rect 2554 3801 2555 3812
rect 2642 3801 2643 3812
rect 2578 3801 2579 3814
rect 2587 3801 2588 3814
rect 2581 3815 2582 4018
rect 2609 3815 2610 4018
rect 2591 3817 2592 4018
rect 2690 3817 2691 4018
rect 2602 3819 2603 4018
rect 2857 3801 2858 3820
rect 2604 3801 2605 3822
rect 2854 3801 2855 3822
rect 2615 3801 2616 3824
rect 2631 3823 2632 4018
rect 2621 3825 2622 4018
rect 2678 3825 2679 4018
rect 2628 3827 2629 4018
rect 2812 3801 2813 3828
rect 2637 3829 2638 4018
rect 2824 3801 2825 3830
rect 2639 3801 2640 3832
rect 2650 3831 2651 4018
rect 2648 3801 2649 3834
rect 2818 3801 2819 3834
rect 2652 3801 2653 3836
rect 2936 3835 2937 4018
rect 2653 3837 2654 4018
rect 2655 3801 2656 3838
rect 2664 3801 2665 3838
rect 2896 3801 2897 3838
rect 2667 3801 2668 3840
rect 2908 3801 2909 3840
rect 2594 3801 2595 3842
rect 2909 3841 2910 4018
rect 2671 3801 2672 3844
rect 2975 3843 2976 4018
rect 2686 3801 2687 3846
rect 2702 3845 2703 4018
rect 2695 3801 2696 3848
rect 2711 3847 2712 4018
rect 2705 3849 2706 4018
rect 2716 3801 2717 3850
rect 2708 3851 2709 4018
rect 2719 3801 2720 3852
rect 2722 3801 2723 3852
rect 2738 3851 2739 4018
rect 2734 3801 2735 3854
rect 3011 3853 3012 4018
rect 2740 3801 2741 3856
rect 2750 3855 2751 4018
rect 2725 3801 2726 3858
rect 2741 3857 2742 4018
rect 2743 3801 2744 3858
rect 2753 3857 2754 4018
rect 2758 3801 2759 3858
rect 2813 3857 2814 4018
rect 2759 3859 2760 4018
rect 2920 3801 2921 3860
rect 2720 3861 2721 4018
rect 2921 3861 2922 4018
rect 2762 3863 2763 4018
rect 2764 3801 2765 3864
rect 2773 3801 2774 3864
rect 2828 3863 2829 4018
rect 2779 3801 2780 3866
rect 2798 3865 2799 4018
rect 2788 3801 2789 3868
rect 2801 3867 2802 4018
rect 2782 3801 2783 3870
rect 2789 3869 2790 4018
rect 2783 3871 2784 4018
rect 2998 3801 2999 3872
rect 2794 3801 2795 3874
rect 2932 3801 2933 3874
rect 2776 3801 2777 3876
rect 2795 3875 2796 4018
rect 2806 3801 2807 3876
rect 2831 3875 2832 4018
rect 2816 3877 2817 4018
rect 2987 3877 2988 4018
rect 2839 3801 2840 3880
rect 2894 3879 2895 4018
rect 2842 3801 2843 3882
rect 2855 3881 2856 4018
rect 2843 3883 2844 4018
rect 2995 3801 2996 3884
rect 2845 3801 2846 3886
rect 2858 3885 2859 4018
rect 2863 3801 2864 3886
rect 2918 3885 2919 4018
rect 2866 3801 2867 3888
rect 2897 3887 2898 4018
rect 2867 3889 2868 4018
rect 3001 3801 3002 3890
rect 2869 3801 2870 3892
rect 2900 3891 2901 4018
rect 2875 3801 2876 3894
rect 2989 3801 2990 3894
rect 2878 3801 2879 3896
rect 2927 3895 2928 4018
rect 2756 3897 2757 4018
rect 2879 3897 2880 4018
rect 2884 3801 2885 3898
rect 2933 3897 2934 4018
rect 2885 3899 2886 4018
rect 3113 3801 3114 3900
rect 2902 3801 2903 3902
rect 2951 3901 2952 4018
rect 2723 3903 2724 4018
rect 2903 3903 2904 4018
rect 2911 3801 2912 3904
rect 2930 3903 2931 4018
rect 2698 3801 2699 3906
rect 2912 3905 2913 4018
rect 2914 3801 2915 3906
rect 2969 3905 2970 4018
rect 2860 3801 2861 3908
rect 2915 3907 2916 4018
rect 2861 3909 2862 4018
rect 2887 3801 2888 3910
rect 2941 3801 2942 3910
rect 2999 3909 3000 4018
rect 2945 3911 2946 4018
rect 3034 3801 3035 3912
rect 2947 3801 2948 3914
rect 2957 3913 2958 4018
rect 2953 3801 2954 3916
rect 2981 3915 2982 4018
rect 2954 3917 2955 4018
rect 3161 3801 3162 3918
rect 2959 3801 2960 3920
rect 3125 3919 3126 4018
rect 2971 3801 2972 3922
rect 3017 3921 3018 4018
rect 2972 3923 2973 4018
rect 3004 3801 3005 3924
rect 2978 3925 2979 4018
rect 3025 3801 3026 3926
rect 3005 3927 3006 4018
rect 3044 3801 3045 3928
rect 3029 3929 3030 4018
rect 3107 3801 3108 3930
rect 3032 3931 3033 4018
rect 3110 3801 3111 3932
rect 3041 3801 3042 3934
rect 3059 3801 3060 3934
rect 3041 3935 3042 4018
rect 3143 3801 3144 3936
rect 2770 3801 2771 3938
rect 3143 3937 3144 4018
rect 2771 3939 2772 4018
rect 3309 3801 3310 3940
rect 3050 3801 3051 3942
rect 3086 3941 3087 4018
rect 3062 3943 3063 4018
rect 3241 3943 3242 4018
rect 3071 3801 3072 3946
rect 3113 3945 3114 4018
rect 3074 3947 3075 4018
rect 3140 3801 3141 3948
rect 3077 3801 3078 3950
rect 3140 3949 3141 4018
rect 3044 3951 3045 4018
rect 3077 3951 3078 4018
rect 3080 3951 3081 4018
rect 3101 3801 3102 3952
rect 3095 3801 3096 3954
rect 3280 3801 3281 3954
rect 3098 3801 3099 3956
rect 3280 3955 3281 4018
rect 3098 3957 3099 4018
rect 3146 3801 3147 3958
rect 3047 3801 3048 3960
rect 3146 3959 3147 4018
rect 3122 3961 3123 4018
rect 3155 3801 3156 3962
rect 3137 3801 3138 3964
rect 3262 3801 3263 3964
rect 3083 3801 3084 3966
rect 3137 3965 3138 4018
rect 3083 3967 3084 4018
rect 3104 3801 3105 3968
rect 3149 3801 3150 3968
rect 3164 3801 3165 3968
rect 3155 3969 3156 4018
rect 3259 3801 3260 3970
rect 3068 3971 3069 4018
rect 3259 3971 3260 4018
rect 3164 3973 3165 4018
rect 3262 3973 3263 4018
rect 3168 3801 3169 3976
rect 3256 3975 3257 4018
rect 3191 3977 3192 4018
rect 3197 3801 3198 3978
rect 3194 3801 3195 3980
rect 3224 3979 3225 4018
rect 3188 3801 3189 3982
rect 3194 3981 3195 4018
rect 3197 3981 3198 4018
rect 3315 3801 3316 3982
rect 3206 3983 3207 4018
rect 3218 3801 3219 3984
rect 3212 3801 3213 3986
rect 3218 3985 3219 4018
rect 3209 3801 3210 3988
rect 3212 3987 3213 4018
rect 3158 3801 3159 3990
rect 3209 3989 3210 4018
rect 2938 3801 2939 3992
rect 3158 3991 3159 4018
rect 2939 3993 2940 4018
rect 3022 3801 3023 3994
rect 2983 3801 2984 3996
rect 3023 3995 3024 4018
rect 2984 3997 2985 4018
rect 2992 3801 2993 3998
rect 3215 3801 3216 3998
rect 3252 3801 3253 3998
rect 3215 3999 3216 4018
rect 3266 3999 3267 4018
rect 3221 4001 3222 4018
rect 3287 3801 3288 4002
rect 3119 3801 3120 4004
rect 3287 4003 3288 4018
rect 3119 4005 3120 4018
rect 3152 3801 3153 4006
rect 3234 3801 3235 4006
rect 3302 4005 3303 4018
rect 3246 3801 3247 4008
rect 3253 4007 3254 4018
rect 3249 3801 3250 4010
rect 3319 3801 3320 4010
rect 3293 4011 3294 4018
rect 3306 3801 3307 4012
rect 3053 3801 3054 4014
rect 3306 4013 3307 4018
rect 3007 3801 3008 4016
rect 3053 4015 3054 4018
rect 3296 4015 3297 4018
rect 3322 3801 3323 4016
rect 2555 4022 2556 4025
rect 2570 4024 2571 4213
rect 2567 4026 2568 4213
rect 2634 4022 2635 4027
rect 2576 4028 2577 4213
rect 2851 4028 2852 4213
rect 2579 4030 2580 4213
rect 2586 4030 2587 4213
rect 2588 4022 2589 4031
rect 2595 4022 2596 4031
rect 2589 4032 2590 4213
rect 2690 4022 2691 4033
rect 2593 4034 2594 4213
rect 2891 4022 2892 4035
rect 2581 4022 2582 4037
rect 2890 4036 2891 4213
rect 2603 4038 2604 4213
rect 2801 4022 2802 4039
rect 2612 4040 2613 4213
rect 2672 4040 2673 4213
rect 2619 4042 2620 4213
rect 2944 4042 2945 4213
rect 2622 4044 2623 4213
rect 2831 4022 2832 4045
rect 2624 4022 2625 4047
rect 2741 4022 2742 4047
rect 2626 4048 2627 4213
rect 2734 4048 2735 4213
rect 2628 4022 2629 4051
rect 2629 4050 2630 4213
rect 2640 4022 2641 4051
rect 2912 4022 2913 4051
rect 2636 4052 2637 4213
rect 2911 4052 2912 4213
rect 2644 4022 2645 4055
rect 2984 4022 2985 4055
rect 2650 4022 2651 4057
rect 2651 4056 2652 4213
rect 2653 4022 2654 4057
rect 2708 4022 2709 4057
rect 2678 4022 2679 4059
rect 2830 4058 2831 4213
rect 2688 4060 2689 4213
rect 2791 4060 2792 4213
rect 2697 4062 2698 4213
rect 2705 4022 2706 4063
rect 2700 4064 2701 4213
rect 2711 4022 2712 4065
rect 2720 4022 2721 4065
rect 2959 4064 2960 4213
rect 2722 4066 2723 4213
rect 3007 4066 3008 4213
rect 2728 4068 2729 4213
rect 2738 4022 2739 4069
rect 2740 4068 2741 4213
rect 2750 4022 2751 4069
rect 2743 4070 2744 4213
rect 2753 4022 2754 4071
rect 2746 4072 2747 4213
rect 2762 4022 2763 4073
rect 2749 4074 2750 4213
rect 2867 4022 2868 4075
rect 2759 4022 2760 4077
rect 3293 4022 3294 4077
rect 2767 4078 2768 4213
rect 2954 4022 2955 4079
rect 2771 4022 2772 4081
rect 2981 4022 2982 4081
rect 2773 4082 2774 4213
rect 2783 4022 2784 4083
rect 2785 4082 2786 4213
rect 2795 4022 2796 4083
rect 2806 4082 2807 4213
rect 2816 4022 2817 4083
rect 2818 4082 2819 4213
rect 2828 4022 2829 4083
rect 2605 4022 2606 4085
rect 2827 4084 2828 4213
rect 2839 4084 2840 4213
rect 2855 4022 2856 4085
rect 2843 4022 2844 4087
rect 3184 4086 3185 4213
rect 2842 4088 2843 4213
rect 2858 4022 2859 4089
rect 2845 4090 2846 4213
rect 2861 4022 2862 4091
rect 2854 4092 2855 4213
rect 2939 4022 2940 4093
rect 2860 4094 2861 4213
rect 2918 4022 2919 4095
rect 2789 4022 2790 4097
rect 2917 4096 2918 4213
rect 2788 4098 2789 4213
rect 2798 4022 2799 4099
rect 2797 4100 2798 4213
rect 2813 4022 2814 4101
rect 2812 4102 2813 4213
rect 2837 4022 2838 4103
rect 2866 4102 2867 4213
rect 2879 4022 2880 4103
rect 2596 4104 2597 4213
rect 2878 4104 2879 4213
rect 2872 4106 2873 4213
rect 2885 4022 2886 4107
rect 2584 4022 2585 4109
rect 2884 4108 2885 4213
rect 2881 4110 2882 4213
rect 2894 4022 2895 4111
rect 2702 4022 2703 4113
rect 2893 4112 2894 4213
rect 2896 4112 2897 4213
rect 2897 4022 2898 4113
rect 2899 4112 2900 4213
rect 2900 4022 2901 4113
rect 2902 4112 2903 4213
rect 2903 4022 2904 4113
rect 2921 4022 2922 4113
rect 2938 4112 2939 4213
rect 2678 4114 2679 4213
rect 2920 4114 2921 4213
rect 2926 4114 2927 4213
rect 2927 4022 2928 4115
rect 2929 4114 2930 4213
rect 2930 4022 2931 4115
rect 2932 4114 2933 4213
rect 2933 4022 2934 4115
rect 2965 4114 2966 4213
rect 2992 4114 2993 4213
rect 2975 4022 2976 4117
rect 2980 4116 2981 4213
rect 2969 4022 2970 4119
rect 2974 4118 2975 4213
rect 2957 4022 2958 4121
rect 2968 4120 2969 4213
rect 2951 4022 2952 4123
rect 2956 4122 2957 4213
rect 2978 4022 2979 4123
rect 2983 4122 2984 4213
rect 2972 4022 2973 4125
rect 2977 4124 2978 4213
rect 2987 4022 2988 4125
rect 3032 4022 3033 4125
rect 2948 4022 2949 4127
rect 2986 4126 2987 4213
rect 2936 4022 2937 4129
rect 2947 4128 2948 4213
rect 2990 4022 2991 4129
rect 3029 4022 3030 4129
rect 2999 4022 3000 4131
rect 3001 4130 3002 4213
rect 3005 4022 3006 4131
rect 3040 4130 3041 4213
rect 3010 4132 3011 4213
rect 3011 4022 3012 4133
rect 3017 4022 3018 4133
rect 3019 4132 3020 4213
rect 3023 4022 3024 4133
rect 3058 4132 3059 4213
rect 3025 4134 3026 4213
rect 3181 4134 3182 4213
rect 3037 4136 3038 4213
rect 3125 4022 3126 4137
rect 3049 4138 3050 4213
rect 3098 4022 3099 4139
rect 3053 4022 3054 4141
rect 3130 4140 3131 4213
rect 3052 4142 3053 4213
rect 3157 4142 3158 4213
rect 3055 4144 3056 4213
rect 3119 4022 3120 4145
rect 3074 4022 3075 4147
rect 3332 4146 3333 4213
rect 3068 4022 3069 4149
rect 3073 4148 3074 4213
rect 3062 4022 3063 4151
rect 3067 4150 3068 4213
rect 3061 4152 3062 4213
rect 3083 4022 3084 4153
rect 3080 4022 3081 4155
rect 3103 4154 3104 4213
rect 3086 4022 3087 4157
rect 3109 4156 3110 4213
rect 3092 4022 3093 4159
rect 3227 4158 3228 4213
rect 3106 4160 3107 4213
rect 3167 4022 3168 4161
rect 3113 4022 3114 4163
rect 3203 4162 3204 4213
rect 3115 4164 3116 4213
rect 3152 4022 3153 4165
rect 3118 4166 3119 4213
rect 3188 4166 3189 4213
rect 3122 4022 3123 4169
rect 3241 4022 3242 4169
rect 3137 4022 3138 4171
rect 3302 4170 3303 4213
rect 3146 4022 3147 4173
rect 3166 4172 3167 4213
rect 3155 4022 3156 4175
rect 3260 4174 3261 4213
rect 3164 4022 3165 4177
rect 3320 4176 3321 4213
rect 3143 4022 3144 4179
rect 3163 4178 3164 4213
rect 3169 4178 3170 4213
rect 3285 4178 3286 4213
rect 3194 4022 3195 4181
rect 3200 4180 3201 4213
rect 3194 4182 3195 4213
rect 3276 4022 3277 4183
rect 3209 4022 3210 4185
rect 3236 4184 3237 4213
rect 2715 4186 2716 4213
rect 3209 4186 3210 4213
rect 3212 4022 3213 4187
rect 3248 4186 3249 4213
rect 3212 4188 3213 4213
rect 3215 4022 3216 4189
rect 3218 4022 3219 4189
rect 3251 4188 3252 4213
rect 3221 4022 3222 4191
rect 3269 4022 3270 4191
rect 3127 4192 3128 4213
rect 3221 4192 3222 4213
rect 3224 4022 3225 4193
rect 3230 4192 3231 4213
rect 3197 4022 3198 4195
rect 3224 4194 3225 4213
rect 3140 4022 3141 4197
rect 3197 4196 3198 4213
rect 3077 4022 3078 4199
rect 3139 4198 3140 4213
rect 3233 4198 3234 4213
rect 3309 4022 3310 4199
rect 3244 4022 3245 4201
rect 3253 4022 3254 4201
rect 3254 4202 3255 4213
rect 3316 4022 3317 4203
rect 3245 4204 3246 4213
rect 3316 4204 3317 4213
rect 3256 4022 3257 4207
rect 3306 4206 3307 4213
rect 3191 4022 3192 4209
rect 3257 4208 3258 4213
rect 3290 4022 3291 4209
rect 3313 4208 3314 4213
rect 3296 4022 3297 4211
rect 3299 4022 3300 4211
rect 2557 4217 2558 4220
rect 2570 4217 2571 4220
rect 2560 4217 2561 4222
rect 2564 4217 2565 4222
rect 2567 4217 2568 4222
rect 2576 4217 2577 4222
rect 2582 4217 2583 4222
rect 2730 4221 2731 4422
rect 2586 4217 2587 4224
rect 2706 4223 2707 4422
rect 2594 4225 2595 4422
rect 2881 4217 2882 4226
rect 2600 4217 2601 4228
rect 2917 4217 2918 4228
rect 2612 4217 2613 4230
rect 2682 4229 2683 4422
rect 2619 4217 2620 4232
rect 2890 4217 2891 4232
rect 2622 4217 2623 4234
rect 2851 4217 2852 4234
rect 2622 4235 2623 4422
rect 2860 4217 2861 4236
rect 2626 4217 2627 4238
rect 2715 4217 2716 4238
rect 2633 4217 2634 4240
rect 2920 4217 2921 4240
rect 2632 4241 2633 4422
rect 2947 4217 2948 4242
rect 2636 4217 2637 4244
rect 2734 4217 2735 4244
rect 2636 4245 2637 4422
rect 2740 4217 2741 4246
rect 2639 4247 2640 4422
rect 3013 4247 3014 4422
rect 2643 4249 2644 4422
rect 2971 4249 2972 4422
rect 2646 4251 2647 4422
rect 2821 4251 2822 4422
rect 2648 4217 2649 4254
rect 2845 4217 2846 4254
rect 2651 4217 2652 4256
rect 2667 4255 2668 4422
rect 2672 4217 2673 4256
rect 2688 4255 2689 4422
rect 2673 4257 2674 4422
rect 2718 4217 2719 4258
rect 2694 4259 2695 4422
rect 2851 4259 2852 4422
rect 2697 4217 2698 4262
rect 2848 4261 2849 4422
rect 2709 4263 2710 4422
rect 2743 4217 2744 4264
rect 2728 4217 2729 4266
rect 2764 4265 2765 4422
rect 2746 4217 2747 4268
rect 2800 4267 2801 4422
rect 2746 4269 2747 4422
rect 3118 4217 3119 4270
rect 2749 4217 2750 4272
rect 2995 4271 2996 4422
rect 2700 4217 2701 4274
rect 2749 4273 2750 4422
rect 2752 4217 2753 4274
rect 2992 4217 2993 4274
rect 2603 4217 2604 4276
rect 2992 4275 2993 4422
rect 2604 4277 2605 4422
rect 2608 4277 2609 4422
rect 2767 4217 2768 4278
rect 2776 4277 2777 4422
rect 2797 4217 2798 4278
rect 2857 4277 2858 4422
rect 2803 4279 2804 4422
rect 2806 4217 2807 4280
rect 2812 4217 2813 4280
rect 2860 4279 2861 4422
rect 2812 4281 2813 4422
rect 2905 4281 2906 4422
rect 2815 4283 2816 4422
rect 2854 4217 2855 4284
rect 2830 4217 2831 4286
rect 2869 4285 2870 4422
rect 2788 4217 2789 4288
rect 2830 4287 2831 4422
rect 2773 4217 2774 4290
rect 2788 4289 2789 4422
rect 2845 4289 2846 4422
rect 2965 4217 2966 4290
rect 2743 4291 2744 4422
rect 2965 4291 2966 4422
rect 2872 4217 2873 4294
rect 3016 4293 3017 4422
rect 2818 4217 2819 4296
rect 2872 4295 2873 4422
rect 2887 4295 2888 4422
rect 2902 4217 2903 4296
rect 2893 4217 2894 4298
rect 2962 4297 2963 4422
rect 2839 4217 2840 4300
rect 2893 4299 2894 4422
rect 2791 4217 2792 4302
rect 2839 4301 2840 4422
rect 2899 4217 2900 4302
rect 2917 4301 2918 4422
rect 2899 4303 2900 4422
rect 2938 4217 2939 4304
rect 2908 4217 2909 4306
rect 2947 4305 2948 4422
rect 2866 4217 2867 4308
rect 2908 4307 2909 4422
rect 2827 4217 2828 4310
rect 2866 4309 2867 4422
rect 2785 4217 2786 4312
rect 2827 4311 2828 4422
rect 2914 4217 2915 4312
rect 2989 4311 2990 4422
rect 2896 4217 2897 4314
rect 2914 4313 2915 4422
rect 2926 4217 2927 4314
rect 2953 4313 2954 4422
rect 2941 4315 2942 4422
rect 2968 4217 2969 4316
rect 2950 4217 2951 4318
rect 2998 4317 2999 4422
rect 2911 4217 2912 4320
rect 2950 4319 2951 4422
rect 2956 4217 2957 4320
rect 3300 4319 3301 4422
rect 2929 4217 2930 4322
rect 2956 4321 2957 4422
rect 2794 4323 2795 4422
rect 2929 4323 2930 4422
rect 2959 4217 2960 4324
rect 2986 4323 2987 4422
rect 2884 4217 2885 4326
rect 2959 4325 2960 4422
rect 2980 4217 2981 4326
rect 3031 4325 3032 4422
rect 2983 4217 2984 4328
rect 3034 4327 3035 4422
rect 2727 4329 2728 4422
rect 2983 4329 2984 4422
rect 3001 4217 3002 4330
rect 3076 4329 3077 4422
rect 2944 4217 2945 4332
rect 3001 4331 3002 4422
rect 3010 4217 3011 4332
rect 3022 4331 3023 4422
rect 3019 4217 3020 4334
rect 3082 4333 3083 4422
rect 3007 4217 3008 4336
rect 3019 4335 3020 4422
rect 3025 4217 3026 4336
rect 3088 4335 3089 4422
rect 3037 4217 3038 4338
rect 3079 4337 3080 4422
rect 3040 4217 3041 4340
rect 3139 4217 3140 4340
rect 3043 4341 3044 4422
rect 3157 4217 3158 4342
rect 3055 4217 3056 4344
rect 3091 4343 3092 4422
rect 3052 4217 3053 4346
rect 3055 4345 3056 4422
rect 2977 4217 2978 4348
rect 3052 4347 3053 4422
rect 2932 4217 2933 4350
rect 2977 4349 2978 4422
rect 2878 4217 2879 4352
rect 2932 4351 2933 4422
rect 3058 4217 3059 4352
rect 3184 4217 3185 4352
rect 3049 4217 3050 4354
rect 3058 4353 3059 4422
rect 2974 4217 2975 4356
rect 3049 4355 3050 4422
rect 2842 4217 2843 4358
rect 2974 4357 2975 4422
rect 3061 4217 3062 4358
rect 3094 4357 3095 4422
rect 3067 4217 3068 4360
rect 3139 4359 3140 4422
rect 3064 4361 3065 4422
rect 3067 4361 3068 4422
rect 3073 4217 3074 4362
rect 3278 4217 3279 4362
rect 3073 4363 3074 4422
rect 3115 4217 3116 4364
rect 3103 4217 3104 4366
rect 3121 4365 3122 4422
rect 3106 4217 3107 4368
rect 3124 4367 3125 4422
rect 3106 4369 3107 4422
rect 3206 4217 3207 4370
rect 3109 4217 3110 4372
rect 3157 4371 3158 4422
rect 3118 4373 3119 4422
rect 3257 4217 3258 4374
rect 3127 4217 3128 4376
rect 3184 4375 3185 4422
rect 3127 4377 3128 4422
rect 3267 4217 3268 4378
rect 3133 4379 3134 4422
rect 3281 4217 3282 4380
rect 3166 4217 3167 4382
rect 3205 4381 3206 4422
rect 3169 4217 3170 4384
rect 3326 4383 3327 4422
rect 3181 4385 3182 4422
rect 3221 4217 3222 4386
rect 3212 4217 3213 4388
rect 3218 4217 3219 4388
rect 2809 4389 2810 4422
rect 3217 4389 3218 4422
rect 3224 4217 3225 4390
rect 3260 4389 3261 4422
rect 3227 4217 3228 4392
rect 3263 4391 3264 4422
rect 3200 4217 3201 4394
rect 3226 4393 3227 4422
rect 3230 4217 3231 4394
rect 3266 4393 3267 4422
rect 3203 4217 3204 4396
rect 3229 4395 3230 4422
rect 3163 4217 3164 4398
rect 3202 4397 3203 4422
rect 3233 4217 3234 4398
rect 3269 4397 3270 4422
rect 3194 4217 3195 4400
rect 3232 4399 3233 4422
rect 3193 4401 3194 4422
rect 3370 4401 3371 4422
rect 3236 4217 3237 4404
rect 3291 4403 3292 4422
rect 3197 4217 3198 4406
rect 3235 4405 3236 4422
rect 3248 4217 3249 4406
rect 3315 4405 3316 4422
rect 3112 4407 3113 4422
rect 3248 4407 3249 4422
rect 3254 4217 3255 4408
rect 3306 4407 3307 4422
rect 3191 4217 3192 4410
rect 3254 4409 3255 4422
rect 3294 4409 3295 4422
rect 3329 4217 3330 4410
rect 3302 4217 3303 4412
rect 3319 4411 3320 4422
rect 3251 4217 3252 4414
rect 3303 4413 3304 4422
rect 3245 4217 3246 4416
rect 3251 4415 3252 4422
rect 3130 4217 3131 4418
rect 3245 4417 3246 4422
rect 3309 4217 3310 4418
rect 3347 4417 3348 4422
rect 3309 4419 3310 4422
rect 3343 4419 3344 4422
rect 3356 4419 3357 4422
rect 3367 4419 3368 4422
rect 2539 4426 2540 4429
rect 2749 4426 2750 4429
rect 2588 4430 2589 4667
rect 2899 4426 2900 4431
rect 2590 4426 2591 4433
rect 2959 4426 2960 4433
rect 2602 4434 2603 4667
rect 2778 4434 2779 4667
rect 2611 4426 2612 4437
rect 2615 4426 2616 4437
rect 2612 4438 2613 4667
rect 2947 4426 2948 4439
rect 2622 4426 2623 4441
rect 2682 4426 2683 4441
rect 2632 4426 2633 4443
rect 2908 4426 2909 4443
rect 2594 4426 2595 4445
rect 2907 4444 2908 4667
rect 2595 4446 2596 4667
rect 2706 4426 2707 4447
rect 2636 4426 2637 4449
rect 2925 4448 2926 4667
rect 2638 4450 2639 4667
rect 2953 4426 2954 4451
rect 2643 4426 2644 4453
rect 2860 4426 2861 4453
rect 2649 4454 2650 4667
rect 3052 4426 3053 4455
rect 2656 4456 2657 4667
rect 2835 4456 2836 4667
rect 2659 4458 2660 4667
rect 2848 4426 2849 4459
rect 2662 4460 2663 4667
rect 2667 4426 2668 4461
rect 2665 4462 2666 4667
rect 2709 4426 2710 4463
rect 2680 4464 2681 4667
rect 2983 4426 2984 4465
rect 2686 4466 2687 4667
rect 2950 4426 2951 4467
rect 2697 4426 2698 4469
rect 2821 4426 2822 4469
rect 2707 4470 2708 4667
rect 2730 4426 2731 4471
rect 2710 4472 2711 4667
rect 2962 4426 2963 4473
rect 2728 4474 2729 4667
rect 2735 4474 2736 4667
rect 2739 4426 2740 4475
rect 2941 4426 2942 4475
rect 2739 4476 2740 4667
rect 2998 4426 2999 4477
rect 2757 4478 2758 4667
rect 2800 4426 2801 4479
rect 2766 4480 2767 4667
rect 2776 4426 2777 4481
rect 2784 4480 2785 4667
rect 2827 4426 2828 4481
rect 2788 4426 2789 4483
rect 2790 4482 2791 4667
rect 2787 4484 2788 4667
rect 2830 4426 2831 4485
rect 2794 4426 2795 4487
rect 2805 4486 2806 4667
rect 2796 4488 2797 4667
rect 2857 4426 2858 4489
rect 2799 4490 2800 4667
rect 2992 4426 2993 4491
rect 2812 4426 2813 4493
rect 2889 4492 2890 4667
rect 2803 4426 2804 4495
rect 2811 4494 2812 4667
rect 2817 4494 2818 4667
rect 2872 4426 2873 4495
rect 2820 4496 2821 4667
rect 2839 4426 2840 4497
rect 2823 4498 2824 4667
rect 2956 4426 2957 4499
rect 2618 4426 2619 4501
rect 2955 4500 2956 4667
rect 2619 4502 2620 4667
rect 2764 4426 2765 4503
rect 2826 4502 2827 4667
rect 2866 4426 2867 4503
rect 2832 4504 2833 4667
rect 2845 4426 2846 4505
rect 2815 4426 2816 4507
rect 2844 4506 2845 4667
rect 2838 4508 2839 4667
rect 2851 4426 2852 4509
rect 2850 4510 2851 4667
rect 2893 4426 2894 4511
rect 2609 4512 2610 4667
rect 2892 4512 2893 4667
rect 2862 4514 2863 4667
rect 2887 4426 2888 4515
rect 2869 4426 2870 4517
rect 2895 4516 2896 4667
rect 2629 4426 2630 4519
rect 2868 4518 2869 4667
rect 2628 4520 2629 4667
rect 2688 4426 2689 4521
rect 2689 4522 2690 4667
rect 2914 4426 2915 4523
rect 2871 4524 2872 4667
rect 2917 4426 2918 4525
rect 2874 4526 2875 4667
rect 2932 4426 2933 4527
rect 2886 4528 2887 4667
rect 2905 4426 2906 4529
rect 2598 4530 2599 4667
rect 2904 4530 2905 4667
rect 2910 4530 2911 4667
rect 2977 4426 2978 4531
rect 2916 4532 2917 4667
rect 2971 4426 2972 4533
rect 2919 4534 2920 4667
rect 2974 4426 2975 4535
rect 2922 4536 2923 4667
rect 2989 4426 2990 4537
rect 2646 4426 2647 4539
rect 2988 4538 2989 4667
rect 2645 4540 2646 4667
rect 2934 4540 2935 4667
rect 2929 4426 2930 4543
rect 3129 4542 3130 4667
rect 2940 4544 2941 4667
rect 2995 4426 2996 4545
rect 2943 4546 2944 4667
rect 3001 4426 3002 4547
rect 2949 4548 2950 4667
rect 3013 4426 3014 4549
rect 2958 4550 2959 4667
rect 3016 4426 3017 4551
rect 2961 4552 2962 4667
rect 2965 4426 2966 4553
rect 2964 4554 2965 4667
rect 2986 4426 2987 4555
rect 2979 4556 2980 4667
rect 3031 4426 3032 4557
rect 2982 4558 2983 4667
rect 3034 4426 3035 4559
rect 2985 4560 2986 4667
rect 3049 4426 3050 4561
rect 2991 4562 2992 4667
rect 3019 4426 3020 4563
rect 2994 4564 2995 4667
rect 3022 4426 3023 4565
rect 3015 4566 3016 4667
rect 3076 4426 3077 4567
rect 3021 4568 3022 4667
rect 3067 4426 3068 4569
rect 3024 4570 3025 4667
rect 3079 4426 3080 4571
rect 3027 4572 3028 4667
rect 3055 4426 3056 4573
rect 3030 4574 3031 4667
rect 3043 4426 3044 4575
rect 3033 4576 3034 4667
rect 3082 4426 3083 4577
rect 3039 4578 3040 4667
rect 3088 4426 3089 4579
rect 3042 4580 3043 4667
rect 3091 4426 3092 4581
rect 3048 4582 3049 4667
rect 3121 4426 3122 4583
rect 3058 4426 3059 4585
rect 3241 4426 3242 4585
rect 3073 4426 3074 4587
rect 3141 4586 3142 4667
rect 3081 4588 3082 4667
rect 3214 4426 3215 4589
rect 3087 4590 3088 4667
rect 3124 4426 3125 4591
rect 3090 4592 3091 4667
rect 3094 4426 3095 4593
rect 3099 4592 3100 4667
rect 3127 4426 3128 4593
rect 3106 4426 3107 4595
rect 3245 4426 3246 4595
rect 3112 4426 3113 4597
rect 3150 4596 3151 4667
rect 3111 4598 3112 4667
rect 3282 4426 3283 4599
rect 3114 4600 3115 4667
rect 3244 4600 3245 4667
rect 3118 4426 3119 4603
rect 3120 4602 3121 4667
rect 3117 4604 3118 4667
rect 3254 4426 3255 4605
rect 3123 4606 3124 4667
rect 3263 4426 3264 4607
rect 3133 4426 3134 4609
rect 3256 4608 3257 4667
rect 3139 4426 3140 4611
rect 3271 4610 3272 4667
rect 3147 4612 3148 4667
rect 3181 4426 3182 4613
rect 3157 4426 3158 4615
rect 3241 4614 3242 4667
rect 3177 4616 3178 4667
rect 3235 4426 3236 4617
rect 3051 4618 3052 4667
rect 3235 4618 3236 4667
rect 3184 4426 3185 4621
rect 3187 4426 3188 4621
rect 3193 4426 3194 4621
rect 3363 4426 3364 4621
rect 3144 4622 3145 4667
rect 3192 4622 3193 4667
rect 3195 4622 3196 4667
rect 3202 4426 3203 4623
rect 3198 4624 3199 4667
rect 3205 4426 3206 4625
rect 3204 4626 3205 4667
rect 3238 4426 3239 4627
rect 3207 4628 3208 4667
rect 3269 4426 3270 4629
rect 3093 4630 3094 4667
rect 3268 4630 3269 4667
rect 3210 4632 3211 4667
rect 3226 4426 3227 4633
rect 3213 4634 3214 4667
rect 3229 4426 3230 4635
rect 3216 4636 3217 4667
rect 3232 4426 3233 4637
rect 3219 4638 3220 4667
rect 3321 4638 3322 4667
rect 3222 4640 3223 4667
rect 3329 4426 3330 4641
rect 3238 4642 3239 4667
rect 3312 4426 3313 4643
rect 3251 4426 3252 4645
rect 3315 4426 3316 4645
rect 3260 4426 3261 4647
rect 3262 4646 3263 4667
rect 3259 4648 3260 4667
rect 3340 4426 3341 4649
rect 3266 4426 3267 4651
rect 3314 4650 3315 4667
rect 3265 4652 3266 4667
rect 3291 4426 3292 4653
rect 3274 4654 3275 4667
rect 3303 4426 3304 4655
rect 3277 4656 3278 4667
rect 3347 4426 3348 4657
rect 3279 4426 3280 4659
rect 3283 4658 3284 4667
rect 3280 4660 3281 4667
rect 3309 4426 3310 4661
rect 3286 4662 3287 4667
rect 3306 4426 3307 4663
rect 3294 4426 3295 4665
rect 3337 4664 3338 4667
rect 2575 4673 2576 4888
rect 2784 4671 2785 4674
rect 2581 4671 2582 4676
rect 2707 4671 2708 4676
rect 2582 4677 2583 4888
rect 2778 4671 2779 4678
rect 2588 4671 2589 4680
rect 2874 4671 2875 4680
rect 2599 4681 2600 4888
rect 2750 4681 2751 4888
rect 2605 4671 2606 4684
rect 2925 4671 2926 4684
rect 2609 4671 2610 4686
rect 2799 4671 2800 4686
rect 2613 4687 2614 4888
rect 2686 4671 2687 4688
rect 2635 4671 2636 4690
rect 2873 4689 2874 4888
rect 2628 4671 2629 4692
rect 2635 4691 2636 4888
rect 2642 4671 2643 4692
rect 2868 4671 2869 4692
rect 2645 4671 2646 4694
rect 2783 4693 2784 4888
rect 2649 4671 2650 4696
rect 2820 4671 2821 4696
rect 2652 4697 2653 4888
rect 2949 4671 2950 4698
rect 2655 4699 2656 4888
rect 2662 4671 2663 4700
rect 2664 4699 2665 4888
rect 2665 4671 2666 4700
rect 2667 4699 2668 4888
rect 2895 4671 2896 4700
rect 2680 4671 2681 4702
rect 2961 4671 2962 4702
rect 2679 4703 2680 4888
rect 2683 4671 2684 4704
rect 2686 4703 2687 4888
rect 2698 4703 2699 4888
rect 2692 4671 2693 4706
rect 2985 4671 2986 4706
rect 2692 4707 2693 4888
rect 2710 4671 2711 4708
rect 2707 4709 2708 4888
rect 2787 4671 2788 4710
rect 2710 4711 2711 4888
rect 2757 4671 2758 4712
rect 2713 4713 2714 4888
rect 2982 4671 2983 4714
rect 2723 4715 2724 4888
rect 2940 4671 2941 4716
rect 2725 4671 2726 4718
rect 2979 4671 2980 4718
rect 2616 4671 2617 4720
rect 2726 4719 2727 4888
rect 2617 4721 2618 4888
rect 2892 4671 2893 4722
rect 2735 4671 2736 4724
rect 3125 4723 3126 4888
rect 2739 4671 2740 4726
rect 2898 4671 2899 4726
rect 2747 4727 2748 4888
rect 2817 4671 2818 4728
rect 2766 4671 2767 4730
rect 2768 4729 2769 4888
rect 2774 4729 2775 4888
rect 2790 4671 2791 4730
rect 2780 4731 2781 4888
rect 2826 4671 2827 4732
rect 2792 4733 2793 4888
rect 2832 4671 2833 4734
rect 2798 4735 2799 4888
rect 2838 4671 2839 4736
rect 2805 4671 2806 4738
rect 2819 4737 2820 4888
rect 2804 4739 2805 4888
rect 2850 4671 2851 4740
rect 2810 4741 2811 4888
rect 2811 4671 2812 4742
rect 2816 4741 2817 4888
rect 2844 4671 2845 4742
rect 2649 4743 2650 4888
rect 2843 4743 2844 4888
rect 2823 4671 2824 4746
rect 3310 4671 3311 4746
rect 2828 4747 2829 4888
rect 2904 4671 2905 4748
rect 2661 4749 2662 4888
rect 2903 4749 2904 4888
rect 2831 4751 2832 4888
rect 2907 4671 2908 4752
rect 2837 4753 2838 4888
rect 2964 4671 2965 4754
rect 2840 4755 2841 4888
rect 2922 4671 2923 4756
rect 2849 4757 2850 4888
rect 2916 4671 2917 4758
rect 2732 4671 2733 4760
rect 2915 4759 2916 4888
rect 2732 4761 2733 4888
rect 2796 4671 2797 4762
rect 2795 4763 2796 4888
rect 2835 4671 2836 4764
rect 2834 4765 2835 4888
rect 2862 4671 2863 4766
rect 2852 4767 2853 4888
rect 2919 4671 2920 4768
rect 2855 4769 2856 4888
rect 2910 4671 2911 4770
rect 2861 4771 2862 4888
rect 2934 4671 2935 4772
rect 2867 4773 2868 4888
rect 2943 4671 2944 4774
rect 2871 4671 2872 4776
rect 2876 4775 2877 4888
rect 2879 4775 2880 4888
rect 2955 4671 2956 4776
rect 2882 4777 2883 4888
rect 2958 4671 2959 4778
rect 2886 4671 2887 4780
rect 2891 4779 2892 4888
rect 2889 4671 2890 4782
rect 2918 4781 2919 4888
rect 2897 4783 2898 4888
rect 2951 4783 2952 4888
rect 2901 4671 2902 4786
rect 2966 4785 2967 4888
rect 2909 4787 2910 4888
rect 2988 4671 2989 4788
rect 2912 4789 2913 4888
rect 3068 4789 3069 4888
rect 2927 4791 2928 4888
rect 2994 4671 2995 4792
rect 2930 4793 2931 4888
rect 2991 4671 2992 4794
rect 2933 4795 2934 4888
rect 3015 4671 3016 4796
rect 2939 4797 2940 4888
rect 3021 4671 3022 4798
rect 2957 4799 2958 4888
rect 3033 4671 3034 4800
rect 2728 4671 2729 4802
rect 3032 4801 3033 4888
rect 2963 4803 2964 4888
rect 3024 4671 3025 4804
rect 2969 4805 2970 4888
rect 3039 4671 3040 4806
rect 2975 4807 2976 4888
rect 3120 4671 3121 4808
rect 2978 4809 2979 4888
rect 3045 4671 3046 4810
rect 2990 4811 2991 4888
rect 3027 4671 3028 4812
rect 2996 4813 2997 4888
rect 3081 4671 3082 4814
rect 3002 4815 3003 4888
rect 3165 4671 3166 4816
rect 3014 4817 3015 4888
rect 3099 4671 3100 4818
rect 3030 4671 3031 4820
rect 3035 4819 3036 4888
rect 3038 4819 3039 4888
rect 3111 4671 3112 4820
rect 3042 4671 3043 4822
rect 3080 4821 3081 4888
rect 3041 4823 3042 4888
rect 3123 4671 3124 4824
rect 3047 4825 3048 4888
rect 3051 4671 3052 4826
rect 3065 4825 3066 4888
rect 3087 4671 3088 4826
rect 3083 4827 3084 4888
rect 3131 4827 3132 4888
rect 3098 4829 3099 4888
rect 3147 4671 3148 4830
rect 3101 4831 3102 4888
rect 3150 4671 3151 4832
rect 3104 4833 3105 4888
rect 3195 4671 3196 4834
rect 3090 4671 3091 4836
rect 3194 4835 3195 4888
rect 3107 4837 3108 4888
rect 3198 4671 3199 4838
rect 3110 4839 3111 4888
rect 3192 4671 3193 4840
rect 3114 4671 3115 4842
rect 3253 4671 3254 4842
rect 3113 4843 3114 4888
rect 3144 4671 3145 4844
rect 3020 4845 3021 4888
rect 3143 4845 3144 4888
rect 3117 4671 3118 4848
rect 3235 4671 3236 4848
rect 3000 4671 3001 4850
rect 3116 4849 3117 4888
rect 3122 4849 3123 4888
rect 3207 4671 3208 4850
rect 3129 4671 3130 4852
rect 3156 4851 3157 4888
rect 3128 4853 3129 4888
rect 3216 4671 3217 4854
rect 3137 4855 3138 4888
rect 3222 4671 3223 4856
rect 3141 4671 3142 4858
rect 3189 4671 3190 4858
rect 3134 4859 3135 4888
rect 3140 4859 3141 4888
rect 3153 4859 3154 4888
rect 3210 4671 3211 4860
rect 3165 4861 3166 4888
rect 3201 4671 3202 4862
rect 3093 4671 3094 4864
rect 3200 4863 3201 4888
rect 3177 4671 3178 4866
rect 3293 4671 3294 4866
rect 3182 4867 3183 4888
rect 3213 4671 3214 4868
rect 3185 4869 3186 4888
rect 3259 4671 3260 4870
rect 3188 4871 3189 4888
rect 3262 4671 3263 4872
rect 3197 4873 3198 4888
rect 3274 4671 3275 4874
rect 3206 4875 3207 4888
rect 3280 4671 3281 4876
rect 3209 4877 3210 4888
rect 3283 4671 3284 4878
rect 3219 4671 3220 4880
rect 3296 4671 3297 4880
rect 3238 4671 3239 4882
rect 3256 4671 3257 4882
rect 3265 4671 3266 4882
rect 3334 4671 3335 4882
rect 3277 4671 3278 4884
rect 3328 4671 3329 4884
rect 3289 4671 3290 4886
rect 3300 4671 3301 4886
rect 3343 4671 3344 4886
rect 3350 4671 3351 4886
rect 2570 4894 2571 5073
rect 2703 4894 2704 5073
rect 2582 4892 2583 4897
rect 2831 4892 2832 4897
rect 2589 4892 2590 4899
rect 2804 4892 2805 4899
rect 2593 4900 2594 5073
rect 2846 4900 2847 5073
rect 2596 4892 2597 4903
rect 2664 4892 2665 4903
rect 2597 4904 2598 5073
rect 2620 4904 2621 5073
rect 2600 4906 2601 5073
rect 2840 4892 2841 4907
rect 2603 4892 2604 4909
rect 2667 4892 2668 4909
rect 2611 4910 2612 5073
rect 2780 4892 2781 4911
rect 2617 4912 2618 5073
rect 2783 4892 2784 4913
rect 2623 4914 2624 5073
rect 2864 4914 2865 5073
rect 2635 4916 2636 5073
rect 2642 4892 2643 4917
rect 2638 4892 2639 4919
rect 2658 4892 2659 4919
rect 2606 4892 2607 4921
rect 2638 4920 2639 5073
rect 2641 4920 2642 5073
rect 2655 4892 2656 4921
rect 2647 4922 2648 5073
rect 2879 4892 2880 4923
rect 2661 4892 2662 4925
rect 2861 4892 2862 4925
rect 2654 4926 2655 5073
rect 2861 4926 2862 5073
rect 2663 4928 2664 5073
rect 2894 4928 2895 5073
rect 2666 4930 2667 5073
rect 2789 4930 2790 5073
rect 2675 4932 2676 5073
rect 2692 4892 2693 4933
rect 2681 4934 2682 5073
rect 2798 4892 2799 4935
rect 2707 4892 2708 4937
rect 2735 4936 2736 5073
rect 2719 4938 2720 5073
rect 2732 4892 2733 4939
rect 2575 4892 2576 4941
rect 2732 4940 2733 5073
rect 2576 4942 2577 5073
rect 2583 4942 2584 5073
rect 2738 4942 2739 5073
rect 2747 4892 2748 4943
rect 2604 4944 2605 5073
rect 2747 4944 2748 5073
rect 2741 4946 2742 5073
rect 2750 4892 2751 4947
rect 2744 4892 2745 4949
rect 2915 4892 2916 4949
rect 2689 4892 2690 4951
rect 2915 4950 2916 5073
rect 2688 4952 2689 5073
rect 2912 4892 2913 4953
rect 2723 4892 2724 4955
rect 2912 4954 2913 5073
rect 2753 4956 2754 5073
rect 2876 4892 2877 4957
rect 2765 4958 2766 5073
rect 2768 4892 2769 4959
rect 2771 4958 2772 5073
rect 2774 4892 2775 4959
rect 2777 4958 2778 5073
rect 2792 4892 2793 4959
rect 2795 4892 2796 4959
rect 2897 4958 2898 5073
rect 2795 4960 2796 5073
rect 2810 4892 2811 4961
rect 2807 4962 2808 5073
rect 2816 4892 2817 4963
rect 2810 4964 2811 5073
rect 2819 4892 2820 4965
rect 2679 4892 2680 4967
rect 2819 4966 2820 5073
rect 2813 4968 2814 5073
rect 2834 4892 2835 4969
rect 2825 4970 2826 5073
rect 2843 4892 2844 4971
rect 2828 4892 2829 4973
rect 2843 4972 2844 5073
rect 2831 4974 2832 5073
rect 2855 4892 2856 4975
rect 2651 4976 2652 5073
rect 2855 4976 2856 5073
rect 2849 4976 2850 5073
rect 2849 4892 2850 4977
rect 2852 4892 2853 4979
rect 2858 4978 2859 5073
rect 2870 4978 2871 5073
rect 2891 4892 2892 4979
rect 2607 4980 2608 5073
rect 2891 4980 2892 5073
rect 2873 4892 2874 4983
rect 2888 4982 2889 5073
rect 2882 4892 2883 4985
rect 2885 4984 2886 5073
rect 2867 4892 2868 4987
rect 2882 4986 2883 5073
rect 2613 4892 2614 4989
rect 2867 4988 2868 5073
rect 2614 4990 2615 5073
rect 2726 4892 2727 4991
rect 2900 4990 2901 5073
rect 2903 4892 2904 4991
rect 2903 4992 2904 5073
rect 2909 4892 2910 4993
rect 2921 4992 2922 5073
rect 2927 4892 2928 4993
rect 2726 4994 2727 5073
rect 2927 4994 2928 5073
rect 2939 4892 2940 4995
rect 2945 4994 2946 5073
rect 2939 4996 2940 5073
rect 2966 4892 2967 4997
rect 2969 4892 2970 4997
rect 2981 4996 2982 5073
rect 2957 4892 2958 4999
rect 2969 4998 2970 5073
rect 2951 4892 2952 5001
rect 2957 5000 2958 5073
rect 2933 4892 2934 5003
rect 2951 5002 2952 5073
rect 2975 4892 2976 5003
rect 2993 5002 2994 5073
rect 2930 4892 2931 5005
rect 2975 5004 2976 5073
rect 2918 4892 2919 5007
rect 2930 5006 2931 5073
rect 2837 4892 2838 5009
rect 2918 5008 2919 5073
rect 2987 5008 2988 5073
rect 3116 4892 3117 5009
rect 2990 4892 2991 5011
rect 3026 5010 3027 5073
rect 2996 4892 2997 5013
rect 3008 5012 3009 5073
rect 2978 4892 2979 5015
rect 2996 5014 2997 5073
rect 2933 5016 2934 5073
rect 2978 5016 2979 5073
rect 3020 4892 3021 5017
rect 3071 4892 3072 5017
rect 3020 5018 3021 5073
rect 3194 4892 3195 5019
rect 2710 4892 2711 5021
rect 3195 5020 3196 5073
rect 3023 5022 3024 5073
rect 3032 4892 3033 5023
rect 3035 4892 3036 5023
rect 3140 5022 3141 5073
rect 3035 5024 3036 5073
rect 3125 4892 3126 5025
rect 3038 4892 3039 5027
rect 3177 5026 3178 5073
rect 3041 4892 3042 5029
rect 3183 5028 3184 5073
rect 3047 4892 3048 5031
rect 3056 5030 3057 5073
rect 3047 5032 3048 5073
rect 3065 4892 3066 5033
rect 3068 5032 3069 5073
rect 3107 4892 3108 5033
rect 3071 5034 3072 5073
rect 3203 4892 3204 5035
rect 3080 4892 3081 5037
rect 3089 5036 3090 5073
rect 2963 4892 2964 5039
rect 3080 5038 3081 5073
rect 2695 4892 2696 5041
rect 2963 5040 2964 5073
rect 3083 4892 3084 5041
rect 3092 5040 3093 5073
rect 3095 5040 3096 5073
rect 3098 4892 3099 5041
rect 3098 5042 3099 5073
rect 3101 4892 3102 5043
rect 3104 4892 3105 5043
rect 3214 5042 3215 5073
rect 3107 5044 3108 5073
rect 3110 4892 3111 5045
rect 3110 5046 3111 5073
rect 3113 4892 3114 5047
rect 3122 4892 3123 5047
rect 3134 5046 3135 5073
rect 3128 4892 3129 5049
rect 3212 4892 3213 5049
rect 3131 5050 3132 5073
rect 3233 4892 3234 5051
rect 3119 5052 3120 5073
rect 3232 5052 3233 5073
rect 3143 5054 3144 5073
rect 3239 5054 3240 5073
rect 3153 4892 3154 5057
rect 3161 5056 3162 5073
rect 3137 4892 3138 5059
rect 3152 5058 3153 5073
rect 3077 5060 3078 5073
rect 3137 5060 3138 5073
rect 3156 4892 3157 5061
rect 3164 5060 3165 5073
rect 2936 5062 2937 5073
rect 3155 5062 3156 5073
rect 3180 5062 3181 5073
rect 3185 4892 3186 5063
rect 3188 4892 3189 5063
rect 3256 4892 3257 5063
rect 3192 5064 3193 5073
rect 3197 4892 3198 5065
rect 3209 4892 3210 5065
rect 3253 5064 3254 5073
rect 3206 4892 3207 5067
rect 3208 5066 3209 5073
rect 3014 4892 3015 5069
rect 3205 5068 3206 5073
rect 3002 4892 3003 5071
rect 3014 5070 3015 5073
rect 2563 5077 2564 5080
rect 2774 5079 2775 5266
rect 2586 5077 2587 5082
rect 2590 5077 2591 5082
rect 2593 5077 2594 5082
rect 2741 5077 2742 5082
rect 2593 5083 2594 5266
rect 2951 5077 2952 5084
rect 2596 5085 2597 5266
rect 2867 5077 2868 5086
rect 2604 5077 2605 5088
rect 2852 5087 2853 5266
rect 2603 5089 2604 5266
rect 2843 5077 2844 5090
rect 2607 5077 2608 5092
rect 2638 5077 2639 5092
rect 2617 5077 2618 5094
rect 2620 5093 2621 5266
rect 2623 5077 2624 5094
rect 2915 5077 2916 5094
rect 2629 5095 2630 5266
rect 2641 5077 2642 5096
rect 2638 5097 2639 5266
rect 2891 5077 2892 5098
rect 2642 5099 2643 5266
rect 2882 5077 2883 5100
rect 2645 5101 2646 5266
rect 2647 5077 2648 5102
rect 2651 5077 2652 5102
rect 2897 5077 2898 5102
rect 2661 5103 2662 5266
rect 2675 5077 2676 5104
rect 2664 5105 2665 5266
rect 2894 5077 2895 5106
rect 2666 5077 2667 5108
rect 2837 5107 2838 5266
rect 2671 5109 2672 5266
rect 2771 5077 2772 5110
rect 2678 5077 2679 5112
rect 2819 5077 2820 5112
rect 2632 5077 2633 5114
rect 2819 5113 2820 5266
rect 2632 5115 2633 5266
rect 2846 5077 2847 5116
rect 2678 5117 2679 5266
rect 2714 5117 2715 5266
rect 2681 5077 2682 5120
rect 2870 5077 2871 5120
rect 2681 5121 2682 5266
rect 2900 5077 2901 5122
rect 2697 5123 2698 5266
rect 2703 5077 2704 5124
rect 2707 5123 2708 5266
rect 2726 5077 2727 5124
rect 2717 5125 2718 5266
rect 2891 5125 2892 5266
rect 2720 5127 2721 5266
rect 2732 5077 2733 5128
rect 2723 5129 2724 5266
rect 2735 5077 2736 5130
rect 2729 5077 2730 5132
rect 2930 5077 2931 5132
rect 2732 5133 2733 5266
rect 2738 5077 2739 5134
rect 2735 5135 2736 5266
rect 2753 5077 2754 5136
rect 2674 5137 2675 5266
rect 2753 5137 2754 5266
rect 2747 5077 2748 5140
rect 2876 5139 2877 5266
rect 2747 5141 2748 5266
rect 2765 5077 2766 5142
rect 2765 5143 2766 5266
rect 2795 5077 2796 5144
rect 2771 5145 2772 5266
rect 2777 5077 2778 5146
rect 2777 5147 2778 5266
rect 2789 5077 2790 5148
rect 2783 5149 2784 5266
rect 2807 5077 2808 5150
rect 2786 5151 2787 5266
rect 2810 5077 2811 5152
rect 2801 5153 2802 5266
rect 2825 5077 2826 5154
rect 2807 5155 2808 5266
rect 2831 5077 2832 5156
rect 2810 5157 2811 5266
rect 2885 5077 2886 5158
rect 2813 5157 2814 5266
rect 2813 5077 2814 5158
rect 2816 5159 2817 5266
rect 2918 5077 2919 5160
rect 2825 5161 2826 5266
rect 3077 5077 3078 5162
rect 2831 5163 2832 5266
rect 2849 5077 2850 5164
rect 2849 5165 2850 5266
rect 2864 5077 2865 5166
rect 2855 5165 2856 5266
rect 2855 5077 2856 5166
rect 2858 5165 2859 5266
rect 2858 5077 2859 5166
rect 2861 5165 2862 5266
rect 2861 5077 2862 5166
rect 2864 5167 2865 5266
rect 3080 5077 3081 5168
rect 2870 5169 2871 5266
rect 2903 5077 2904 5170
rect 2873 5171 2874 5266
rect 2888 5077 2889 5172
rect 2897 5171 2898 5266
rect 2933 5077 2934 5172
rect 2900 5173 2901 5266
rect 2936 5077 2937 5174
rect 2903 5175 2904 5266
rect 2984 5175 2985 5266
rect 2909 5177 2910 5266
rect 2927 5077 2928 5178
rect 2912 5077 2913 5180
rect 2915 5179 2916 5266
rect 2703 5181 2704 5266
rect 2912 5181 2913 5266
rect 2918 5181 2919 5266
rect 2939 5077 2940 5182
rect 2921 5077 2922 5184
rect 2978 5077 2979 5184
rect 2924 5185 2925 5266
rect 2957 5077 2958 5186
rect 2930 5187 2931 5266
rect 2945 5077 2946 5188
rect 2933 5189 2934 5266
rect 3116 5077 3117 5190
rect 2936 5191 2937 5266
rect 2987 5077 2988 5192
rect 2942 5193 2943 5266
rect 2969 5077 2970 5194
rect 2948 5195 2949 5266
rect 2981 5077 2982 5196
rect 2960 5197 2961 5266
rect 3023 5077 3024 5198
rect 2963 5077 2964 5200
rect 3137 5077 3138 5200
rect 2963 5201 2964 5266
rect 2996 5077 2997 5202
rect 2966 5203 2967 5266
rect 3177 5077 3178 5204
rect 2987 5205 2988 5266
rect 3056 5077 3057 5206
rect 2999 5207 3000 5266
rect 3092 5077 3093 5208
rect 3002 5209 3003 5266
rect 3014 5077 3015 5210
rect 3008 5077 3009 5212
rect 3014 5211 3015 5266
rect 3011 5213 3012 5266
rect 3164 5077 3165 5214
rect 3017 5215 3018 5266
rect 3068 5077 3069 5216
rect 3020 5077 3021 5218
rect 3205 5077 3206 5218
rect 3026 5077 3027 5220
rect 3158 5077 3159 5220
rect 3032 5221 3033 5266
rect 3107 5077 3108 5222
rect 3035 5077 3036 5224
rect 3067 5223 3068 5266
rect 3035 5225 3036 5266
rect 3071 5077 3072 5226
rect 3038 5227 3039 5266
rect 3095 5077 3096 5228
rect 3047 5077 3048 5230
rect 3174 5077 3175 5230
rect 2993 5077 2994 5232
rect 3048 5231 3049 5266
rect 3064 5231 3065 5266
rect 3119 5077 3120 5232
rect 3070 5233 3071 5266
rect 3086 5233 3087 5266
rect 3073 5235 3074 5266
rect 3083 5235 3084 5266
rect 3089 5077 3090 5236
rect 3146 5077 3147 5236
rect 3095 5237 3096 5266
rect 3161 5077 3162 5238
rect 3098 5077 3099 5240
rect 3202 5077 3203 5240
rect 3105 5241 3106 5266
rect 3262 5077 3263 5242
rect 3108 5243 3109 5266
rect 3180 5077 3181 5244
rect 3110 5077 3111 5246
rect 3170 5077 3171 5246
rect 3089 5247 3090 5266
rect 3170 5247 3171 5266
rect 3111 5249 3112 5266
rect 3183 5077 3184 5250
rect 3120 5251 3121 5266
rect 3192 5077 3193 5252
rect 3123 5253 3124 5266
rect 3152 5077 3153 5254
rect 3131 5077 3132 5256
rect 3235 5077 3236 5256
rect 3134 5077 3135 5258
rect 3232 5077 3233 5258
rect 3140 5259 3141 5266
rect 3246 5077 3247 5260
rect 3143 5077 3144 5262
rect 3253 5077 3254 5262
rect 3164 5263 3165 5266
rect 3208 5077 3209 5264
rect 2576 5270 2577 5273
rect 2720 5270 2721 5273
rect 2573 5274 2574 5443
rect 2576 5274 2577 5443
rect 2605 5274 2606 5443
rect 2629 5270 2630 5275
rect 2610 5270 2611 5277
rect 2849 5270 2850 5277
rect 2617 5270 2618 5279
rect 2620 5270 2621 5279
rect 2623 5270 2624 5279
rect 2664 5278 2665 5443
rect 2626 5270 2627 5281
rect 2831 5270 2832 5281
rect 2632 5270 2633 5283
rect 2635 5282 2636 5443
rect 2632 5284 2633 5443
rect 2876 5270 2877 5285
rect 2638 5286 2639 5443
rect 2810 5270 2811 5287
rect 2625 5288 2626 5443
rect 2811 5288 2812 5443
rect 2649 5270 2650 5291
rect 2753 5270 2754 5291
rect 2655 5292 2656 5443
rect 3120 5270 3121 5293
rect 2661 5270 2662 5295
rect 2688 5270 2689 5295
rect 2569 5270 2570 5297
rect 2689 5296 2690 5443
rect 2570 5298 2571 5443
rect 2774 5270 2775 5299
rect 2671 5270 2672 5301
rect 2747 5270 2748 5301
rect 2641 5302 2642 5443
rect 2748 5302 2749 5443
rect 2671 5304 2672 5443
rect 2692 5304 2693 5443
rect 2674 5270 2675 5307
rect 2816 5270 2817 5307
rect 2677 5308 2678 5443
rect 2723 5270 2724 5309
rect 2681 5270 2682 5311
rect 2870 5270 2871 5311
rect 2683 5312 2684 5443
rect 2765 5270 2766 5313
rect 2686 5314 2687 5443
rect 2697 5270 2698 5315
rect 2695 5316 2696 5443
rect 2732 5270 2733 5317
rect 2704 5318 2705 5443
rect 2735 5270 2736 5319
rect 2717 5270 2718 5321
rect 2900 5270 2901 5321
rect 2680 5322 2681 5443
rect 2717 5322 2718 5443
rect 2720 5322 2721 5443
rect 2835 5322 2836 5443
rect 2724 5324 2725 5443
rect 2871 5324 2872 5443
rect 2736 5326 2737 5443
rect 2783 5270 2784 5327
rect 2739 5328 2740 5443
rect 2786 5270 2787 5329
rect 2751 5330 2752 5443
rect 2771 5270 2772 5331
rect 2760 5332 2761 5443
rect 2777 5270 2778 5333
rect 2766 5334 2767 5443
rect 2868 5334 2869 5443
rect 2769 5336 2770 5443
rect 2918 5270 2919 5337
rect 2784 5338 2785 5443
rect 2807 5270 2808 5339
rect 2787 5340 2788 5443
rect 2801 5270 2802 5341
rect 2790 5342 2791 5443
rect 2819 5270 2820 5343
rect 2796 5344 2797 5443
rect 2837 5270 2838 5345
rect 2802 5346 2803 5443
rect 2855 5270 2856 5347
rect 2808 5348 2809 5443
rect 2852 5270 2853 5349
rect 2813 5270 2814 5351
rect 2817 5350 2818 5443
rect 2814 5352 2815 5443
rect 2858 5270 2859 5353
rect 2820 5354 2821 5443
rect 2861 5270 2862 5355
rect 2823 5356 2824 5443
rect 2873 5270 2874 5357
rect 2700 5270 2701 5359
rect 2874 5358 2875 5443
rect 2825 5270 2826 5361
rect 2984 5270 2985 5361
rect 2629 5362 2630 5443
rect 2826 5362 2827 5443
rect 2841 5362 2842 5443
rect 2891 5270 2892 5363
rect 2847 5364 2848 5443
rect 2915 5270 2916 5365
rect 2850 5366 2851 5443
rect 2903 5270 2904 5367
rect 2856 5368 2857 5443
rect 2897 5270 2898 5369
rect 2862 5370 2863 5443
rect 2909 5270 2910 5371
rect 2864 5270 2865 5373
rect 2981 5270 2982 5373
rect 2710 5270 2711 5375
rect 2865 5374 2866 5443
rect 2877 5374 2878 5443
rect 3009 5374 3010 5443
rect 2880 5376 2881 5443
rect 2930 5270 2931 5377
rect 2883 5378 2884 5443
rect 2933 5270 2934 5379
rect 2886 5380 2887 5443
rect 2924 5270 2925 5381
rect 2892 5382 2893 5443
rect 2942 5270 2943 5383
rect 2898 5384 2899 5443
rect 2936 5270 2937 5385
rect 2910 5386 2911 5443
rect 2960 5270 2961 5387
rect 2922 5388 2923 5443
rect 2999 5270 3000 5389
rect 2912 5270 2913 5391
rect 2999 5390 3000 5443
rect 2913 5392 2914 5443
rect 2963 5270 2964 5393
rect 2925 5394 2926 5443
rect 3002 5270 3003 5395
rect 2934 5396 2935 5443
rect 2987 5270 2988 5397
rect 2940 5398 2941 5443
rect 3035 5270 3036 5399
rect 2946 5400 2947 5443
rect 3037 5400 3038 5443
rect 2948 5270 2949 5403
rect 3002 5402 3003 5443
rect 2955 5404 2956 5443
rect 3067 5270 3068 5405
rect 2958 5406 2959 5443
rect 3011 5270 3012 5407
rect 2961 5408 2962 5443
rect 3014 5270 3015 5409
rect 2964 5410 2965 5443
rect 3017 5270 3018 5411
rect 2966 5270 2967 5413
rect 3048 5270 3049 5413
rect 2979 5414 2980 5443
rect 3032 5270 3033 5415
rect 2982 5416 2983 5443
rect 3045 5270 3046 5417
rect 3026 5270 3027 5419
rect 3154 5270 3155 5419
rect 3040 5420 3041 5443
rect 3147 5270 3148 5421
rect 3043 5422 3044 5443
rect 3089 5270 3090 5423
rect 3052 5424 3053 5443
rect 3108 5270 3109 5425
rect 3055 5270 3056 5427
rect 3076 5270 3077 5427
rect 3055 5428 3056 5443
rect 3111 5270 3112 5429
rect 3061 5430 3062 5443
rect 3143 5270 3144 5431
rect 3064 5270 3065 5433
rect 3140 5270 3141 5433
rect 3070 5270 3071 5435
rect 3102 5270 3103 5435
rect 3073 5270 3074 5437
rect 3079 5270 3080 5437
rect 3085 5436 3086 5443
rect 3123 5270 3124 5437
rect 3088 5438 3089 5443
rect 3170 5270 3171 5439
rect 3105 5270 3106 5441
rect 3167 5270 3168 5441
rect 2563 5447 2564 5450
rect 2576 5447 2577 5450
rect 2563 5451 2564 5600
rect 2566 5447 2567 5452
rect 2566 5453 2567 5600
rect 2605 5447 2606 5454
rect 2570 5447 2571 5456
rect 2686 5447 2687 5456
rect 2573 5447 2574 5458
rect 2689 5447 2690 5458
rect 2575 5459 2576 5600
rect 2582 5459 2583 5600
rect 2596 5447 2597 5460
rect 2635 5447 2636 5460
rect 2611 5447 2612 5462
rect 2638 5447 2639 5462
rect 2615 5463 2616 5600
rect 2823 5447 2824 5464
rect 2618 5447 2619 5466
rect 2702 5465 2703 5600
rect 2622 5447 2623 5468
rect 2802 5447 2803 5468
rect 2625 5447 2626 5470
rect 2796 5447 2797 5470
rect 2632 5447 2633 5472
rect 2650 5471 2651 5600
rect 2644 5473 2645 5600
rect 2677 5447 2678 5474
rect 2648 5447 2649 5476
rect 2820 5447 2821 5476
rect 2653 5477 2654 5600
rect 2695 5447 2696 5478
rect 2662 5479 2663 5600
rect 2771 5479 2772 5600
rect 2667 5447 2668 5482
rect 2692 5447 2693 5482
rect 2674 5447 2675 5484
rect 2710 5447 2711 5484
rect 2679 5485 2680 5600
rect 2736 5447 2737 5486
rect 2683 5447 2684 5488
rect 2739 5447 2740 5488
rect 2686 5489 2687 5600
rect 2795 5489 2796 5600
rect 2693 5491 2694 5600
rect 2883 5447 2884 5492
rect 2704 5447 2705 5494
rect 2720 5447 2721 5494
rect 2705 5495 2706 5600
rect 2748 5447 2749 5496
rect 2612 5497 2613 5600
rect 2747 5497 2748 5600
rect 2708 5499 2709 5600
rect 2751 5447 2752 5500
rect 2711 5501 2712 5600
rect 2865 5447 2866 5502
rect 2714 5503 2715 5600
rect 2760 5447 2761 5504
rect 2738 5505 2739 5600
rect 2808 5447 2809 5506
rect 2741 5507 2742 5600
rect 2784 5447 2785 5508
rect 2744 5509 2745 5600
rect 2787 5447 2788 5510
rect 2750 5511 2751 5600
rect 2811 5447 2812 5512
rect 2753 5513 2754 5600
rect 2814 5447 2815 5514
rect 2756 5515 2757 5600
rect 2790 5447 2791 5516
rect 2759 5517 2760 5600
rect 2826 5447 2827 5518
rect 2762 5519 2763 5600
rect 2862 5447 2863 5520
rect 2766 5447 2767 5522
rect 2847 5447 2848 5522
rect 2765 5523 2766 5600
rect 2880 5447 2881 5524
rect 2769 5447 2770 5526
rect 2856 5447 2857 5526
rect 2768 5527 2769 5600
rect 2817 5447 2818 5528
rect 2780 5529 2781 5600
rect 2835 5447 2836 5530
rect 2786 5531 2787 5600
rect 2841 5447 2842 5532
rect 2792 5533 2793 5600
rect 2850 5447 2851 5534
rect 2801 5535 2802 5600
rect 2910 5447 2911 5536
rect 2804 5537 2805 5600
rect 2868 5447 2869 5538
rect 2807 5539 2808 5600
rect 2871 5447 2872 5540
rect 2822 5541 2823 5600
rect 2967 5447 2968 5542
rect 2825 5543 2826 5600
rect 2886 5447 2887 5544
rect 2828 5545 2829 5600
rect 2992 5447 2993 5546
rect 2834 5547 2835 5600
rect 2925 5447 2926 5548
rect 2837 5549 2838 5600
rect 2922 5447 2923 5550
rect 2840 5551 2841 5600
rect 2892 5447 2893 5552
rect 2843 5553 2844 5600
rect 2913 5447 2914 5554
rect 2846 5555 2847 5600
rect 2919 5555 2920 5600
rect 2852 5557 2853 5600
rect 2891 5557 2892 5600
rect 2864 5559 2865 5600
rect 2934 5447 2935 5560
rect 2882 5561 2883 5600
rect 2982 5447 2983 5562
rect 2885 5563 2886 5600
rect 2940 5447 2941 5564
rect 2888 5565 2889 5600
rect 2964 5447 2965 5566
rect 2898 5447 2899 5568
rect 2995 5447 2996 5568
rect 2849 5569 2850 5600
rect 2898 5569 2899 5600
rect 2901 5569 2902 5600
rect 2985 5447 2986 5570
rect 2910 5571 2911 5600
rect 2923 5571 2924 5600
rect 2913 5573 2914 5600
rect 2933 5573 2934 5600
rect 2930 5575 2931 5600
rect 2961 5447 2962 5576
rect 2937 5577 2938 5600
rect 2946 5447 2947 5578
rect 2947 5579 2948 5600
rect 3040 5447 3041 5580
rect 2955 5447 2956 5582
rect 2960 5581 2961 5600
rect 2958 5447 2959 5584
rect 3013 5447 3014 5584
rect 2957 5585 2958 5600
rect 3058 5447 3059 5586
rect 2969 5587 2970 5600
rect 3094 5447 3095 5588
rect 2972 5589 2973 5600
rect 3052 5447 3053 5590
rect 2975 5591 2976 5600
rect 3055 5447 3056 5592
rect 2979 5447 2980 5594
rect 3002 5447 3003 5594
rect 3014 5593 3015 5600
rect 3018 5593 3019 5600
rect 3027 5593 3028 5600
rect 3085 5447 3086 5594
rect 3043 5447 3044 5596
rect 3108 5447 3109 5596
rect 3088 5447 3089 5598
rect 3098 5447 3099 5598
rect 2563 5604 2564 5607
rect 2578 5604 2579 5607
rect 2581 5606 2582 5707
rect 2653 5604 2654 5607
rect 2599 5604 2600 5609
rect 2702 5604 2703 5609
rect 2602 5604 2603 5611
rect 2768 5604 2769 5611
rect 2606 5604 2607 5613
rect 2684 5612 2685 5707
rect 2612 5604 2613 5615
rect 2759 5604 2760 5615
rect 2566 5604 2567 5617
rect 2760 5616 2761 5707
rect 2615 5604 2616 5619
rect 2756 5604 2757 5619
rect 2619 5604 2620 5621
rect 2714 5604 2715 5621
rect 2619 5622 2620 5707
rect 2644 5604 2645 5623
rect 2626 5604 2627 5625
rect 2741 5604 2742 5625
rect 2629 5604 2630 5627
rect 2744 5604 2745 5627
rect 2642 5628 2643 5707
rect 2705 5604 2706 5629
rect 2645 5630 2646 5707
rect 2708 5604 2709 5631
rect 2650 5604 2651 5633
rect 2717 5632 2718 5707
rect 2662 5604 2663 5635
rect 2705 5634 2706 5707
rect 2665 5604 2666 5637
rect 2714 5636 2715 5707
rect 2675 5638 2676 5707
rect 2676 5604 2677 5639
rect 2678 5638 2679 5707
rect 2679 5604 2680 5639
rect 2681 5638 2682 5707
rect 2738 5604 2739 5639
rect 2687 5640 2688 5707
rect 2792 5604 2793 5641
rect 2690 5604 2691 5643
rect 2795 5604 2796 5643
rect 2693 5604 2694 5645
rect 2837 5604 2838 5645
rect 2693 5646 2694 5707
rect 2747 5604 2748 5647
rect 2696 5648 2697 5707
rect 2750 5604 2751 5649
rect 2711 5604 2712 5651
rect 2798 5604 2799 5651
rect 2711 5652 2712 5707
rect 2771 5604 2772 5653
rect 2739 5654 2740 5707
rect 2780 5604 2781 5655
rect 2745 5656 2746 5707
rect 2786 5604 2787 5657
rect 2751 5658 2752 5707
rect 2804 5604 2805 5659
rect 2763 5660 2764 5707
rect 2825 5604 2826 5661
rect 2769 5662 2770 5707
rect 2840 5604 2841 5663
rect 2772 5664 2773 5707
rect 2828 5604 2829 5665
rect 2775 5666 2776 5707
rect 2852 5604 2853 5667
rect 2782 5668 2783 5707
rect 2882 5604 2883 5669
rect 2801 5604 2802 5671
rect 2822 5604 2823 5671
rect 2766 5672 2767 5707
rect 2800 5672 2801 5707
rect 2803 5672 2804 5707
rect 2849 5604 2850 5673
rect 2815 5674 2816 5707
rect 2846 5604 2847 5675
rect 2830 5676 2831 5707
rect 2888 5604 2889 5677
rect 2834 5604 2835 5679
rect 2916 5604 2917 5679
rect 2812 5680 2813 5707
rect 2833 5680 2834 5707
rect 2836 5680 2837 5707
rect 2913 5604 2914 5681
rect 2840 5682 2841 5707
rect 2937 5604 2938 5683
rect 2843 5684 2844 5707
rect 2947 5604 2948 5685
rect 2864 5604 2865 5687
rect 2891 5604 2892 5687
rect 2865 5688 2866 5707
rect 2957 5604 2958 5689
rect 2868 5690 2869 5707
rect 2960 5604 2961 5691
rect 2877 5692 2878 5707
rect 2972 5604 2973 5693
rect 2880 5694 2881 5707
rect 2975 5604 2976 5695
rect 2885 5604 2886 5697
rect 2894 5604 2895 5697
rect 2753 5604 2754 5699
rect 2893 5698 2894 5707
rect 2754 5700 2755 5707
rect 2807 5604 2808 5701
rect 2806 5702 2807 5707
rect 2818 5702 2819 5707
rect 2910 5604 2911 5703
rect 2919 5604 2920 5703
rect 2969 5604 2970 5703
rect 3021 5604 3022 5703
rect 3001 5604 3002 5705
rect 3008 5604 3009 5705
rect 2575 5711 2576 5714
rect 2619 5711 2620 5714
rect 2599 5711 2600 5716
rect 2606 5711 2607 5716
rect 2602 5711 2603 5718
rect 2684 5711 2685 5718
rect 2613 5711 2614 5720
rect 2693 5711 2694 5720
rect 2635 5711 2636 5722
rect 2696 5711 2697 5722
rect 2642 5711 2643 5724
rect 2675 5711 2676 5724
rect 2652 5711 2653 5726
rect 2714 5711 2715 5726
rect 2581 5711 2582 5728
rect 2713 5727 2714 5778
rect 2656 5711 2657 5730
rect 2681 5711 2682 5730
rect 2648 5731 2649 5778
rect 2655 5731 2656 5778
rect 2658 5731 2659 5778
rect 2685 5731 2686 5778
rect 2661 5733 2662 5778
rect 2711 5711 2712 5734
rect 2664 5735 2665 5778
rect 2717 5711 2718 5736
rect 2666 5711 2667 5738
rect 2705 5711 2706 5738
rect 2678 5711 2679 5740
rect 2694 5739 2695 5778
rect 2641 5741 2642 5778
rect 2679 5741 2680 5778
rect 2682 5741 2683 5778
rect 2697 5741 2698 5778
rect 2690 5711 2691 5744
rect 2754 5711 2755 5744
rect 2687 5711 2688 5746
rect 2691 5745 2692 5778
rect 2707 5745 2708 5778
rect 2739 5711 2740 5746
rect 2719 5747 2720 5778
rect 2734 5747 2735 5778
rect 2723 5711 2724 5750
rect 2745 5711 2746 5750
rect 2728 5751 2729 5778
rect 2772 5711 2773 5752
rect 2730 5711 2731 5754
rect 2751 5711 2752 5754
rect 2731 5755 2732 5778
rect 2775 5711 2776 5756
rect 2737 5757 2738 5778
rect 2755 5757 2756 5778
rect 2740 5759 2741 5778
rect 2800 5711 2801 5760
rect 2746 5761 2747 5778
rect 2815 5711 2816 5762
rect 2761 5763 2762 5778
rect 2806 5711 2807 5764
rect 2763 5711 2764 5766
rect 2769 5711 2770 5766
rect 2764 5767 2765 5778
rect 2847 5711 2848 5768
rect 2773 5769 2774 5778
rect 2830 5711 2831 5770
rect 2779 5771 2780 5778
rect 2812 5711 2813 5772
rect 2789 5773 2790 5778
rect 2877 5711 2878 5774
rect 2803 5711 2804 5776
rect 2833 5711 2834 5776
rect 2836 5711 2837 5776
rect 2843 5711 2844 5776
rect 2862 5711 2863 5776
rect 2865 5711 2866 5776
rect 2868 5711 2869 5776
rect 2874 5711 2875 5776
rect 2880 5711 2881 5776
rect 2883 5711 2884 5776
rect 2617 5782 2618 5785
rect 2761 5782 2762 5785
rect 2644 5782 2645 5787
rect 2664 5782 2665 5787
rect 2648 5782 2649 5789
rect 2789 5782 2790 5789
rect 2651 5782 2652 5791
rect 2661 5782 2662 5791
rect 2655 5782 2656 5793
rect 2656 5792 2657 5811
rect 2665 5792 2666 5811
rect 2685 5782 2686 5793
rect 2667 5782 2668 5795
rect 2668 5794 2669 5811
rect 2674 5794 2675 5811
rect 2691 5782 2692 5795
rect 2677 5796 2678 5811
rect 2697 5782 2698 5797
rect 2694 5782 2695 5799
rect 2703 5782 2704 5799
rect 2707 5798 2708 5811
rect 2728 5782 2729 5799
rect 2710 5800 2711 5811
rect 2731 5782 2732 5801
rect 2713 5782 2714 5803
rect 2719 5782 2720 5803
rect 2737 5802 2738 5811
rect 2773 5782 2774 5803
rect 2740 5782 2741 5805
rect 2767 5782 2768 5805
rect 2746 5782 2747 5807
rect 2786 5782 2787 5807
rect 2764 5782 2765 5809
rect 2770 5782 2771 5809
rect 2623 5815 2624 5818
rect 2737 5815 2738 5818
rect 2653 5815 2654 5820
rect 2677 5815 2678 5820
rect 2656 5815 2657 5822
rect 2668 5815 2669 5822
rect 2665 5815 2666 5824
rect 2674 5815 2675 5824
rect 2707 5815 2708 5824
rect 2716 5815 2717 5824
rect 2710 5815 2711 5826
rect 2713 5815 2714 5826
<< via >>
rect 2641 1271 2642 1272
rect 2737 1271 2738 1272
rect 2644 1273 2645 1274
rect 2647 1273 2648 1274
rect 2671 1273 2672 1274
rect 2684 1273 2685 1274
rect 2678 1275 2679 1276
rect 2687 1275 2688 1276
rect 2690 1275 2691 1276
rect 2693 1275 2694 1276
rect 2699 1275 2700 1276
rect 2708 1275 2709 1276
rect 2702 1277 2703 1278
rect 2705 1277 2706 1278
rect 2527 1287 2528 1288
rect 2533 1287 2534 1288
rect 2605 1287 2606 1288
rect 2839 1287 2840 1288
rect 2626 1289 2627 1290
rect 2645 1289 2646 1290
rect 2633 1291 2634 1292
rect 2662 1291 2663 1292
rect 2641 1293 2642 1294
rect 2677 1293 2678 1294
rect 2642 1295 2643 1296
rect 2655 1295 2656 1296
rect 2647 1297 2648 1298
rect 2674 1297 2675 1298
rect 2684 1297 2685 1298
rect 2714 1297 2715 1298
rect 2687 1299 2688 1300
rect 2721 1299 2722 1300
rect 2680 1301 2681 1302
rect 2686 1301 2687 1302
rect 2690 1301 2691 1302
rect 2727 1301 2728 1302
rect 2692 1303 2693 1304
rect 2730 1303 2731 1304
rect 2696 1305 2697 1306
rect 2711 1305 2712 1306
rect 2699 1307 2700 1308
rect 2751 1307 2752 1308
rect 2699 1309 2700 1310
rect 2708 1309 2709 1310
rect 2702 1311 2703 1312
rect 2748 1311 2749 1312
rect 2737 1313 2738 1314
rect 2827 1313 2828 1314
rect 2754 1315 2755 1316
rect 2815 1315 2816 1316
rect 2757 1317 2758 1318
rect 2851 1317 2852 1318
rect 2760 1319 2761 1320
rect 2775 1319 2776 1320
rect 2769 1321 2770 1322
rect 2794 1321 2795 1322
rect 2772 1323 2773 1324
rect 2791 1323 2792 1324
rect 2781 1325 2782 1326
rect 2845 1325 2846 1326
rect 2784 1327 2785 1328
rect 2824 1327 2825 1328
rect 2798 1329 2799 1330
rect 2830 1329 2831 1330
rect 2521 1338 2522 1339
rect 2539 1338 2540 1339
rect 2533 1340 2534 1341
rect 2545 1340 2546 1341
rect 2533 1342 2534 1343
rect 2542 1342 2543 1343
rect 2587 1342 2588 1343
rect 2596 1342 2597 1343
rect 2593 1344 2594 1345
rect 2648 1344 2649 1345
rect 2626 1346 2627 1347
rect 2689 1346 2690 1347
rect 2630 1348 2631 1349
rect 2642 1348 2643 1349
rect 2633 1350 2634 1351
rect 2645 1350 2646 1351
rect 2617 1352 2618 1353
rect 2646 1352 2647 1353
rect 2665 1352 2666 1353
rect 2711 1352 2712 1353
rect 2668 1354 2669 1355
rect 2674 1354 2675 1355
rect 2623 1356 2624 1357
rect 2674 1356 2675 1357
rect 2671 1358 2672 1359
rect 2677 1358 2678 1359
rect 2680 1358 2681 1359
rect 2686 1358 2687 1359
rect 2704 1358 2705 1359
rect 2708 1358 2709 1359
rect 2723 1358 2724 1359
rect 2798 1358 2799 1359
rect 2741 1360 2742 1361
rect 2751 1360 2752 1361
rect 2744 1362 2745 1363
rect 2754 1362 2755 1363
rect 2750 1364 2751 1365
rect 2757 1364 2758 1365
rect 2753 1366 2754 1367
rect 2760 1366 2761 1367
rect 2756 1368 2757 1369
rect 2772 1368 2773 1369
rect 2769 1370 2770 1371
rect 2771 1370 2772 1371
rect 2768 1372 2769 1373
rect 2794 1372 2795 1373
rect 2781 1374 2782 1375
rect 2866 1374 2867 1375
rect 2792 1376 2793 1377
rect 2805 1376 2806 1377
rect 2808 1376 2809 1377
rect 2863 1376 2864 1377
rect 2815 1378 2816 1379
rect 2836 1378 2837 1379
rect 2827 1380 2828 1381
rect 2833 1380 2834 1381
rect 2827 1382 2828 1383
rect 2839 1382 2840 1383
rect 2875 1382 2876 1383
rect 2895 1382 2896 1383
rect 2539 1391 2540 1392
rect 2620 1391 2621 1392
rect 2542 1393 2543 1394
rect 2561 1393 2562 1394
rect 2533 1395 2534 1396
rect 2543 1395 2544 1396
rect 2549 1395 2550 1396
rect 2558 1395 2559 1396
rect 2564 1395 2565 1396
rect 2861 1395 2862 1396
rect 2593 1397 2594 1398
rect 2611 1397 2612 1398
rect 2608 1399 2609 1400
rect 2661 1399 2662 1400
rect 2614 1401 2615 1402
rect 2721 1401 2722 1402
rect 2617 1403 2618 1404
rect 2682 1403 2683 1404
rect 2623 1405 2624 1406
rect 2643 1405 2644 1406
rect 2623 1407 2624 1408
rect 2715 1407 2716 1408
rect 2626 1409 2627 1410
rect 2709 1409 2710 1410
rect 2629 1411 2630 1412
rect 2706 1411 2707 1412
rect 2630 1413 2631 1414
rect 2739 1413 2740 1414
rect 2633 1415 2634 1416
rect 2697 1415 2698 1416
rect 2637 1417 2638 1418
rect 2736 1417 2737 1418
rect 2652 1419 2653 1420
rect 2664 1419 2665 1420
rect 2668 1419 2669 1420
rect 2703 1419 2704 1420
rect 2671 1421 2672 1422
rect 2685 1421 2686 1422
rect 2700 1421 2701 1422
rect 2766 1421 2767 1422
rect 2711 1423 2712 1424
rect 2782 1423 2783 1424
rect 2646 1425 2647 1426
rect 2712 1425 2713 1426
rect 2545 1427 2546 1428
rect 2646 1427 2647 1428
rect 2723 1427 2724 1428
rect 2800 1427 2801 1428
rect 2726 1429 2727 1430
rect 2803 1429 2804 1430
rect 2741 1431 2742 1432
rect 2857 1431 2858 1432
rect 2747 1433 2748 1434
rect 2868 1433 2869 1434
rect 2750 1435 2751 1436
rect 2806 1435 2807 1436
rect 2753 1437 2754 1438
rect 2809 1437 2810 1438
rect 2754 1439 2755 1440
rect 2760 1439 2761 1440
rect 2756 1441 2757 1442
rect 2839 1441 2840 1442
rect 2757 1443 2758 1444
rect 2836 1443 2837 1444
rect 2763 1445 2764 1446
rect 2768 1445 2769 1446
rect 2769 1447 2770 1448
rect 2909 1447 2910 1448
rect 2771 1449 2772 1450
rect 2818 1449 2819 1450
rect 2680 1451 2681 1452
rect 2772 1451 2773 1452
rect 2679 1453 2680 1454
rect 2877 1453 2878 1454
rect 2778 1455 2779 1456
rect 2821 1455 2822 1456
rect 2792 1457 2793 1458
rect 2848 1457 2849 1458
rect 2824 1459 2825 1460
rect 2916 1459 2917 1460
rect 2744 1461 2745 1462
rect 2824 1461 2825 1462
rect 2827 1461 2828 1462
rect 2904 1461 2905 1462
rect 2830 1463 2831 1464
rect 2886 1463 2887 1464
rect 2833 1465 2834 1466
rect 2889 1465 2890 1466
rect 2798 1467 2799 1468
rect 2833 1467 2834 1468
rect 2851 1467 2852 1468
rect 2907 1467 2908 1468
rect 2863 1469 2864 1470
rect 2939 1469 2940 1470
rect 2866 1471 2867 1472
rect 2945 1471 2946 1472
rect 2875 1473 2876 1474
rect 2956 1473 2957 1474
rect 2815 1475 2816 1476
rect 2874 1475 2875 1476
rect 2910 1475 2911 1476
rect 2913 1475 2914 1476
rect 2551 1484 2552 1485
rect 2558 1484 2559 1485
rect 2611 1484 2612 1485
rect 2636 1484 2637 1485
rect 2617 1486 2618 1487
rect 2780 1486 2781 1487
rect 2620 1488 2621 1489
rect 2659 1488 2660 1489
rect 2623 1490 2624 1491
rect 2712 1490 2713 1491
rect 2626 1492 2627 1493
rect 2677 1492 2678 1493
rect 2630 1494 2631 1495
rect 2715 1494 2716 1495
rect 2649 1496 2650 1497
rect 2706 1496 2707 1497
rect 2661 1498 2662 1499
rect 2783 1498 2784 1499
rect 2643 1500 2644 1501
rect 2662 1500 2663 1501
rect 2674 1500 2675 1501
rect 2762 1500 2763 1501
rect 2679 1502 2680 1503
rect 2968 1502 2969 1503
rect 2685 1504 2686 1505
rect 2711 1504 2712 1505
rect 2689 1506 2690 1507
rect 2965 1506 2966 1507
rect 2693 1508 2694 1509
rect 2754 1508 2755 1509
rect 2697 1510 2698 1511
rect 2729 1510 2730 1511
rect 2696 1512 2697 1513
rect 2798 1512 2799 1513
rect 2703 1514 2704 1515
rect 2717 1514 2718 1515
rect 2709 1516 2710 1517
rect 2747 1516 2748 1517
rect 2739 1518 2740 1519
rect 2789 1518 2790 1519
rect 2800 1518 2801 1519
rect 2846 1518 2847 1519
rect 2671 1520 2672 1521
rect 2801 1520 2802 1521
rect 2803 1520 2804 1521
rect 2840 1520 2841 1521
rect 2806 1522 2807 1523
rect 2831 1522 2832 1523
rect 2818 1524 2819 1525
rect 2864 1524 2865 1525
rect 2809 1526 2810 1527
rect 2819 1526 2820 1527
rect 2766 1528 2767 1529
rect 2810 1528 2811 1529
rect 2682 1530 2683 1531
rect 2765 1530 2766 1531
rect 2824 1530 2825 1531
rect 2858 1530 2859 1531
rect 2772 1532 2773 1533
rect 2825 1532 2826 1533
rect 2848 1532 2849 1533
rect 2900 1532 2901 1533
rect 2785 1534 2786 1535
rect 2849 1534 2850 1535
rect 2736 1536 2737 1537
rect 2786 1536 2787 1537
rect 2735 1538 2736 1539
rect 2778 1538 2779 1539
rect 2868 1538 2869 1539
rect 2892 1538 2893 1539
rect 2646 1540 2647 1541
rect 2891 1540 2892 1541
rect 2646 1542 2647 1543
rect 2652 1542 2653 1543
rect 2874 1542 2875 1543
rect 2987 1542 2988 1543
rect 2833 1544 2834 1545
rect 2873 1544 2874 1545
rect 2775 1546 2776 1547
rect 2834 1546 2835 1547
rect 2757 1548 2758 1549
rect 2774 1548 2775 1549
rect 2686 1550 2687 1551
rect 2756 1550 2757 1551
rect 2877 1550 2878 1551
rect 2897 1550 2898 1551
rect 2721 1552 2722 1553
rect 2876 1552 2877 1553
rect 2664 1554 2665 1555
rect 2720 1554 2721 1555
rect 2886 1554 2887 1555
rect 2953 1554 2954 1555
rect 2821 1556 2822 1557
rect 2885 1556 2886 1557
rect 2769 1558 2770 1559
rect 2822 1558 2823 1559
rect 2904 1558 2905 1559
rect 2944 1558 2945 1559
rect 2851 1560 2852 1561
rect 2903 1560 2904 1561
rect 2913 1560 2914 1561
rect 2959 1560 2960 1561
rect 2916 1562 2917 1563
rect 2962 1562 2963 1563
rect 2939 1564 2940 1565
rect 3004 1564 3005 1565
rect 2956 1566 2957 1567
rect 3007 1566 3008 1567
rect 2889 1568 2890 1569
rect 2956 1568 2957 1569
rect 2760 1570 2761 1571
rect 2888 1570 2889 1571
rect 2971 1570 2972 1571
rect 2980 1570 2981 1571
rect 2974 1572 2975 1573
rect 2977 1572 2978 1573
rect 2560 1581 2561 1582
rect 2651 1581 2652 1582
rect 2563 1583 2564 1584
rect 2654 1583 2655 1584
rect 2605 1585 2606 1586
rect 3104 1585 3105 1586
rect 2656 1587 2657 1588
rect 2762 1587 2763 1588
rect 2659 1589 2660 1590
rect 2713 1589 2714 1590
rect 2662 1591 2663 1592
rect 2685 1591 2686 1592
rect 2667 1593 2668 1594
rect 2765 1593 2766 1594
rect 2693 1595 2694 1596
rect 2791 1595 2792 1596
rect 2711 1597 2712 1598
rect 2758 1597 2759 1598
rect 2717 1599 2718 1600
rect 2764 1599 2765 1600
rect 2677 1601 2678 1602
rect 2716 1601 2717 1602
rect 2636 1603 2637 1604
rect 2676 1603 2677 1604
rect 2720 1603 2721 1604
rect 2794 1603 2795 1604
rect 2722 1605 2723 1606
rect 2864 1605 2865 1606
rect 2729 1607 2730 1608
rect 2806 1607 2807 1608
rect 2747 1609 2748 1610
rect 2803 1609 2804 1610
rect 2746 1611 2747 1612
rect 2756 1611 2757 1612
rect 2768 1611 2769 1612
rect 2861 1611 2862 1612
rect 2780 1613 2781 1614
rect 2828 1613 2829 1614
rect 2631 1615 2632 1616
rect 2779 1615 2780 1616
rect 2783 1615 2784 1616
rect 2831 1615 2832 1616
rect 2626 1617 2627 1618
rect 2782 1617 2783 1618
rect 2798 1617 2799 1618
rect 2855 1617 2856 1618
rect 2789 1619 2790 1620
rect 2797 1619 2798 1620
rect 2810 1619 2811 1620
rect 2812 1619 2813 1620
rect 2837 1619 2838 1620
rect 2867 1619 2868 1620
rect 2638 1621 2639 1622
rect 2837 1621 2838 1622
rect 2846 1621 2847 1622
rect 2891 1621 2892 1622
rect 2708 1623 2709 1624
rect 2846 1623 2847 1624
rect 2623 1625 2624 1626
rect 2707 1625 2708 1626
rect 2849 1625 2850 1626
rect 2894 1625 2895 1626
rect 2774 1627 2775 1628
rect 2849 1627 2850 1628
rect 2634 1629 2635 1630
rect 2773 1629 2774 1630
rect 2873 1629 2874 1630
rect 2913 1629 2914 1630
rect 2819 1631 2820 1632
rect 2912 1631 2913 1632
rect 2819 1633 2820 1634
rect 2840 1633 2841 1634
rect 2822 1635 2823 1636
rect 2873 1635 2874 1636
rect 2876 1635 2877 1636
rect 2948 1635 2949 1636
rect 2825 1637 2826 1638
rect 2876 1637 2877 1638
rect 2649 1639 2650 1640
rect 2825 1639 2826 1640
rect 2885 1639 2886 1640
rect 2927 1639 2928 1640
rect 2834 1641 2835 1642
rect 2885 1641 2886 1642
rect 2786 1643 2787 1644
rect 2834 1643 2835 1644
rect 2888 1643 2889 1644
rect 2930 1643 2931 1644
rect 2771 1645 2772 1646
rect 2888 1645 2889 1646
rect 2735 1647 2736 1648
rect 2770 1647 2771 1648
rect 2612 1649 2613 1650
rect 2734 1649 2735 1650
rect 2897 1649 2898 1650
rect 2951 1649 2952 1650
rect 2916 1651 2917 1652
rect 2980 1651 2981 1652
rect 2858 1653 2859 1654
rect 2915 1653 2916 1654
rect 2801 1655 2802 1656
rect 2858 1655 2859 1656
rect 2953 1655 2954 1656
rect 3020 1655 3021 1656
rect 2909 1657 2910 1658
rect 2954 1657 2955 1658
rect 2956 1657 2957 1658
rect 3023 1657 3024 1658
rect 2959 1659 2960 1660
rect 3014 1659 3015 1660
rect 2900 1661 2901 1662
rect 2960 1661 2961 1662
rect 2962 1661 2963 1662
rect 3002 1661 3003 1662
rect 2903 1663 2904 1664
rect 2963 1663 2964 1664
rect 2965 1663 2966 1664
rect 3026 1663 3027 1664
rect 2968 1665 2969 1666
rect 3029 1665 3030 1666
rect 2971 1667 2972 1668
rect 2998 1667 2999 1668
rect 2944 1669 2945 1670
rect 2999 1669 3000 1670
rect 2921 1671 2922 1672
rect 2945 1671 2946 1672
rect 2974 1671 2975 1672
rect 2984 1671 2985 1672
rect 3004 1671 3005 1672
rect 3063 1671 3064 1672
rect 3007 1673 3008 1674
rect 3066 1673 3067 1674
rect 3044 1675 3045 1676
rect 3055 1675 3056 1676
rect 3047 1677 3048 1678
rect 3052 1677 3053 1678
rect 2533 1686 2534 1687
rect 2654 1686 2655 1687
rect 2551 1688 2552 1689
rect 2593 1688 2594 1689
rect 2575 1690 2576 1691
rect 2663 1690 2664 1691
rect 2590 1692 2591 1693
rect 2625 1692 2626 1693
rect 2605 1694 2606 1695
rect 2734 1694 2735 1695
rect 2605 1696 2606 1697
rect 2904 1696 2905 1697
rect 2619 1698 2620 1699
rect 2773 1698 2774 1699
rect 2619 1700 2620 1701
rect 2803 1700 2804 1701
rect 2612 1702 2613 1703
rect 2802 1702 2803 1703
rect 2628 1704 2629 1705
rect 2667 1704 2668 1705
rect 2634 1706 2635 1707
rect 2679 1706 2680 1707
rect 2643 1708 2644 1709
rect 2764 1708 2765 1709
rect 2660 1710 2661 1711
rect 2676 1710 2677 1711
rect 2696 1710 2697 1711
rect 2713 1710 2714 1711
rect 2699 1712 2700 1713
rect 2707 1712 2708 1713
rect 2705 1714 2706 1715
rect 2716 1714 2717 1715
rect 2730 1714 2731 1715
rect 3018 1714 3019 1715
rect 2748 1716 2749 1717
rect 2758 1716 2759 1717
rect 2766 1716 2767 1717
rect 2779 1716 2780 1717
rect 2772 1718 2773 1719
rect 2837 1718 2838 1719
rect 2770 1720 2771 1721
rect 2838 1720 2839 1721
rect 2769 1722 2770 1723
rect 2782 1722 2783 1723
rect 2778 1724 2779 1725
rect 2791 1724 2792 1725
rect 2781 1726 2782 1727
rect 2794 1726 2795 1727
rect 2784 1728 2785 1729
rect 2797 1728 2798 1729
rect 2746 1730 2747 1731
rect 2796 1730 2797 1731
rect 2790 1732 2791 1733
rect 2806 1732 2807 1733
rect 2685 1734 2686 1735
rect 2805 1734 2806 1735
rect 2684 1736 2685 1737
rect 2888 1736 2889 1737
rect 2808 1738 2809 1739
rect 2828 1738 2829 1739
rect 2669 1740 2670 1741
rect 2829 1740 2830 1741
rect 2812 1742 2813 1743
rect 2919 1742 2920 1743
rect 2811 1744 2812 1745
rect 2831 1744 2832 1745
rect 2820 1746 2821 1747
rect 2825 1746 2826 1747
rect 2638 1748 2639 1749
rect 2826 1748 2827 1749
rect 2637 1750 2638 1751
rect 2651 1750 2652 1751
rect 2622 1752 2623 1753
rect 2650 1752 2651 1753
rect 2823 1752 2824 1753
rect 2834 1752 2835 1753
rect 2631 1754 2632 1755
rect 2835 1754 2836 1755
rect 2853 1754 2854 1755
rect 2873 1754 2874 1755
rect 2855 1756 2856 1757
rect 2865 1756 2866 1757
rect 2856 1758 2857 1759
rect 2876 1758 2877 1759
rect 2861 1760 2862 1761
rect 2901 1760 2902 1761
rect 2867 1762 2868 1763
rect 2877 1762 2878 1763
rect 2858 1764 2859 1765
rect 2868 1764 2869 1765
rect 2849 1766 2850 1767
rect 2859 1766 2860 1767
rect 2733 1768 2734 1769
rect 2850 1768 2851 1769
rect 2883 1768 2884 1769
rect 2885 1768 2886 1769
rect 2894 1768 2895 1769
rect 2925 1768 2926 1769
rect 2907 1770 2908 1771
rect 2930 1770 2931 1771
rect 2909 1772 2910 1773
rect 2967 1772 2968 1773
rect 2921 1774 2922 1775
rect 3012 1774 3013 1775
rect 2931 1776 2932 1777
rect 2948 1776 2949 1777
rect 2726 1778 2727 1779
rect 2949 1778 2950 1779
rect 2937 1780 2938 1781
rect 2945 1780 2946 1781
rect 2951 1780 2952 1781
rect 3089 1780 3090 1781
rect 2952 1782 2953 1783
rect 2969 1782 2970 1783
rect 2955 1784 2956 1785
rect 2976 1784 2977 1785
rect 2958 1786 2959 1787
rect 2960 1786 2961 1787
rect 2961 1788 2962 1789
rect 2963 1788 2964 1789
rect 2973 1788 2974 1789
rect 3113 1788 3114 1789
rect 2976 1790 2977 1791
rect 3002 1790 3003 1791
rect 2983 1792 2984 1793
rect 2990 1792 2991 1793
rect 2994 1792 2995 1793
rect 3014 1792 3015 1793
rect 2927 1794 2928 1795
rect 3015 1794 3016 1795
rect 2891 1796 2892 1797
rect 2928 1796 2929 1797
rect 3003 1796 3004 1797
rect 3097 1796 3098 1797
rect 3006 1798 3007 1799
rect 3151 1798 3152 1799
rect 3020 1800 3021 1801
rect 3055 1800 3056 1801
rect 3021 1802 3022 1803
rect 3026 1802 3027 1803
rect 2915 1804 2916 1805
rect 3027 1804 3028 1805
rect 3023 1806 3024 1807
rect 3058 1806 3059 1807
rect 3029 1808 3030 1809
rect 3074 1808 3075 1809
rect 3063 1810 3064 1811
rect 3112 1810 3113 1811
rect 2964 1812 2965 1813
rect 3064 1812 3065 1813
rect 3066 1812 3067 1813
rect 3072 1812 3073 1813
rect 2912 1814 2913 1815
rect 3071 1814 3072 1815
rect 3083 1814 3084 1815
rect 3119 1814 3120 1815
rect 3106 1816 3107 1817
rect 3109 1816 3110 1817
rect 2548 1825 2549 1826
rect 2578 1825 2579 1826
rect 2552 1827 2553 1828
rect 2575 1827 2576 1828
rect 2587 1827 2588 1828
rect 2663 1827 2664 1828
rect 2593 1829 2594 1830
rect 2599 1829 2600 1830
rect 2593 1831 2594 1832
rect 2714 1831 2715 1832
rect 2605 1833 2606 1834
rect 2817 1833 2818 1834
rect 2619 1835 2620 1836
rect 2705 1835 2706 1836
rect 2622 1837 2623 1838
rect 2625 1837 2626 1838
rect 2637 1837 2638 1838
rect 2652 1837 2653 1838
rect 2634 1839 2635 1840
rect 2636 1839 2637 1840
rect 2640 1839 2641 1840
rect 2823 1839 2824 1840
rect 2647 1841 2648 1842
rect 2865 1841 2866 1842
rect 2657 1843 2658 1844
rect 2778 1843 2779 1844
rect 2664 1845 2665 1846
rect 2676 1845 2677 1846
rect 2667 1847 2668 1848
rect 2850 1847 2851 1848
rect 2683 1849 2684 1850
rect 2796 1849 2797 1850
rect 2687 1851 2688 1852
rect 2772 1851 2773 1852
rect 2615 1853 2616 1854
rect 2772 1853 2773 1854
rect 2690 1855 2691 1856
rect 2781 1855 2782 1856
rect 2696 1857 2697 1858
rect 2717 1857 2718 1858
rect 2699 1859 2700 1860
rect 2702 1859 2703 1860
rect 2723 1859 2724 1860
rect 2823 1859 2824 1860
rect 2730 1861 2731 1862
rect 2847 1861 2848 1862
rect 2733 1863 2734 1864
rect 2892 1863 2893 1864
rect 2748 1865 2749 1866
rect 2751 1865 2752 1866
rect 2766 1865 2767 1866
rect 2778 1865 2779 1866
rect 2655 1867 2656 1868
rect 2766 1867 2767 1868
rect 2769 1867 2770 1868
rect 2781 1867 2782 1868
rect 2784 1867 2785 1868
rect 2793 1867 2794 1868
rect 2790 1869 2791 1870
rect 2799 1869 2800 1870
rect 2790 1871 2791 1872
rect 2820 1871 2821 1872
rect 2805 1873 2806 1874
rect 2832 1873 2833 1874
rect 2829 1875 2830 1876
rect 2841 1875 2842 1876
rect 2802 1877 2803 1878
rect 2829 1877 2830 1878
rect 2838 1877 2839 1878
rect 2862 1877 2863 1878
rect 2811 1879 2812 1880
rect 2838 1879 2839 1880
rect 2726 1881 2727 1882
rect 2811 1881 2812 1882
rect 2847 1881 2848 1882
rect 3140 1881 3141 1882
rect 2856 1883 2857 1884
rect 2886 1883 2887 1884
rect 2826 1885 2827 1886
rect 2856 1885 2857 1886
rect 2859 1885 2860 1886
rect 2871 1885 2872 1886
rect 2835 1887 2836 1888
rect 2859 1887 2860 1888
rect 2808 1889 2809 1890
rect 2835 1889 2836 1890
rect 2868 1889 2869 1890
rect 2874 1889 2875 1890
rect 2877 1889 2878 1890
rect 2895 1889 2896 1890
rect 2877 1891 2878 1892
rect 2904 1891 2905 1892
rect 2889 1893 2890 1894
rect 2967 1893 2968 1894
rect 2901 1895 2902 1896
rect 2910 1895 2911 1896
rect 2904 1897 2905 1898
rect 2907 1897 2908 1898
rect 2883 1899 2884 1900
rect 2907 1899 2908 1900
rect 2853 1901 2854 1902
rect 2883 1901 2884 1902
rect 2643 1903 2644 1904
rect 2853 1903 2854 1904
rect 2913 1903 2914 1904
rect 2928 1903 2929 1904
rect 2916 1905 2917 1906
rect 2925 1905 2926 1906
rect 2919 1907 2920 1908
rect 2922 1907 2923 1908
rect 2919 1909 2920 1910
rect 2949 1909 2950 1910
rect 2931 1911 2932 1912
rect 2934 1911 2935 1912
rect 2937 1911 2938 1912
rect 2985 1911 2986 1912
rect 2940 1913 2941 1914
rect 2961 1913 2962 1914
rect 2949 1915 2950 1916
rect 3015 1915 3016 1916
rect 2958 1917 2959 1918
rect 2970 1917 2971 1918
rect 2955 1919 2956 1920
rect 2958 1919 2959 1920
rect 2952 1921 2953 1922
rect 2955 1921 2956 1922
rect 2952 1923 2953 1924
rect 3018 1923 3019 1924
rect 2964 1925 2965 1926
rect 2982 1925 2983 1926
rect 2967 1927 2968 1928
rect 3100 1927 3101 1928
rect 2979 1929 2980 1930
rect 3071 1929 3072 1930
rect 2991 1931 2992 1932
rect 3012 1931 3013 1932
rect 2994 1933 2995 1934
rect 3018 1933 3019 1934
rect 2994 1935 2995 1936
rect 3003 1935 3004 1936
rect 3000 1937 3001 1938
rect 3135 1937 3136 1938
rect 2973 1939 2974 1940
rect 3000 1939 3001 1940
rect 3006 1939 3007 1940
rect 3024 1939 3025 1940
rect 2976 1941 2977 1942
rect 3006 1941 3007 1942
rect 3021 1941 3022 1942
rect 3036 1941 3037 1942
rect 3034 1943 3035 1944
rect 3064 1943 3065 1944
rect 3043 1945 3044 1946
rect 3129 1945 3130 1946
rect 3046 1947 3047 1948
rect 3048 1947 3049 1948
rect 3045 1949 3046 1950
rect 3083 1949 3084 1950
rect 3055 1951 3056 1952
rect 3066 1951 3067 1952
rect 3058 1953 3059 1954
rect 3069 1953 3070 1954
rect 3074 1953 3075 1954
rect 3093 1953 3094 1954
rect 3092 1955 3093 1956
rect 3106 1955 3107 1956
rect 3114 1955 3115 1956
rect 3154 1955 3155 1956
rect 3117 1957 3118 1958
rect 3154 1957 3155 1958
rect 3126 1959 3127 1960
rect 3164 1959 3165 1960
rect 3132 1961 3133 1962
rect 3150 1961 3151 1962
rect 3144 1963 3145 1964
rect 3147 1963 3148 1964
rect 3144 1965 3145 1966
rect 3170 1965 3171 1966
rect 2596 1974 2597 1975
rect 2707 1974 2708 1975
rect 2609 1976 2610 1977
rect 2702 1976 2703 1977
rect 2587 1978 2588 1979
rect 2609 1978 2610 1979
rect 2615 1978 2616 1979
rect 2619 1978 2620 1979
rect 2619 1980 2620 1981
rect 2692 1980 2693 1981
rect 2623 1982 2624 1983
rect 2856 1982 2857 1983
rect 2626 1984 2627 1985
rect 2719 1984 2720 1985
rect 2629 1986 2630 1987
rect 2814 1986 2815 1987
rect 2633 1988 2634 1989
rect 2646 1988 2647 1989
rect 2636 1990 2637 1991
rect 2680 1990 2681 1991
rect 2649 1992 2650 1993
rect 2766 1992 2767 1993
rect 2656 1994 2657 1995
rect 2859 1994 2860 1995
rect 2658 1996 2659 1997
rect 2664 1996 2665 1997
rect 2661 1998 2662 1999
rect 2704 1998 2705 1999
rect 2683 2000 2684 2001
rect 2874 2000 2875 2001
rect 2652 2002 2653 2003
rect 2683 2002 2684 2003
rect 2642 2004 2643 2005
rect 2653 2004 2654 2005
rect 2690 2004 2691 2005
rect 2769 2004 2770 2005
rect 2695 2006 2696 2007
rect 3141 2006 3142 2007
rect 2714 2008 2715 2009
rect 2745 2008 2746 2009
rect 2717 2010 2718 2011
rect 2748 2010 2749 2011
rect 2725 2012 2726 2013
rect 2790 2012 2791 2013
rect 2732 2014 2733 2015
rect 2892 2014 2893 2015
rect 2633 2016 2634 2017
rect 2892 2016 2893 2017
rect 2772 2018 2773 2019
rect 2904 2018 2905 2019
rect 2802 2020 2803 2021
rect 2865 2020 2866 2021
rect 2823 2022 2824 2023
rect 2859 2022 2860 2023
rect 2829 2024 2830 2025
rect 2865 2024 2866 2025
rect 2647 2026 2648 2027
rect 2829 2026 2830 2027
rect 2832 2026 2833 2027
rect 2868 2026 2869 2027
rect 2742 2028 2743 2029
rect 2832 2028 2833 2029
rect 2838 2028 2839 2029
rect 2880 2028 2881 2029
rect 2886 2028 2887 2029
rect 2925 2028 2926 2029
rect 2862 2030 2863 2031
rect 2886 2030 2887 2031
rect 2901 2030 2902 2031
rect 3081 2030 3082 2031
rect 2871 2032 2872 2033
rect 2901 2032 2902 2033
rect 2847 2034 2848 2035
rect 2871 2034 2872 2035
rect 2811 2036 2812 2037
rect 2847 2036 2848 2037
rect 2778 2038 2779 2039
rect 2811 2038 2812 2039
rect 2910 2038 2911 2039
rect 2943 2038 2944 2039
rect 2913 2040 2914 2041
rect 2946 2040 2947 2041
rect 2895 2042 2896 2043
rect 2913 2042 2914 2043
rect 2735 2044 2736 2045
rect 2895 2044 2896 2045
rect 2686 2046 2687 2047
rect 2735 2046 2736 2047
rect 2605 2048 2606 2049
rect 2686 2048 2687 2049
rect 2919 2048 2920 2049
rect 2928 2048 2929 2049
rect 2889 2050 2890 2051
rect 2919 2050 2920 2051
rect 2853 2052 2854 2053
rect 2889 2052 2890 2053
rect 2817 2054 2818 2055
rect 2853 2054 2854 2055
rect 2934 2054 2935 2055
rect 2976 2054 2977 2055
rect 2940 2056 2941 2057
rect 3015 2056 3016 2057
rect 2907 2058 2908 2059
rect 2940 2058 2941 2059
rect 2877 2060 2878 2061
rect 2907 2060 2908 2061
rect 2835 2062 2836 2063
rect 2877 2062 2878 2063
rect 2793 2064 2794 2065
rect 2835 2064 2836 2065
rect 2751 2066 2752 2067
rect 2793 2066 2794 2067
rect 2751 2068 2752 2069
rect 2781 2068 2782 2069
rect 2781 2070 2782 2071
rect 2964 2070 2965 2071
rect 2967 2070 2968 2071
rect 3003 2070 3004 2071
rect 2952 2072 2953 2073
rect 2967 2072 2968 2073
rect 2979 2072 2980 2073
rect 3102 2072 3103 2073
rect 2988 2074 2989 2075
rect 3039 2074 3040 2075
rect 2955 2076 2956 2077
rect 2988 2076 2989 2077
rect 2916 2078 2917 2079
rect 2955 2078 2956 2079
rect 3000 2078 3001 2079
rect 3191 2078 3192 2079
rect 3006 2080 3007 2081
rect 3039 2080 3040 2081
rect 3012 2082 3013 2083
rect 3084 2082 3085 2083
rect 3015 2084 3016 2085
rect 3098 2084 3099 2085
rect 2982 2086 2983 2087
rect 3099 2086 3100 2087
rect 2949 2088 2950 2089
rect 2982 2088 2983 2089
rect 3018 2088 3019 2089
rect 3195 2088 3196 2089
rect 2991 2090 2992 2091
rect 3018 2090 3019 2091
rect 2958 2092 2959 2093
rect 2991 2092 2992 2093
rect 2922 2094 2923 2095
rect 2958 2094 2959 2095
rect 2883 2096 2884 2097
rect 2922 2096 2923 2097
rect 2841 2098 2842 2099
rect 2883 2098 2884 2099
rect 2799 2100 2800 2101
rect 2841 2100 2842 2101
rect 2799 2102 2800 2103
rect 2952 2102 2953 2103
rect 3027 2102 3028 2103
rect 3120 2102 3121 2103
rect 3033 2104 3034 2105
rect 3135 2104 3136 2105
rect 3036 2106 3037 2107
rect 3159 2106 3160 2107
rect 3045 2108 3046 2109
rect 3105 2108 3106 2109
rect 3024 2110 3025 2111
rect 3045 2110 3046 2111
rect 3048 2110 3049 2111
rect 3063 2110 3064 2111
rect 3075 2110 3076 2111
rect 3089 2110 3090 2111
rect 3092 2110 3093 2111
rect 3095 2110 3096 2111
rect 3066 2112 3067 2113
rect 3093 2112 3094 2113
rect 3069 2114 3070 2115
rect 3096 2114 3097 2115
rect 3114 2114 3115 2115
rect 3157 2114 3158 2115
rect 3117 2116 3118 2117
rect 3135 2116 3136 2117
rect 3122 2118 3123 2119
rect 3156 2118 3157 2119
rect 3129 2120 3130 2121
rect 3147 2120 3148 2121
rect 3132 2122 3133 2123
rect 3171 2122 3172 2123
rect 3144 2124 3145 2125
rect 3177 2124 3178 2125
rect 3126 2126 3127 2127
rect 3144 2126 3145 2127
rect 3150 2126 3151 2127
rect 3168 2126 3169 2127
rect 2994 2128 2995 2129
rect 3150 2128 3151 2129
rect 2994 2130 2995 2131
rect 3021 2130 3022 2131
rect 3174 2130 3175 2131
rect 3184 2130 3185 2131
rect 3204 2130 3205 2131
rect 3208 2130 3209 2131
rect 2594 2139 2595 2140
rect 2851 2139 2852 2140
rect 2587 2141 2588 2142
rect 2594 2141 2595 2142
rect 2603 2141 2604 2142
rect 2853 2141 2854 2142
rect 2604 2143 2605 2144
rect 2617 2143 2618 2144
rect 2619 2143 2620 2144
rect 2686 2143 2687 2144
rect 2620 2145 2621 2146
rect 2692 2145 2693 2146
rect 2622 2147 2623 2148
rect 2695 2147 2696 2148
rect 2626 2149 2627 2150
rect 2854 2149 2855 2150
rect 2633 2151 2634 2152
rect 2899 2151 2900 2152
rect 2633 2153 2634 2154
rect 2707 2153 2708 2154
rect 2637 2155 2638 2156
rect 2751 2155 2752 2156
rect 2640 2157 2641 2158
rect 2865 2157 2866 2158
rect 2643 2159 2644 2160
rect 2687 2159 2688 2160
rect 2644 2161 2645 2162
rect 2935 2161 2936 2162
rect 2650 2163 2651 2164
rect 2821 2163 2822 2164
rect 2650 2165 2651 2166
rect 2653 2165 2654 2166
rect 2653 2167 2654 2168
rect 2776 2167 2777 2168
rect 2660 2169 2661 2170
rect 2793 2169 2794 2170
rect 2666 2171 2667 2172
rect 2868 2171 2869 2172
rect 2669 2173 2670 2174
rect 2680 2173 2681 2174
rect 2672 2175 2673 2176
rect 2683 2175 2684 2176
rect 2681 2177 2682 2178
rect 2892 2177 2893 2178
rect 2693 2179 2694 2180
rect 2704 2179 2705 2180
rect 2702 2181 2703 2182
rect 2719 2181 2720 2182
rect 2733 2181 2734 2182
rect 2745 2181 2746 2182
rect 2742 2183 2743 2184
rect 2880 2183 2881 2184
rect 2748 2185 2749 2186
rect 2754 2185 2755 2186
rect 2748 2187 2749 2188
rect 2769 2187 2770 2188
rect 2794 2187 2795 2188
rect 2904 2187 2905 2188
rect 2735 2189 2736 2190
rect 2905 2189 2906 2190
rect 2809 2191 2810 2192
rect 2811 2191 2812 2192
rect 2814 2191 2815 2192
rect 2893 2191 2894 2192
rect 2827 2193 2828 2194
rect 2835 2193 2836 2194
rect 2829 2195 2830 2196
rect 2839 2195 2840 2196
rect 2845 2195 2846 2196
rect 2847 2195 2848 2196
rect 2866 2195 2867 2196
rect 2871 2195 2872 2196
rect 2872 2197 2873 2198
rect 2943 2197 2944 2198
rect 2881 2199 2882 2200
rect 2886 2199 2887 2200
rect 2597 2201 2598 2202
rect 2887 2201 2888 2202
rect 2895 2201 2896 2202
rect 2950 2201 2951 2202
rect 2889 2203 2890 2204
rect 2896 2203 2897 2204
rect 2606 2205 2607 2206
rect 2890 2205 2891 2206
rect 2600 2207 2601 2208
rect 2607 2207 2608 2208
rect 2601 2209 2602 2210
rect 2609 2209 2610 2210
rect 2610 2211 2611 2212
rect 2800 2211 2801 2212
rect 2925 2211 2926 2212
rect 2932 2211 2933 2212
rect 2919 2213 2920 2214
rect 2926 2213 2927 2214
rect 2715 2215 2716 2216
rect 2920 2215 2921 2216
rect 2928 2215 2929 2216
rect 2985 2215 2986 2216
rect 2922 2217 2923 2218
rect 2929 2217 2930 2218
rect 2955 2217 2956 2218
rect 2962 2217 2963 2218
rect 2964 2217 2965 2218
rect 2971 2217 2972 2218
rect 2958 2219 2959 2220
rect 2965 2219 2966 2220
rect 2952 2221 2953 2222
rect 2959 2221 2960 2222
rect 2946 2223 2947 2224
rect 2953 2223 2954 2224
rect 2940 2225 2941 2226
rect 2947 2225 2948 2226
rect 2967 2225 2968 2226
rect 2974 2225 2975 2226
rect 2976 2225 2977 2226
rect 3009 2225 3010 2226
rect 2991 2227 2992 2228
rect 2998 2227 2999 2228
rect 3000 2227 3001 2228
rect 3075 2227 3076 2228
rect 2994 2229 2995 2230
rect 3001 2229 3002 2230
rect 2988 2231 2989 2232
rect 2995 2231 2996 2232
rect 3015 2231 3016 2232
rect 3115 2231 3116 2232
rect 3018 2233 3019 2234
rect 3031 2233 3032 2234
rect 3027 2235 3028 2236
rect 3076 2235 3077 2236
rect 3033 2237 3034 2238
rect 3067 2237 3068 2238
rect 3037 2239 3038 2240
rect 3215 2239 3216 2240
rect 3039 2241 3040 2242
rect 3055 2241 3056 2242
rect 3045 2243 3046 2244
rect 3061 2243 3062 2244
rect 3012 2245 3013 2246
rect 3046 2245 3047 2246
rect 3003 2247 3004 2248
rect 3013 2247 3014 2248
rect 3004 2249 3005 2250
rect 3150 2249 3151 2250
rect 3063 2251 3064 2252
rect 3088 2251 3089 2252
rect 3073 2253 3074 2254
rect 3159 2253 3160 2254
rect 3079 2255 3080 2256
rect 3257 2255 3258 2256
rect 3096 2257 3097 2258
rect 3139 2257 3140 2258
rect 3105 2259 3106 2260
rect 3160 2259 3161 2260
rect 3106 2261 3107 2262
rect 3151 2261 3152 2262
rect 3112 2263 3113 2264
rect 3178 2263 3179 2264
rect 3118 2265 3119 2266
rect 3141 2265 3142 2266
rect 3081 2267 3082 2268
rect 3142 2267 3143 2268
rect 3082 2269 3083 2270
rect 3166 2269 3167 2270
rect 3125 2271 3126 2272
rect 3163 2271 3164 2272
rect 3135 2273 3136 2274
rect 3194 2273 3195 2274
rect 3093 2275 3094 2276
rect 3136 2275 3137 2276
rect 3147 2275 3148 2276
rect 3184 2275 3185 2276
rect 3099 2277 3100 2278
rect 3148 2277 3149 2278
rect 3154 2277 3155 2278
rect 3204 2277 3205 2278
rect 3156 2279 3157 2280
rect 3174 2279 3175 2280
rect 3157 2281 3158 2282
rect 3263 2281 3264 2282
rect 3168 2283 3169 2284
rect 3227 2283 3228 2284
rect 3171 2285 3172 2286
rect 3230 2285 3231 2286
rect 2612 2287 2613 2288
rect 3172 2287 3173 2288
rect 3181 2287 3182 2288
rect 3191 2287 3192 2288
rect 3144 2289 3145 2290
rect 3181 2289 3182 2290
rect 3084 2291 3085 2292
rect 3145 2291 3146 2292
rect 3201 2291 3202 2292
rect 3240 2291 3241 2292
rect 3270 2291 3271 2292
rect 3277 2291 3278 2292
rect 2587 2300 2588 2301
rect 2607 2300 2608 2301
rect 2610 2300 2611 2301
rect 2884 2300 2885 2301
rect 2611 2302 2612 2303
rect 2887 2302 2888 2303
rect 2623 2304 2624 2305
rect 2896 2304 2897 2305
rect 2625 2306 2626 2307
rect 2839 2306 2840 2307
rect 2628 2308 2629 2309
rect 2869 2308 2870 2309
rect 2633 2310 2634 2311
rect 2687 2310 2688 2311
rect 2632 2312 2633 2313
rect 2890 2312 2891 2313
rect 2640 2314 2641 2315
rect 2815 2314 2816 2315
rect 2650 2316 2651 2317
rect 2676 2316 2677 2317
rect 2656 2318 2657 2319
rect 2881 2318 2882 2319
rect 2679 2320 2680 2321
rect 2693 2320 2694 2321
rect 2681 2322 2682 2323
rect 2848 2322 2849 2323
rect 2694 2324 2695 2325
rect 2702 2324 2703 2325
rect 2718 2324 2719 2325
rect 2860 2324 2861 2325
rect 2721 2326 2722 2327
rect 2728 2326 2729 2327
rect 2731 2326 2732 2327
rect 2733 2326 2734 2327
rect 2604 2328 2605 2329
rect 2734 2328 2735 2329
rect 2757 2328 2758 2329
rect 2899 2328 2900 2329
rect 2661 2330 2662 2331
rect 2758 2330 2759 2331
rect 2760 2330 2761 2331
rect 2788 2330 2789 2331
rect 2764 2332 2765 2333
rect 2914 2332 2915 2333
rect 2782 2334 2783 2335
rect 2794 2334 2795 2335
rect 2791 2336 2792 2337
rect 3207 2336 3208 2337
rect 2797 2338 2798 2339
rect 2926 2338 2927 2339
rect 2812 2340 2813 2341
rect 2893 2340 2894 2341
rect 2833 2342 2834 2343
rect 2839 2342 2840 2343
rect 2821 2344 2822 2345
rect 2833 2344 2834 2345
rect 2620 2346 2621 2347
rect 2821 2346 2822 2347
rect 2836 2346 2837 2347
rect 2842 2346 2843 2347
rect 2851 2346 2852 2347
rect 2857 2346 2858 2347
rect 2590 2348 2591 2349
rect 2851 2348 2852 2349
rect 2590 2350 2591 2351
rect 2712 2350 2713 2351
rect 2854 2350 2855 2351
rect 2863 2350 2864 2351
rect 2593 2352 2594 2353
rect 2854 2352 2855 2353
rect 2872 2352 2873 2353
rect 2981 2352 2982 2353
rect 2600 2354 2601 2355
rect 2872 2354 2873 2355
rect 2878 2354 2879 2355
rect 2900 2354 2901 2355
rect 2666 2356 2667 2357
rect 2878 2356 2879 2357
rect 2891 2356 2892 2357
rect 2927 2356 2928 2357
rect 2902 2358 2903 2359
rect 2918 2358 2919 2359
rect 2653 2360 2654 2361
rect 2903 2360 2904 2361
rect 2630 2362 2631 2363
rect 2654 2362 2655 2363
rect 2905 2362 2906 2363
rect 2939 2362 2940 2363
rect 2866 2364 2867 2365
rect 2906 2364 2907 2365
rect 2742 2366 2743 2367
rect 2866 2366 2867 2367
rect 2743 2368 2744 2369
rect 2748 2368 2749 2369
rect 2924 2368 2925 2369
rect 3254 2368 3255 2369
rect 2947 2370 2948 2371
rect 3178 2370 3179 2371
rect 2884 2372 2885 2373
rect 2948 2372 2949 2373
rect 2962 2372 2963 2373
rect 2978 2372 2979 2373
rect 2971 2374 2972 2375
rect 3026 2374 3027 2375
rect 2908 2376 2909 2377
rect 2972 2376 2973 2377
rect 2984 2376 2985 2377
rect 3059 2376 3060 2377
rect 2987 2378 2988 2379
rect 3099 2378 3100 2379
rect 2998 2380 2999 2381
rect 3017 2380 3018 2381
rect 3001 2382 3002 2383
rect 3047 2382 3048 2383
rect 3004 2384 3005 2385
rect 3050 2384 3051 2385
rect 2965 2386 2966 2387
rect 3005 2386 3006 2387
rect 2953 2388 2954 2389
rect 2966 2388 2967 2389
rect 2935 2390 2936 2391
rect 2954 2390 2955 2391
rect 2845 2392 2846 2393
rect 2936 2392 2937 2393
rect 2635 2394 2636 2395
rect 2845 2394 2846 2395
rect 3007 2394 3008 2395
rect 3190 2394 3191 2395
rect 2827 2396 2828 2397
rect 3189 2396 3190 2397
rect 2682 2398 2683 2399
rect 2827 2398 2828 2399
rect 3013 2398 3014 2399
rect 3029 2398 3030 2399
rect 3019 2400 3020 2401
rect 3053 2400 3054 2401
rect 3022 2402 3023 2403
rect 3043 2402 3044 2403
rect 2974 2404 2975 2405
rect 3023 2404 3024 2405
rect 2920 2406 2921 2407
rect 2975 2406 2976 2407
rect 3037 2406 3038 2407
rect 3243 2406 3244 2407
rect 3041 2408 3042 2409
rect 3197 2408 3198 2409
rect 3055 2410 3056 2411
rect 3266 2410 3267 2411
rect 2995 2412 2996 2413
rect 3056 2412 3057 2413
rect 3067 2412 3068 2413
rect 3071 2412 3072 2413
rect 3073 2412 3074 2413
rect 3086 2412 3087 2413
rect 3076 2414 3077 2415
rect 3245 2414 3246 2415
rect 3077 2416 3078 2417
rect 3280 2416 3281 2417
rect 3079 2418 3080 2419
rect 3290 2418 3291 2419
rect 3088 2420 3089 2421
rect 3102 2420 3103 2421
rect 2950 2422 2951 2423
rect 3089 2422 3090 2423
rect 2794 2424 2795 2425
rect 2951 2424 2952 2425
rect 3106 2424 3107 2425
rect 3126 2424 3127 2425
rect 3108 2426 3109 2427
rect 3184 2426 3185 2427
rect 3112 2428 3113 2429
rect 3132 2428 3133 2429
rect 3120 2430 3121 2431
rect 3129 2430 3130 2431
rect 3142 2430 3143 2431
rect 3151 2430 3152 2431
rect 3031 2432 3032 2433
rect 3141 2432 3142 2433
rect 3136 2434 3137 2435
rect 3150 2434 3151 2435
rect 3115 2436 3116 2437
rect 3135 2436 3136 2437
rect 3145 2436 3146 2437
rect 3148 2436 3149 2437
rect 3154 2436 3155 2437
rect 3187 2436 3188 2437
rect 3139 2438 3140 2439
rect 3153 2438 3154 2439
rect 3138 2440 3139 2441
rect 3157 2440 3158 2441
rect 2875 2442 2876 2443
rect 3156 2442 3157 2443
rect 2621 2444 2622 2445
rect 2875 2444 2876 2445
rect 3163 2444 3164 2445
rect 3166 2444 3167 2445
rect 3082 2446 3083 2447
rect 3165 2446 3166 2447
rect 3160 2448 3161 2449
rect 3162 2448 3163 2449
rect 3061 2450 3062 2451
rect 3159 2450 3160 2451
rect 3172 2450 3173 2451
rect 3186 2450 3187 2451
rect 3183 2452 3184 2453
rect 3269 2452 3270 2453
rect 3201 2454 3202 2455
rect 3211 2454 3212 2455
rect 3181 2456 3182 2457
rect 3210 2456 3211 2457
rect 3218 2456 3219 2457
rect 3247 2456 3248 2457
rect 3227 2458 3228 2459
rect 3239 2458 3240 2459
rect 3174 2460 3175 2461
rect 3227 2460 3228 2461
rect 3230 2460 3231 2461
rect 3242 2460 3243 2461
rect 2593 2469 2594 2470
rect 2915 2469 2916 2470
rect 2600 2471 2601 2472
rect 2851 2471 2852 2472
rect 2600 2473 2601 2474
rect 2731 2473 2732 2474
rect 2604 2475 2605 2476
rect 2848 2475 2849 2476
rect 2603 2477 2604 2478
rect 2771 2477 2772 2478
rect 2607 2479 2608 2480
rect 2912 2479 2913 2480
rect 2587 2481 2588 2482
rect 2606 2481 2607 2482
rect 2618 2481 2619 2482
rect 2849 2481 2850 2482
rect 2625 2483 2626 2484
rect 2857 2483 2858 2484
rect 2630 2485 2631 2486
rect 2640 2485 2641 2486
rect 2635 2487 2636 2488
rect 2852 2487 2853 2488
rect 2642 2489 2643 2490
rect 2897 2489 2898 2490
rect 2658 2491 2659 2492
rect 2743 2491 2744 2492
rect 2661 2493 2662 2494
rect 2836 2493 2837 2494
rect 2670 2495 2671 2496
rect 2696 2495 2697 2496
rect 2673 2497 2674 2498
rect 2705 2497 2706 2498
rect 2676 2499 2677 2500
rect 2819 2499 2820 2500
rect 2679 2501 2680 2502
rect 2687 2501 2688 2502
rect 2682 2503 2683 2504
rect 2815 2503 2816 2504
rect 2626 2505 2627 2506
rect 2816 2505 2817 2506
rect 2681 2507 2682 2508
rect 2878 2507 2879 2508
rect 2694 2509 2695 2510
rect 2738 2509 2739 2510
rect 2702 2511 2703 2512
rect 2918 2511 2919 2512
rect 2712 2513 2713 2514
rect 2732 2513 2733 2514
rect 2714 2515 2715 2516
rect 2812 2515 2813 2516
rect 2726 2517 2727 2518
rect 2854 2517 2855 2518
rect 2728 2519 2729 2520
rect 3253 2519 3254 2520
rect 2734 2521 2735 2522
rect 2774 2521 2775 2522
rect 2750 2523 2751 2524
rect 2948 2523 2949 2524
rect 2776 2525 2777 2526
rect 2804 2525 2805 2526
rect 2619 2527 2620 2528
rect 2777 2527 2778 2528
rect 2800 2527 2801 2528
rect 2909 2527 2910 2528
rect 2755 2529 2756 2530
rect 2801 2529 2802 2530
rect 2581 2531 2582 2532
rect 2756 2531 2757 2532
rect 2827 2531 2828 2532
rect 2858 2531 2859 2532
rect 2839 2533 2840 2534
rect 2882 2533 2883 2534
rect 2845 2535 2846 2536
rect 2894 2535 2895 2536
rect 2809 2537 2810 2538
rect 2846 2537 2847 2538
rect 2869 2537 2870 2538
rect 2918 2537 2919 2538
rect 2833 2539 2834 2540
rect 2870 2539 2871 2540
rect 2872 2539 2873 2540
rect 2921 2539 2922 2540
rect 2758 2541 2759 2542
rect 2873 2541 2874 2542
rect 2759 2543 2760 2544
rect 2782 2543 2783 2544
rect 2888 2543 2889 2544
rect 2966 2543 2967 2544
rect 2633 2545 2634 2546
rect 2888 2545 2889 2546
rect 2900 2545 2901 2546
rect 2948 2545 2949 2546
rect 2863 2547 2864 2548
rect 2900 2547 2901 2548
rect 2821 2549 2822 2550
rect 2864 2549 2865 2550
rect 2924 2549 2925 2550
rect 2984 2549 2985 2550
rect 2875 2551 2876 2552
rect 2924 2551 2925 2552
rect 2930 2551 2931 2552
rect 2990 2551 2991 2552
rect 2685 2553 2686 2554
rect 2930 2553 2931 2554
rect 2933 2553 2934 2554
rect 2993 2553 2994 2554
rect 2936 2555 2937 2556
rect 2966 2555 2967 2556
rect 2831 2557 2832 2558
rect 2936 2557 2937 2558
rect 2939 2557 2940 2558
rect 2969 2557 2970 2558
rect 2954 2559 2955 2560
rect 2996 2559 2997 2560
rect 2623 2561 2624 2562
rect 2954 2561 2955 2562
rect 2972 2561 2973 2562
rect 3002 2561 3003 2562
rect 2975 2563 2976 2564
rect 3011 2563 3012 2564
rect 2978 2565 2979 2566
rect 3020 2565 3021 2566
rect 2951 2567 2952 2568
rect 2978 2567 2979 2568
rect 2903 2569 2904 2570
rect 2951 2569 2952 2570
rect 2866 2571 2867 2572
rect 2903 2571 2904 2572
rect 2987 2571 2988 2572
rect 3113 2571 3114 2572
rect 2927 2573 2928 2574
rect 2987 2573 2988 2574
rect 2584 2575 2585 2576
rect 2927 2575 2928 2576
rect 3005 2575 3006 2576
rect 3035 2575 3036 2576
rect 2891 2577 2892 2578
rect 3005 2577 3006 2578
rect 3017 2577 3018 2578
rect 3092 2577 3093 2578
rect 2960 2579 2961 2580
rect 3017 2579 3018 2580
rect 2906 2581 2907 2582
rect 2960 2581 2961 2582
rect 2596 2583 2597 2584
rect 2906 2583 2907 2584
rect 3023 2583 3024 2584
rect 3062 2583 3063 2584
rect 3026 2585 3027 2586
rect 3059 2585 3060 2586
rect 3029 2587 3030 2588
rect 3083 2587 3084 2588
rect 3041 2589 3042 2590
rect 3234 2589 3235 2590
rect 3044 2591 3045 2592
rect 3099 2591 3100 2592
rect 3047 2593 3048 2594
rect 3155 2593 3156 2594
rect 3050 2595 3051 2596
rect 3179 2595 3180 2596
rect 2981 2597 2982 2598
rect 3050 2597 3051 2598
rect 2753 2599 2754 2600
rect 2981 2599 2982 2600
rect 3053 2599 3054 2600
rect 3089 2599 3090 2600
rect 2654 2601 2655 2602
rect 3053 2601 3054 2602
rect 3056 2601 3057 2602
rect 3092 2601 3093 2602
rect 3056 2603 3057 2604
rect 3129 2603 3130 2604
rect 3071 2605 3072 2606
rect 3122 2605 3123 2606
rect 3077 2607 3078 2608
rect 3287 2607 3288 2608
rect 3077 2609 3078 2610
rect 3262 2609 3263 2610
rect 3086 2611 3087 2612
rect 3146 2611 3147 2612
rect 3102 2613 3103 2614
rect 3158 2613 3159 2614
rect 3038 2615 3039 2616
rect 3101 2615 3102 2616
rect 3119 2615 3120 2616
rect 3141 2615 3142 2616
rect 3126 2617 3127 2618
rect 3201 2617 3202 2618
rect 3128 2619 3129 2620
rect 3135 2619 3136 2620
rect 3132 2621 3133 2622
rect 3213 2621 3214 2622
rect 3131 2623 3132 2624
rect 3259 2623 3260 2624
rect 3134 2625 3135 2626
rect 3273 2625 3274 2626
rect 3138 2627 3139 2628
rect 3269 2627 3270 2628
rect 3143 2629 3144 2630
rect 3290 2629 3291 2630
rect 3150 2631 3151 2632
rect 3194 2631 3195 2632
rect 3149 2633 3150 2634
rect 3248 2633 3249 2634
rect 3153 2635 3154 2636
rect 3197 2635 3198 2636
rect 2876 2637 2877 2638
rect 3152 2637 3153 2638
rect 3174 2637 3175 2638
rect 3225 2637 3226 2638
rect 3204 2639 3205 2640
rect 3220 2639 3221 2640
rect 3168 2641 3169 2642
rect 3203 2641 3204 2642
rect 3183 2643 3184 2644
rect 3219 2643 3220 2644
rect 3162 2645 3163 2646
rect 3182 2645 3183 2646
rect 3207 2645 3208 2646
rect 3272 2645 3273 2646
rect 3210 2647 3211 2648
rect 3275 2647 3276 2648
rect 3041 2649 3042 2650
rect 3210 2649 3211 2650
rect 3216 2649 3217 2650
rect 3244 2649 3245 2650
rect 3223 2651 3224 2652
rect 3281 2651 3282 2652
rect 3186 2653 3187 2654
rect 3222 2653 3223 2654
rect 3165 2655 3166 2656
rect 3185 2655 3186 2656
rect 3108 2657 3109 2658
rect 3164 2657 3165 2658
rect 3228 2657 3229 2658
rect 3278 2657 3279 2658
rect 3239 2659 3240 2660
rect 3290 2659 3291 2660
rect 3242 2661 3243 2662
rect 3293 2661 3294 2662
rect 3303 2661 3304 2662
rect 3317 2661 3318 2662
rect 2584 2670 2585 2671
rect 2765 2670 2766 2671
rect 2596 2672 2597 2673
rect 2918 2672 2919 2673
rect 2606 2674 2607 2675
rect 2613 2674 2614 2675
rect 2581 2676 2582 2677
rect 2607 2676 2608 2677
rect 2609 2676 2610 2677
rect 2822 2676 2823 2677
rect 2616 2678 2617 2679
rect 2921 2678 2922 2679
rect 2619 2680 2620 2681
rect 2714 2680 2715 2681
rect 2603 2682 2604 2683
rect 2619 2682 2620 2683
rect 2623 2682 2624 2683
rect 2900 2682 2901 2683
rect 2633 2684 2634 2685
rect 2677 2684 2678 2685
rect 2637 2686 2638 2687
rect 3116 2686 3117 2687
rect 2647 2688 2648 2689
rect 2858 2688 2859 2689
rect 2654 2690 2655 2691
rect 2945 2690 2946 2691
rect 2658 2692 2659 2693
rect 2900 2692 2901 2693
rect 2672 2694 2673 2695
rect 2966 2694 2967 2695
rect 2683 2696 2684 2697
rect 2687 2696 2688 2697
rect 2681 2698 2682 2699
rect 2686 2698 2687 2699
rect 2693 2698 2694 2699
rect 2870 2698 2871 2699
rect 2692 2700 2693 2701
rect 2696 2700 2697 2701
rect 2702 2700 2703 2701
rect 2852 2700 2853 2701
rect 2705 2702 2706 2703
rect 2714 2702 2715 2703
rect 2723 2702 2724 2703
rect 2726 2702 2727 2703
rect 2729 2702 2730 2703
rect 2732 2702 2733 2703
rect 2738 2702 2739 2703
rect 2741 2702 2742 2703
rect 2747 2702 2748 2703
rect 2954 2702 2955 2703
rect 2669 2704 2670 2705
rect 2954 2704 2955 2705
rect 2668 2706 2669 2707
rect 2972 2706 2973 2707
rect 2756 2708 2757 2709
rect 2762 2708 2763 2709
rect 2768 2708 2769 2709
rect 2777 2708 2778 2709
rect 2771 2710 2772 2711
rect 2780 2710 2781 2711
rect 2774 2712 2775 2713
rect 3296 2712 3297 2713
rect 2786 2714 2787 2715
rect 3014 2714 3015 2715
rect 2789 2716 2790 2717
rect 2873 2716 2874 2717
rect 2792 2718 2793 2719
rect 2951 2718 2952 2719
rect 2798 2720 2799 2721
rect 2801 2720 2802 2721
rect 2801 2722 2802 2723
rect 2903 2722 2904 2723
rect 2600 2724 2601 2725
rect 2903 2724 2904 2725
rect 2831 2726 2832 2727
rect 2930 2726 2931 2727
rect 2840 2728 2841 2729
rect 2846 2728 2847 2729
rect 2849 2728 2850 2729
rect 2921 2728 2922 2729
rect 2849 2730 2850 2731
rect 3002 2730 3003 2731
rect 2661 2732 2662 2733
rect 3002 2732 3003 2733
rect 2852 2734 2853 2735
rect 2864 2734 2865 2735
rect 2870 2734 2871 2735
rect 2882 2734 2883 2735
rect 2876 2736 2877 2737
rect 2894 2736 2895 2737
rect 2654 2738 2655 2739
rect 2894 2738 2895 2739
rect 2879 2740 2880 2741
rect 3005 2740 3006 2741
rect 2882 2742 2883 2743
rect 2906 2742 2907 2743
rect 2885 2744 2886 2745
rect 2909 2744 2910 2745
rect 2888 2746 2889 2747
rect 2930 2746 2931 2747
rect 2888 2748 2889 2749
rect 2912 2748 2913 2749
rect 2637 2750 2638 2751
rect 2912 2750 2913 2751
rect 2891 2752 2892 2753
rect 2915 2752 2916 2753
rect 2906 2754 2907 2755
rect 2924 2754 2925 2755
rect 2909 2756 2910 2757
rect 2927 2756 2928 2757
rect 2942 2756 2943 2757
rect 2948 2756 2949 2757
rect 2951 2756 2952 2757
rect 3191 2756 3192 2757
rect 2960 2758 2961 2759
rect 3008 2758 3009 2759
rect 2960 2760 2961 2761
rect 2984 2760 2985 2761
rect 2834 2762 2835 2763
rect 2984 2762 2985 2763
rect 2966 2764 2967 2765
rect 2990 2764 2991 2765
rect 2837 2766 2838 2767
rect 2990 2766 2991 2767
rect 2981 2768 2982 2769
rect 3047 2768 3048 2769
rect 2981 2770 2982 2771
rect 3059 2770 3060 2771
rect 2993 2772 2994 2773
rect 3215 2772 3216 2773
rect 3011 2774 3012 2775
rect 3074 2774 3075 2775
rect 3020 2776 3021 2777
rect 3173 2776 3174 2777
rect 3020 2778 3021 2779
rect 3038 2778 3039 2779
rect 2996 2780 2997 2781
rect 3038 2780 3039 2781
rect 2996 2782 2997 2783
rect 3017 2782 3018 2783
rect 2969 2784 2970 2785
rect 3017 2784 3018 2785
rect 2699 2786 2700 2787
rect 2969 2786 2970 2787
rect 2698 2788 2699 2789
rect 2978 2788 2979 2789
rect 2978 2790 2979 2791
rect 2987 2790 2988 2791
rect 3035 2790 3036 2791
rect 3107 2790 3108 2791
rect 3044 2792 3045 2793
rect 3068 2792 3069 2793
rect 2750 2794 2751 2795
rect 3044 2794 3045 2795
rect 3056 2794 3057 2795
rect 3265 2794 3266 2795
rect 3041 2796 3042 2797
rect 3056 2796 3057 2797
rect 3059 2796 3060 2797
rect 3104 2796 3105 2797
rect 3083 2798 3084 2799
rect 3110 2798 3111 2799
rect 3104 2800 3105 2801
rect 3176 2800 3177 2801
rect 2936 2802 2937 2803
rect 3176 2802 3177 2803
rect 3125 2804 3126 2805
rect 3155 2804 3156 2805
rect 3119 2806 3120 2807
rect 3155 2806 3156 2807
rect 3128 2808 3129 2809
rect 3262 2808 3263 2809
rect 3134 2810 3135 2811
rect 3330 2810 3331 2811
rect 3137 2812 3138 2813
rect 3206 2812 3207 2813
rect 3143 2814 3144 2815
rect 3170 2814 3171 2815
rect 3131 2816 3132 2817
rect 3143 2816 3144 2817
rect 3149 2816 3150 2817
rect 3188 2816 3189 2817
rect 3089 2818 3090 2819
rect 3149 2818 3150 2819
rect 3158 2818 3159 2819
rect 3234 2818 3235 2819
rect 3182 2820 3183 2821
rect 3240 2820 3241 2821
rect 3194 2822 3195 2823
rect 3317 2822 3318 2823
rect 3053 2824 3054 2825
rect 3194 2824 3195 2825
rect 2759 2826 2760 2827
rect 3053 2826 3054 2827
rect 2644 2828 2645 2829
rect 2759 2828 2760 2829
rect 2644 2830 2645 2831
rect 2918 2830 2919 2831
rect 3197 2830 3198 2831
rect 3314 2830 3315 2831
rect 3164 2832 3165 2833
rect 3197 2832 3198 2833
rect 3122 2834 3123 2835
rect 3164 2834 3165 2835
rect 3203 2834 3204 2835
rect 3234 2834 3235 2835
rect 3225 2836 3226 2837
rect 3278 2836 3279 2837
rect 3228 2838 3229 2839
rect 3281 2838 3282 2839
rect 3231 2840 3232 2841
rect 3268 2840 3269 2841
rect 3238 2842 3239 2843
rect 3246 2842 3247 2843
rect 3152 2844 3153 2845
rect 3237 2844 3238 2845
rect 3092 2846 3093 2847
rect 3152 2846 3153 2847
rect 3092 2848 3093 2849
rect 3324 2848 3325 2849
rect 3244 2850 3245 2851
rect 3381 2850 3382 2851
rect 3185 2852 3186 2853
rect 3243 2852 3244 2853
rect 3146 2854 3147 2855
rect 3185 2854 3186 2855
rect 3077 2856 3078 2857
rect 3146 2856 3147 2857
rect 3253 2856 3254 2857
rect 3308 2856 3309 2857
rect 3252 2858 3253 2859
rect 3339 2858 3340 2859
rect 3272 2860 3273 2861
rect 3333 2860 3334 2861
rect 3210 2862 3211 2863
rect 3272 2862 3273 2863
rect 3275 2862 3276 2863
rect 3336 2862 3337 2863
rect 3290 2864 3291 2865
rect 3358 2864 3359 2865
rect 3219 2866 3220 2867
rect 3290 2866 3291 2867
rect 3293 2866 3294 2867
rect 3361 2866 3362 2867
rect 3222 2868 3223 2869
rect 3293 2868 3294 2869
rect 3113 2870 3114 2871
rect 3222 2870 3223 2871
rect 3050 2872 3051 2873
rect 3113 2872 3114 2873
rect 2846 2874 2847 2875
rect 3050 2874 3051 2875
rect 3299 2874 3300 2875
rect 3303 2874 3304 2875
rect 3388 2874 3389 2875
rect 3395 2874 3396 2875
rect 2539 2883 2540 2884
rect 2546 2883 2547 2884
rect 2588 2883 2589 2884
rect 2765 2883 2766 2884
rect 2591 2885 2592 2886
rect 2888 2885 2889 2886
rect 2590 2887 2591 2888
rect 2762 2887 2763 2888
rect 2598 2889 2599 2890
rect 2932 2889 2933 2890
rect 2602 2891 2603 2892
rect 2761 2891 2762 2892
rect 2605 2893 2606 2894
rect 2607 2893 2608 2894
rect 2608 2895 2609 2896
rect 2613 2895 2614 2896
rect 2611 2897 2612 2898
rect 2719 2897 2720 2898
rect 2623 2899 2624 2900
rect 2891 2899 2892 2900
rect 2630 2901 2631 2902
rect 2909 2901 2910 2902
rect 2640 2903 2641 2904
rect 2737 2903 2738 2904
rect 2644 2905 2645 2906
rect 2912 2905 2913 2906
rect 2644 2907 2645 2908
rect 2759 2907 2760 2908
rect 2651 2909 2652 2910
rect 2866 2909 2867 2910
rect 2647 2911 2648 2912
rect 2651 2911 2652 2912
rect 2647 2913 2648 2914
rect 2872 2913 2873 2914
rect 2654 2915 2655 2916
rect 2876 2915 2877 2916
rect 2658 2917 2659 2918
rect 2852 2917 2853 2918
rect 2658 2919 2659 2920
rect 2974 2919 2975 2920
rect 2661 2921 2662 2922
rect 2914 2921 2915 2922
rect 2661 2923 2662 2924
rect 2741 2923 2742 2924
rect 2665 2925 2666 2926
rect 2897 2925 2898 2926
rect 2673 2927 2674 2928
rect 2894 2927 2895 2928
rect 2677 2929 2678 2930
rect 2911 2929 2912 2930
rect 2683 2931 2684 2932
rect 2688 2931 2689 2932
rect 2682 2933 2683 2934
rect 2686 2933 2687 2934
rect 2692 2933 2693 2934
rect 2694 2933 2695 2934
rect 2575 2935 2576 2936
rect 2691 2935 2692 2936
rect 2698 2935 2699 2936
rect 2935 2935 2936 2936
rect 2700 2937 2701 2938
rect 2926 2937 2927 2938
rect 2702 2939 2703 2940
rect 2969 2939 2970 2940
rect 2710 2941 2711 2942
rect 2714 2941 2715 2942
rect 2723 2941 2724 2942
rect 2734 2941 2735 2942
rect 2729 2943 2730 2944
rect 2731 2943 2732 2944
rect 2747 2943 2748 2944
rect 2978 2943 2979 2944
rect 2750 2945 2751 2946
rect 2801 2945 2802 2946
rect 2768 2947 2769 2948
rect 2785 2947 2786 2948
rect 2767 2949 2768 2950
rect 2903 2949 2904 2950
rect 2773 2951 2774 2952
rect 2780 2951 2781 2952
rect 2792 2951 2793 2952
rect 2800 2951 2801 2952
rect 2791 2953 2792 2954
rect 2798 2953 2799 2954
rect 2804 2953 2805 2954
rect 2836 2953 2837 2954
rect 2806 2955 2807 2956
rect 2816 2955 2817 2956
rect 2812 2957 2813 2958
rect 2822 2957 2823 2958
rect 2819 2959 2820 2960
rect 2821 2959 2822 2960
rect 2752 2961 2753 2962
rect 2818 2961 2819 2962
rect 2830 2961 2831 2962
rect 2840 2961 2841 2962
rect 2834 2963 2835 2964
rect 3002 2963 3003 2964
rect 2870 2965 2871 2966
rect 2875 2965 2876 2966
rect 2878 2965 2879 2966
rect 2930 2965 2931 2966
rect 2882 2967 2883 2968
rect 2890 2967 2891 2968
rect 2885 2969 2886 2970
rect 2893 2969 2894 2970
rect 2884 2971 2885 2972
rect 2918 2971 2919 2972
rect 2887 2973 2888 2974
rect 2921 2973 2922 2974
rect 2900 2975 2901 2976
rect 2902 2975 2903 2976
rect 2906 2975 2907 2976
rect 2908 2975 2909 2976
rect 2616 2977 2617 2978
rect 2905 2977 2906 2978
rect 2920 2977 2921 2978
rect 2942 2977 2943 2978
rect 2923 2979 2924 2980
rect 2945 2979 2946 2980
rect 2941 2981 2942 2982
rect 3008 2981 3009 2982
rect 2947 2983 2948 2984
rect 3014 2983 3015 2984
rect 2951 2985 2952 2986
rect 3007 2985 3008 2986
rect 2966 2987 2967 2988
rect 2977 2987 2978 2988
rect 2960 2989 2961 2990
rect 2965 2989 2966 2990
rect 2954 2991 2955 2992
rect 2959 2991 2960 2992
rect 2984 2991 2985 2992
rect 3268 2991 3269 2992
rect 2848 2993 2849 2994
rect 2983 2993 2984 2994
rect 2992 2993 2993 2994
rect 3017 2993 3018 2994
rect 2996 2995 2997 2996
rect 3013 2995 3014 2996
rect 2990 2997 2991 2998
rect 2995 2997 2996 2998
rect 2749 2999 2750 3000
rect 2989 2999 2990 3000
rect 3020 2999 3021 3000
rect 3031 2999 3032 3000
rect 3019 3001 3020 3002
rect 3044 3001 3045 3002
rect 3022 3003 3023 3004
rect 3047 3003 3048 3004
rect 3025 3005 3026 3006
rect 3050 3005 3051 3006
rect 3028 3007 3029 3008
rect 3053 3007 3054 3008
rect 3038 3009 3039 3010
rect 3094 3009 3095 3010
rect 3037 3011 3038 3012
rect 3116 3011 3117 3012
rect 3043 3013 3044 3014
rect 3265 3013 3266 3014
rect 3056 3015 3057 3016
rect 3064 3015 3065 3016
rect 3055 3017 3056 3018
rect 3364 3017 3365 3018
rect 3059 3019 3060 3020
rect 3225 3019 3226 3020
rect 3061 3021 3062 3022
rect 3215 3021 3216 3022
rect 3074 3023 3075 3024
rect 3076 3023 3077 3024
rect 3079 3023 3080 3024
rect 3367 3023 3368 3024
rect 3085 3025 3086 3026
rect 3107 3025 3108 3026
rect 3104 3027 3105 3028
rect 3121 3027 3122 3028
rect 3092 3029 3093 3030
rect 3103 3029 3104 3030
rect 3091 3031 3092 3032
rect 3173 3031 3174 3032
rect 3125 3033 3126 3034
rect 3339 3033 3340 3034
rect 3124 3035 3125 3036
rect 3208 3035 3209 3036
rect 3133 3037 3134 3038
rect 3149 3037 3150 3038
rect 3137 3039 3138 3040
rect 3139 3039 3140 3040
rect 3136 3041 3137 3042
rect 3152 3041 3153 3042
rect 3146 3043 3147 3044
rect 3324 3043 3325 3044
rect 3143 3045 3144 3046
rect 3145 3045 3146 3046
rect 3148 3045 3149 3046
rect 3321 3045 3322 3046
rect 3155 3047 3156 3048
rect 3342 3047 3343 3048
rect 3164 3049 3165 3050
rect 3166 3049 3167 3050
rect 3163 3051 3164 3052
rect 3330 3051 3331 3052
rect 3170 3053 3171 3054
rect 3407 3053 3408 3054
rect 3172 3055 3173 3056
rect 3194 3055 3195 3056
rect 3176 3057 3177 3058
rect 3206 3057 3207 3058
rect 3113 3059 3114 3060
rect 3175 3059 3176 3060
rect 3202 3059 3203 3060
rect 3243 3059 3244 3060
rect 3218 3061 3219 3062
rect 3222 3061 3223 3062
rect 3157 3063 3158 3064
rect 3222 3063 3223 3064
rect 3232 3063 3233 3064
rect 3283 3063 3284 3064
rect 3234 3065 3235 3066
rect 3261 3065 3262 3066
rect 3235 3067 3236 3068
rect 3317 3067 3318 3068
rect 3237 3069 3238 3070
rect 3258 3069 3259 3070
rect 3110 3071 3111 3072
rect 3238 3071 3239 3072
rect 3252 3071 3253 3072
rect 3298 3071 3299 3072
rect 3259 3073 3260 3074
rect 3319 3073 3320 3074
rect 3265 3075 3266 3076
rect 3331 3075 3332 3076
rect 3286 3077 3287 3078
rect 3314 3077 3315 3078
rect 3290 3079 3291 3080
rect 3313 3079 3314 3080
rect 3278 3081 3279 3082
rect 3289 3081 3290 3082
rect 3272 3083 3273 3084
rect 3277 3083 3278 3084
rect 3293 3083 3294 3084
rect 3302 3083 3303 3084
rect 3292 3085 3293 3086
rect 3355 3085 3356 3086
rect 3295 3087 3296 3088
rect 3336 3087 3337 3088
rect 3305 3089 3306 3090
rect 3316 3089 3317 3090
rect 3308 3091 3309 3092
rect 3325 3091 3326 3092
rect 3281 3093 3282 3094
rect 3307 3093 3308 3094
rect 3240 3095 3241 3096
rect 3280 3095 3281 3096
rect 3327 3095 3328 3096
rect 3370 3095 3371 3096
rect 3333 3097 3334 3098
rect 3385 3097 3386 3098
rect 3358 3099 3359 3100
rect 3364 3099 3365 3100
rect 3361 3101 3362 3102
rect 3367 3101 3368 3102
rect 3374 3101 3375 3102
rect 3384 3101 3385 3102
rect 3381 3103 3382 3104
rect 3394 3103 3395 3104
rect 3391 3105 3392 3106
rect 3398 3105 3399 3106
rect 2578 3114 2579 3115
rect 2599 3114 2600 3115
rect 2582 3116 2583 3117
rect 2691 3116 2692 3117
rect 2587 3118 2588 3119
rect 2665 3118 2666 3119
rect 2589 3120 2590 3121
rect 2777 3120 2778 3121
rect 2596 3122 2597 3123
rect 2893 3122 2894 3123
rect 2602 3124 2603 3125
rect 2611 3124 2612 3125
rect 2605 3126 2606 3127
rect 2668 3126 2669 3127
rect 2608 3128 2609 3129
rect 2616 3128 2617 3129
rect 2610 3130 2611 3131
rect 2855 3130 2856 3131
rect 2613 3132 2614 3133
rect 2884 3132 2885 3133
rect 2623 3134 2624 3135
rect 2812 3134 2813 3135
rect 2603 3136 2604 3137
rect 2813 3136 2814 3137
rect 2626 3138 2627 3139
rect 2825 3138 2826 3139
rect 2631 3140 2632 3141
rect 2767 3140 2768 3141
rect 2640 3142 2641 3143
rect 2887 3142 2888 3143
rect 2645 3144 2646 3145
rect 2951 3144 2952 3145
rect 2662 3146 2663 3147
rect 2885 3146 2886 3147
rect 2677 3148 2678 3149
rect 2905 3148 2906 3149
rect 2686 3150 2687 3151
rect 2882 3150 2883 3151
rect 2688 3152 2689 3153
rect 2704 3152 2705 3153
rect 2700 3154 2701 3155
rect 2914 3154 2915 3155
rect 2694 3156 2695 3157
rect 2701 3156 2702 3157
rect 2682 3158 2683 3159
rect 2695 3158 2696 3159
rect 2683 3160 2684 3161
rect 3031 3160 3032 3161
rect 2707 3162 2708 3163
rect 2783 3162 2784 3163
rect 2707 3164 2708 3165
rect 2878 3164 2879 3165
rect 2710 3166 2711 3167
rect 2726 3166 2727 3167
rect 2714 3168 2715 3169
rect 3011 3168 3012 3169
rect 2719 3170 2720 3171
rect 2741 3170 2742 3171
rect 2737 3172 2738 3173
rect 2840 3172 2841 3173
rect 2734 3174 2735 3175
rect 2738 3174 2739 3175
rect 2731 3176 2732 3177
rect 2735 3176 2736 3177
rect 2752 3176 2753 3177
rect 3022 3176 3023 3177
rect 2761 3178 2762 3179
rect 2768 3178 2769 3179
rect 2765 3180 2766 3181
rect 2791 3180 2792 3181
rect 2773 3182 2774 3183
rect 2795 3182 2796 3183
rect 2527 3184 2528 3185
rect 2774 3184 2775 3185
rect 2785 3184 2786 3185
rect 2789 3184 2790 3185
rect 2786 3186 2787 3187
rect 2923 3186 2924 3187
rect 2800 3188 2801 3189
rect 2906 3188 2907 3189
rect 2804 3190 2805 3191
rect 2963 3190 2964 3191
rect 2818 3192 2819 3193
rect 2846 3192 2847 3193
rect 2647 3194 2648 3195
rect 2819 3194 2820 3195
rect 2633 3196 2634 3197
rect 2648 3196 2649 3197
rect 2821 3196 2822 3197
rect 2888 3196 2889 3197
rect 2641 3198 2642 3199
rect 2822 3198 2823 3199
rect 2828 3198 2829 3199
rect 2911 3198 2912 3199
rect 2836 3200 2837 3201
rect 2864 3200 2865 3201
rect 2830 3202 2831 3203
rect 2837 3202 2838 3203
rect 2806 3204 2807 3205
rect 2831 3204 2832 3205
rect 2843 3204 2844 3205
rect 2890 3204 2891 3205
rect 2848 3206 2849 3207
rect 2947 3206 2948 3207
rect 2852 3208 2853 3209
rect 2902 3208 2903 3209
rect 2866 3210 2867 3211
rect 2870 3210 2871 3211
rect 2872 3210 2873 3211
rect 2879 3210 2880 3211
rect 2897 3210 2898 3211
rect 3007 3210 3008 3211
rect 2903 3212 2904 3213
rect 2920 3212 2921 3213
rect 2908 3214 2909 3215
rect 3370 3214 3371 3215
rect 2909 3216 2910 3217
rect 2959 3216 2960 3217
rect 2915 3218 2916 3219
rect 2965 3218 2966 3219
rect 2921 3220 2922 3221
rect 2977 3220 2978 3221
rect 2930 3222 2931 3223
rect 2980 3222 2981 3223
rect 2658 3224 2659 3225
rect 2981 3224 2982 3225
rect 2652 3226 2653 3227
rect 2659 3226 2660 3227
rect 2935 3226 2936 3227
rect 3041 3226 3042 3227
rect 2939 3228 2940 3229
rect 2971 3228 2972 3229
rect 2941 3230 2942 3231
rect 2978 3230 2979 3231
rect 2954 3232 2955 3233
rect 2974 3232 2975 3233
rect 2957 3234 2958 3235
rect 3013 3234 3014 3235
rect 2975 3236 2976 3237
rect 2992 3236 2993 3237
rect 2983 3238 2984 3239
rect 2987 3238 2988 3239
rect 2993 3238 2994 3239
rect 3019 3238 3020 3239
rect 2999 3240 3000 3241
rect 3043 3240 3044 3241
rect 3023 3242 3024 3243
rect 3025 3242 3026 3243
rect 3028 3242 3029 3243
rect 3050 3242 3051 3243
rect 3029 3244 3030 3245
rect 3037 3244 3038 3245
rect 3035 3246 3036 3247
rect 3067 3246 3068 3247
rect 3047 3248 3048 3249
rect 3155 3248 3156 3249
rect 3055 3250 3056 3251
rect 3310 3250 3311 3251
rect 3059 3252 3060 3253
rect 3061 3252 3062 3253
rect 3064 3252 3065 3253
rect 3215 3252 3216 3253
rect 3073 3254 3074 3255
rect 3193 3254 3194 3255
rect 3077 3256 3078 3257
rect 3133 3256 3134 3257
rect 3079 3258 3080 3259
rect 3352 3258 3353 3259
rect 3080 3260 3081 3261
rect 3136 3260 3137 3261
rect 3083 3262 3084 3263
rect 3232 3262 3233 3263
rect 3094 3264 3095 3265
rect 3107 3264 3108 3265
rect 3095 3266 3096 3267
rect 3225 3266 3226 3267
rect 3098 3268 3099 3269
rect 3157 3268 3158 3269
rect 3103 3270 3104 3271
rect 3271 3270 3272 3271
rect 3091 3272 3092 3273
rect 3104 3272 3105 3273
rect 3092 3274 3093 3275
rect 3145 3274 3146 3275
rect 3121 3276 3122 3277
rect 3208 3276 3209 3277
rect 3122 3278 3123 3279
rect 3184 3278 3185 3279
rect 3128 3280 3129 3281
rect 3172 3280 3173 3281
rect 3131 3282 3132 3283
rect 3175 3282 3176 3283
rect 3134 3284 3135 3285
rect 3196 3284 3197 3285
rect 3146 3286 3147 3287
rect 3195 3286 3196 3287
rect 3148 3288 3149 3289
rect 3348 3288 3349 3289
rect 3124 3290 3125 3291
rect 3149 3290 3150 3291
rect 3125 3292 3126 3293
rect 3187 3292 3188 3293
rect 3152 3294 3153 3295
rect 3259 3294 3260 3295
rect 3163 3296 3164 3297
rect 3373 3296 3374 3297
rect 3085 3298 3086 3299
rect 3162 3298 3163 3299
rect 3086 3300 3087 3301
rect 3139 3300 3140 3301
rect 3140 3302 3141 3303
rect 3202 3302 3203 3303
rect 3168 3304 3169 3305
rect 3238 3304 3239 3305
rect 3177 3306 3178 3307
rect 3384 3306 3385 3307
rect 3186 3308 3187 3309
rect 3247 3308 3248 3309
rect 3190 3310 3191 3311
rect 3256 3310 3257 3311
rect 3216 3312 3217 3313
rect 3277 3312 3278 3313
rect 3219 3314 3220 3315
rect 3280 3314 3281 3315
rect 3229 3316 3230 3317
rect 3307 3316 3308 3317
rect 3238 3318 3239 3319
rect 3298 3318 3299 3319
rect 3241 3320 3242 3321
rect 3289 3320 3290 3321
rect 3253 3322 3254 3323
rect 3259 3322 3260 3323
rect 3262 3322 3263 3323
rect 3313 3322 3314 3323
rect 3265 3324 3266 3325
rect 3322 3324 3323 3325
rect 3265 3326 3266 3327
rect 3325 3326 3326 3327
rect 2875 3328 2876 3329
rect 3324 3328 3325 3329
rect 2876 3330 2877 3331
rect 2932 3330 2933 3331
rect 2933 3332 2934 3333
rect 2989 3332 2990 3333
rect 3304 3332 3305 3333
rect 3364 3332 3365 3333
rect 3307 3334 3308 3335
rect 3367 3334 3368 3335
rect 3310 3336 3311 3337
rect 3331 3336 3332 3337
rect 3316 3338 3317 3339
rect 3380 3338 3381 3339
rect 3166 3340 3167 3341
rect 3317 3340 3318 3341
rect 3165 3342 3166 3343
rect 3235 3342 3236 3343
rect 3235 3344 3236 3345
rect 3295 3344 3296 3345
rect 3244 3346 3245 3347
rect 3295 3346 3296 3347
rect 2588 3355 2589 3356
rect 2749 3355 2750 3356
rect 2602 3357 2603 3358
rect 2627 3357 2628 3358
rect 2609 3359 2610 3360
rect 2876 3359 2877 3360
rect 2631 3361 2632 3362
rect 2825 3361 2826 3362
rect 2634 3363 2635 3364
rect 2948 3363 2949 3364
rect 2616 3365 2617 3366
rect 2633 3365 2634 3366
rect 2638 3365 2639 3366
rect 2698 3365 2699 3366
rect 2648 3367 2649 3368
rect 2791 3367 2792 3368
rect 2652 3369 2653 3370
rect 2879 3369 2880 3370
rect 2659 3371 2660 3372
rect 2906 3371 2907 3372
rect 2658 3373 2659 3374
rect 2789 3373 2790 3374
rect 2662 3375 2663 3376
rect 2924 3375 2925 3376
rect 2665 3377 2666 3378
rect 2680 3377 2681 3378
rect 2668 3379 2669 3380
rect 2683 3379 2684 3380
rect 2674 3381 2675 3382
rect 2722 3381 2723 3382
rect 2677 3383 2678 3384
rect 2692 3383 2693 3384
rect 2686 3385 2687 3386
rect 2909 3385 2910 3386
rect 2701 3387 2702 3388
rect 2716 3387 2717 3388
rect 2710 3389 2711 3390
rect 2918 3389 2919 3390
rect 2695 3391 2696 3392
rect 2710 3391 2711 3392
rect 2719 3391 2720 3392
rect 2731 3391 2732 3392
rect 2735 3391 2736 3392
rect 2746 3391 2747 3392
rect 2734 3393 2735 3394
rect 3026 3393 3027 3394
rect 2765 3395 2766 3396
rect 2809 3395 2810 3396
rect 2770 3397 2771 3398
rect 2828 3397 2829 3398
rect 2777 3399 2778 3400
rect 2797 3399 2798 3400
rect 2779 3401 2780 3402
rect 2875 3401 2876 3402
rect 2783 3403 2784 3404
rect 2927 3403 2928 3404
rect 2782 3405 2783 3406
rect 2857 3405 2858 3406
rect 2786 3407 2787 3408
rect 3017 3407 3018 3408
rect 2768 3409 2769 3410
rect 2785 3409 2786 3410
rect 2741 3411 2742 3412
rect 2767 3411 2768 3412
rect 2738 3413 2739 3414
rect 2740 3413 2741 3414
rect 2737 3415 2738 3416
rect 2759 3415 2760 3416
rect 2726 3417 2727 3418
rect 2758 3417 2759 3418
rect 2795 3417 2796 3418
rect 2827 3417 2828 3418
rect 2704 3419 2705 3420
rect 2794 3419 2795 3420
rect 2803 3419 2804 3420
rect 2993 3419 2994 3420
rect 2815 3421 2816 3422
rect 2975 3421 2976 3422
rect 2831 3423 2832 3424
rect 2833 3423 2834 3424
rect 2840 3423 2841 3424
rect 2872 3423 2873 3424
rect 2839 3425 2840 3426
rect 2846 3425 2847 3426
rect 2813 3427 2814 3428
rect 2845 3427 2846 3428
rect 2852 3427 2853 3428
rect 2912 3427 2913 3428
rect 2819 3429 2820 3430
rect 2851 3429 2852 3430
rect 2774 3431 2775 3432
rect 2818 3431 2819 3432
rect 2885 3431 2886 3432
rect 2936 3431 2937 3432
rect 2897 3433 2898 3434
rect 3020 3433 3021 3434
rect 2900 3435 2901 3436
rect 2987 3435 2988 3436
rect 2843 3437 2844 3438
rect 2900 3437 2901 3438
rect 2903 3437 2904 3438
rect 2960 3437 2961 3438
rect 2595 3439 2596 3440
rect 2903 3439 2904 3440
rect 2915 3439 2916 3440
rect 2990 3439 2991 3440
rect 2855 3441 2856 3442
rect 2915 3441 2916 3442
rect 2822 3443 2823 3444
rect 2854 3443 2855 3444
rect 2933 3443 2934 3444
rect 3014 3443 3015 3444
rect 2882 3445 2883 3446
rect 2933 3445 2934 3446
rect 2942 3445 2943 3446
rect 2951 3445 2952 3446
rect 2954 3445 2955 3446
rect 2993 3445 2994 3446
rect 2613 3447 2614 3448
rect 2954 3447 2955 3448
rect 2957 3447 2958 3448
rect 3032 3447 3033 3448
rect 2585 3449 2586 3450
rect 2957 3449 2958 3450
rect 2963 3449 2964 3450
rect 3059 3449 3060 3450
rect 2864 3451 2865 3452
rect 2963 3451 2964 3452
rect 2966 3451 2967 3452
rect 3062 3451 3063 3452
rect 2978 3453 2979 3454
rect 2984 3453 2985 3454
rect 2939 3455 2940 3456
rect 2978 3455 2979 3456
rect 2888 3457 2889 3458
rect 2939 3457 2940 3458
rect 2999 3457 3000 3458
rect 3195 3457 3196 3458
rect 2930 3459 2931 3460
rect 2999 3459 3000 3460
rect 2870 3461 2871 3462
rect 2930 3461 2931 3462
rect 2837 3463 2838 3464
rect 2869 3463 2870 3464
rect 3008 3463 3009 3464
rect 3023 3463 3024 3464
rect 2996 3465 2997 3466
rect 3023 3465 3024 3466
rect 2921 3467 2922 3468
rect 2996 3467 2997 3468
rect 3011 3467 3012 3468
rect 3062 3467 3063 3468
rect 3029 3469 3030 3470
rect 3155 3469 3156 3470
rect 3041 3471 3042 3472
rect 3071 3471 3072 3472
rect 3047 3473 3048 3474
rect 3068 3473 3069 3474
rect 3050 3475 3051 3476
rect 3232 3475 3233 3476
rect 2981 3477 2982 3478
rect 3050 3477 3051 3478
rect 3083 3477 3084 3478
rect 3116 3477 3117 3478
rect 3086 3479 3087 3480
rect 3179 3479 3180 3480
rect 3086 3481 3087 3482
rect 3162 3481 3163 3482
rect 3095 3483 3096 3484
rect 3155 3483 3156 3484
rect 3098 3485 3099 3486
rect 3119 3485 3120 3486
rect 3125 3485 3126 3486
rect 3331 3485 3332 3486
rect 3092 3487 3093 3488
rect 3125 3487 3126 3488
rect 3134 3487 3135 3488
rect 3269 3487 3270 3488
rect 3140 3489 3141 3490
rect 3170 3489 3171 3490
rect 3146 3491 3147 3492
rect 3182 3491 3183 3492
rect 3104 3493 3105 3494
rect 3146 3493 3147 3494
rect 3077 3495 3078 3496
rect 3104 3495 3105 3496
rect 3152 3495 3153 3496
rect 3327 3495 3328 3496
rect 3165 3497 3166 3498
rect 3206 3497 3207 3498
rect 3128 3499 3129 3500
rect 3164 3499 3165 3500
rect 3128 3501 3129 3502
rect 3345 3501 3346 3502
rect 3168 3503 3169 3504
rect 3209 3503 3210 3504
rect 3131 3505 3132 3506
rect 3167 3505 3168 3506
rect 3177 3505 3178 3506
rect 3224 3505 3225 3506
rect 3122 3507 3123 3508
rect 3176 3507 3177 3508
rect 3188 3507 3189 3508
rect 3192 3507 3193 3508
rect 3044 3509 3045 3510
rect 3191 3509 3192 3510
rect 3216 3509 3217 3510
rect 3272 3509 3273 3510
rect 3238 3511 3239 3512
rect 3334 3511 3335 3512
rect 3241 3513 3242 3514
rect 3278 3513 3279 3514
rect 3244 3515 3245 3516
rect 3281 3515 3282 3516
rect 3253 3517 3254 3518
rect 3291 3517 3292 3518
rect 3259 3519 3260 3520
rect 3312 3519 3313 3520
rect 3256 3521 3257 3522
rect 3260 3521 3261 3522
rect 3257 3523 3258 3524
rect 3274 3523 3275 3524
rect 3219 3525 3220 3526
rect 3275 3525 3276 3526
rect 3186 3527 3187 3528
rect 3218 3527 3219 3528
rect 3149 3529 3150 3530
rect 3185 3529 3186 3530
rect 3107 3531 3108 3532
rect 3149 3531 3150 3532
rect 3080 3533 3081 3534
rect 3107 3533 3108 3534
rect 3035 3535 3036 3536
rect 3080 3535 3081 3536
rect 3263 3535 3264 3536
rect 3370 3535 3371 3536
rect 3265 3537 3266 3538
rect 3318 3537 3319 3538
rect 3235 3539 3236 3540
rect 3266 3539 3267 3540
rect 3304 3539 3305 3540
rect 3357 3539 3358 3540
rect 3239 3541 3240 3542
rect 3305 3541 3306 3542
rect 3307 3541 3308 3542
rect 3360 3541 3361 3542
rect 3373 3541 3374 3542
rect 3377 3541 3378 3542
rect 2530 3550 2531 3551
rect 2761 3550 2762 3551
rect 2541 3552 2542 3553
rect 2677 3552 2678 3553
rect 2561 3554 2562 3555
rect 2642 3554 2643 3555
rect 2564 3556 2565 3557
rect 2575 3556 2576 3557
rect 2581 3556 2582 3557
rect 2680 3556 2681 3557
rect 2584 3558 2585 3559
rect 2686 3558 2687 3559
rect 2588 3560 2589 3561
rect 2683 3560 2684 3561
rect 2595 3562 2596 3563
rect 3170 3562 3171 3563
rect 2594 3564 2595 3565
rect 2900 3564 2901 3565
rect 2605 3566 2606 3567
rect 2915 3566 2916 3567
rect 2604 3568 2605 3569
rect 2836 3568 2837 3569
rect 2609 3570 2610 3571
rect 2698 3570 2699 3571
rect 2608 3572 2609 3573
rect 2863 3572 2864 3573
rect 2612 3574 2613 3575
rect 2954 3574 2955 3575
rect 2615 3576 2616 3577
rect 2636 3576 2637 3577
rect 2639 3576 2640 3577
rect 2767 3576 2768 3577
rect 2633 3578 2634 3579
rect 2639 3578 2640 3579
rect 2648 3578 2649 3579
rect 2842 3578 2843 3579
rect 2651 3580 2652 3581
rect 2851 3580 2852 3581
rect 2652 3582 2653 3583
rect 2887 3582 2888 3583
rect 2667 3584 2668 3585
rect 2933 3584 2934 3585
rect 2667 3586 2668 3587
rect 2890 3586 2891 3587
rect 2670 3588 2671 3589
rect 2725 3588 2726 3589
rect 2671 3590 2672 3591
rect 2924 3590 2925 3591
rect 2674 3592 2675 3593
rect 2740 3592 2741 3593
rect 2674 3594 2675 3595
rect 2930 3594 2931 3595
rect 2692 3596 2693 3597
rect 2698 3596 2699 3597
rect 2695 3598 2696 3599
rect 2716 3598 2717 3599
rect 2658 3600 2659 3601
rect 2716 3600 2717 3601
rect 2710 3602 2711 3603
rect 2722 3602 2723 3603
rect 2719 3604 2720 3605
rect 2731 3604 2732 3605
rect 2734 3604 2735 3605
rect 2948 3604 2949 3605
rect 2734 3606 2735 3607
rect 2770 3606 2771 3607
rect 2737 3608 2738 3609
rect 2767 3608 2768 3609
rect 2740 3610 2741 3611
rect 2746 3610 2747 3611
rect 2743 3612 2744 3613
rect 2749 3612 2750 3613
rect 2758 3612 2759 3613
rect 2764 3612 2765 3613
rect 2758 3614 2759 3615
rect 2809 3614 2810 3615
rect 2773 3616 2774 3617
rect 2818 3616 2819 3617
rect 2655 3618 2656 3619
rect 2818 3618 2819 3619
rect 2776 3620 2777 3621
rect 2791 3620 2792 3621
rect 2779 3622 2780 3623
rect 2794 3622 2795 3623
rect 2782 3624 2783 3625
rect 2999 3624 3000 3625
rect 2782 3626 2783 3627
rect 2785 3626 2786 3627
rect 2788 3626 2789 3627
rect 2797 3626 2798 3627
rect 2797 3628 2798 3629
rect 3239 3628 3240 3629
rect 2806 3630 2807 3631
rect 2978 3630 2979 3631
rect 2806 3632 2807 3633
rect 2827 3632 2828 3633
rect 2812 3634 2813 3635
rect 3014 3634 3015 3635
rect 2636 3636 2637 3637
rect 2812 3636 2813 3637
rect 2824 3636 2825 3637
rect 2845 3636 2846 3637
rect 2833 3638 2834 3639
rect 2908 3638 2909 3639
rect 2845 3640 2846 3641
rect 2854 3640 2855 3641
rect 2854 3642 2855 3643
rect 2912 3642 2913 3643
rect 2857 3644 2858 3645
rect 3004 3644 3005 3645
rect 2627 3646 2628 3647
rect 2857 3646 2858 3647
rect 2860 3646 2861 3647
rect 2957 3646 2958 3647
rect 2866 3648 2867 3649
rect 2869 3648 2870 3649
rect 2869 3650 2870 3651
rect 2872 3650 2873 3651
rect 2875 3650 2876 3651
rect 3001 3650 3002 3651
rect 2875 3652 2876 3653
rect 3017 3652 3018 3653
rect 2878 3654 2879 3655
rect 2936 3654 2937 3655
rect 2884 3656 2885 3657
rect 3284 3656 3285 3657
rect 2894 3658 2895 3659
rect 3026 3658 3027 3659
rect 2897 3660 2898 3661
rect 3212 3660 3213 3661
rect 2839 3662 2840 3663
rect 2896 3662 2897 3663
rect 2839 3664 2840 3665
rect 2903 3664 2904 3665
rect 2902 3666 2903 3667
rect 2960 3666 2961 3667
rect 2911 3668 2912 3669
rect 2939 3668 2940 3669
rect 2914 3670 2915 3671
rect 2996 3670 2997 3671
rect 2918 3672 2919 3673
rect 3188 3672 3189 3673
rect 2920 3674 2921 3675
rect 2990 3674 2991 3675
rect 2932 3676 2933 3677
rect 2966 3676 2967 3677
rect 2938 3678 2939 3679
rect 3023 3678 3024 3679
rect 2815 3680 2816 3681
rect 3022 3680 3023 3681
rect 2942 3682 2943 3683
rect 2947 3682 2948 3683
rect 2941 3684 2942 3685
rect 3032 3684 3033 3685
rect 2953 3686 2954 3687
rect 2984 3686 2985 3687
rect 2959 3688 2960 3689
rect 3044 3688 3045 3689
rect 2963 3690 2964 3691
rect 2995 3690 2996 3691
rect 2971 3692 2972 3693
rect 3050 3692 3051 3693
rect 2983 3694 2984 3695
rect 3062 3694 3063 3695
rect 2993 3696 2994 3697
rect 3025 3696 3026 3697
rect 2872 3698 2873 3699
rect 2992 3698 2993 3699
rect 2998 3698 2999 3699
rect 3171 3698 3172 3699
rect 3008 3700 3009 3701
rect 3059 3700 3060 3701
rect 3020 3702 3021 3703
rect 3034 3702 3035 3703
rect 3044 3702 3045 3703
rect 3185 3702 3186 3703
rect 3047 3704 3048 3705
rect 3209 3704 3210 3705
rect 3053 3706 3054 3707
rect 3128 3706 3129 3707
rect 3071 3708 3072 3709
rect 3110 3708 3111 3709
rect 3071 3710 3072 3711
rect 3119 3710 3120 3711
rect 3077 3712 3078 3713
rect 3155 3712 3156 3713
rect 3086 3714 3087 3715
rect 3155 3714 3156 3715
rect 3095 3716 3096 3717
rect 3149 3716 3150 3717
rect 3095 3718 3096 3719
rect 3152 3718 3153 3719
rect 3098 3720 3099 3721
rect 3283 3720 3284 3721
rect 3101 3722 3102 3723
rect 3104 3722 3105 3723
rect 3080 3724 3081 3725
rect 3104 3724 3105 3725
rect 3107 3724 3108 3725
rect 3230 3724 3231 3725
rect 3068 3726 3069 3727
rect 3107 3726 3108 3727
rect 3116 3726 3117 3727
rect 3287 3726 3288 3727
rect 3119 3728 3120 3729
rect 3176 3728 3177 3729
rect 2989 3730 2990 3731
rect 3175 3730 3176 3731
rect 3125 3732 3126 3733
rect 3324 3732 3325 3733
rect 3137 3734 3138 3735
rect 3327 3734 3328 3735
rect 3140 3736 3141 3737
rect 3146 3736 3147 3737
rect 3146 3738 3147 3739
rect 3164 3738 3165 3739
rect 3143 3740 3144 3741
rect 3164 3740 3165 3741
rect 3149 3742 3150 3743
rect 3167 3742 3168 3743
rect 3007 3744 3008 3745
rect 3168 3744 3169 3745
rect 3152 3746 3153 3747
rect 3182 3746 3183 3747
rect 3158 3748 3159 3749
rect 3224 3748 3225 3749
rect 3179 3750 3180 3751
rect 3348 3750 3349 3751
rect 3178 3752 3179 3753
rect 3291 3752 3292 3753
rect 3182 3754 3183 3755
rect 3278 3754 3279 3755
rect 3188 3756 3189 3757
rect 3275 3756 3276 3757
rect 3194 3758 3195 3759
rect 3281 3758 3282 3759
rect 3083 3760 3084 3761
rect 3280 3760 3281 3761
rect 3197 3762 3198 3763
rect 3272 3762 3273 3763
rect 3206 3764 3207 3765
rect 3377 3764 3378 3765
rect 3209 3766 3210 3767
rect 3334 3766 3335 3767
rect 3212 3768 3213 3769
rect 3266 3768 3267 3769
rect 3218 3770 3219 3771
rect 3363 3770 3364 3771
rect 3218 3772 3219 3773
rect 3252 3772 3253 3773
rect 3221 3774 3222 3775
rect 3269 3774 3270 3775
rect 3050 3776 3051 3777
rect 3269 3776 3270 3777
rect 3234 3778 3235 3779
rect 3318 3778 3319 3779
rect 3246 3780 3247 3781
rect 3297 3780 3298 3781
rect 3249 3782 3250 3783
rect 3294 3782 3295 3783
rect 3257 3784 3258 3785
rect 3308 3784 3309 3785
rect 3260 3786 3261 3787
rect 3305 3786 3306 3787
rect 3215 3788 3216 3789
rect 3259 3788 3260 3789
rect 3263 3788 3264 3789
rect 3329 3788 3330 3789
rect 3306 3790 3307 3791
rect 3357 3790 3358 3791
rect 3309 3792 3310 3793
rect 3360 3792 3361 3793
rect 3319 3794 3320 3795
rect 3366 3794 3367 3795
rect 2527 3803 2528 3804
rect 3092 3803 3093 3804
rect 2534 3805 2535 3806
rect 2761 3805 2762 3806
rect 2545 3807 2546 3808
rect 2634 3807 2635 3808
rect 2551 3809 2552 3810
rect 2677 3809 2678 3810
rect 2554 3811 2555 3812
rect 2642 3811 2643 3812
rect 2578 3813 2579 3814
rect 2587 3813 2588 3814
rect 2581 3815 2582 3816
rect 2609 3815 2610 3816
rect 2591 3817 2592 3818
rect 2690 3817 2691 3818
rect 2602 3819 2603 3820
rect 2857 3819 2858 3820
rect 2604 3821 2605 3822
rect 2854 3821 2855 3822
rect 2615 3823 2616 3824
rect 2631 3823 2632 3824
rect 2621 3825 2622 3826
rect 2678 3825 2679 3826
rect 2628 3827 2629 3828
rect 2812 3827 2813 3828
rect 2637 3829 2638 3830
rect 2824 3829 2825 3830
rect 2639 3831 2640 3832
rect 2650 3831 2651 3832
rect 2648 3833 2649 3834
rect 2818 3833 2819 3834
rect 2652 3835 2653 3836
rect 2936 3835 2937 3836
rect 2653 3837 2654 3838
rect 2655 3837 2656 3838
rect 2664 3837 2665 3838
rect 2896 3837 2897 3838
rect 2667 3839 2668 3840
rect 2908 3839 2909 3840
rect 2594 3841 2595 3842
rect 2909 3841 2910 3842
rect 2671 3843 2672 3844
rect 2975 3843 2976 3844
rect 2686 3845 2687 3846
rect 2702 3845 2703 3846
rect 2695 3847 2696 3848
rect 2711 3847 2712 3848
rect 2705 3849 2706 3850
rect 2716 3849 2717 3850
rect 2708 3851 2709 3852
rect 2719 3851 2720 3852
rect 2722 3851 2723 3852
rect 2738 3851 2739 3852
rect 2734 3853 2735 3854
rect 3011 3853 3012 3854
rect 2740 3855 2741 3856
rect 2750 3855 2751 3856
rect 2725 3857 2726 3858
rect 2741 3857 2742 3858
rect 2743 3857 2744 3858
rect 2753 3857 2754 3858
rect 2758 3857 2759 3858
rect 2813 3857 2814 3858
rect 2759 3859 2760 3860
rect 2920 3859 2921 3860
rect 2720 3861 2721 3862
rect 2921 3861 2922 3862
rect 2762 3863 2763 3864
rect 2764 3863 2765 3864
rect 2773 3863 2774 3864
rect 2828 3863 2829 3864
rect 2779 3865 2780 3866
rect 2798 3865 2799 3866
rect 2788 3867 2789 3868
rect 2801 3867 2802 3868
rect 2782 3869 2783 3870
rect 2789 3869 2790 3870
rect 2783 3871 2784 3872
rect 2998 3871 2999 3872
rect 2794 3873 2795 3874
rect 2932 3873 2933 3874
rect 2776 3875 2777 3876
rect 2795 3875 2796 3876
rect 2806 3875 2807 3876
rect 2831 3875 2832 3876
rect 2816 3877 2817 3878
rect 2987 3877 2988 3878
rect 2839 3879 2840 3880
rect 2894 3879 2895 3880
rect 2842 3881 2843 3882
rect 2855 3881 2856 3882
rect 2843 3883 2844 3884
rect 2995 3883 2996 3884
rect 2845 3885 2846 3886
rect 2858 3885 2859 3886
rect 2863 3885 2864 3886
rect 2918 3885 2919 3886
rect 2866 3887 2867 3888
rect 2897 3887 2898 3888
rect 2867 3889 2868 3890
rect 3001 3889 3002 3890
rect 2869 3891 2870 3892
rect 2900 3891 2901 3892
rect 2875 3893 2876 3894
rect 2989 3893 2990 3894
rect 2878 3895 2879 3896
rect 2927 3895 2928 3896
rect 2756 3897 2757 3898
rect 2879 3897 2880 3898
rect 2884 3897 2885 3898
rect 2933 3897 2934 3898
rect 2885 3899 2886 3900
rect 3113 3899 3114 3900
rect 2902 3901 2903 3902
rect 2951 3901 2952 3902
rect 2723 3903 2724 3904
rect 2903 3903 2904 3904
rect 2911 3903 2912 3904
rect 2930 3903 2931 3904
rect 2698 3905 2699 3906
rect 2912 3905 2913 3906
rect 2914 3905 2915 3906
rect 2969 3905 2970 3906
rect 2860 3907 2861 3908
rect 2915 3907 2916 3908
rect 2861 3909 2862 3910
rect 2887 3909 2888 3910
rect 2941 3909 2942 3910
rect 2999 3909 3000 3910
rect 2945 3911 2946 3912
rect 3034 3911 3035 3912
rect 2947 3913 2948 3914
rect 2957 3913 2958 3914
rect 2953 3915 2954 3916
rect 2981 3915 2982 3916
rect 2954 3917 2955 3918
rect 3161 3917 3162 3918
rect 2959 3919 2960 3920
rect 3125 3919 3126 3920
rect 2971 3921 2972 3922
rect 3017 3921 3018 3922
rect 2972 3923 2973 3924
rect 3004 3923 3005 3924
rect 2978 3925 2979 3926
rect 3025 3925 3026 3926
rect 3005 3927 3006 3928
rect 3044 3927 3045 3928
rect 3029 3929 3030 3930
rect 3107 3929 3108 3930
rect 3032 3931 3033 3932
rect 3110 3931 3111 3932
rect 3041 3933 3042 3934
rect 3059 3933 3060 3934
rect 3041 3935 3042 3936
rect 3143 3935 3144 3936
rect 2770 3937 2771 3938
rect 3143 3937 3144 3938
rect 2771 3939 2772 3940
rect 3309 3939 3310 3940
rect 3050 3941 3051 3942
rect 3086 3941 3087 3942
rect 3062 3943 3063 3944
rect 3241 3943 3242 3944
rect 3071 3945 3072 3946
rect 3113 3945 3114 3946
rect 3074 3947 3075 3948
rect 3140 3947 3141 3948
rect 3077 3949 3078 3950
rect 3140 3949 3141 3950
rect 3044 3951 3045 3952
rect 3077 3951 3078 3952
rect 3080 3951 3081 3952
rect 3101 3951 3102 3952
rect 3095 3953 3096 3954
rect 3280 3953 3281 3954
rect 3098 3955 3099 3956
rect 3280 3955 3281 3956
rect 3098 3957 3099 3958
rect 3146 3957 3147 3958
rect 3047 3959 3048 3960
rect 3146 3959 3147 3960
rect 3122 3961 3123 3962
rect 3155 3961 3156 3962
rect 3137 3963 3138 3964
rect 3262 3963 3263 3964
rect 3083 3965 3084 3966
rect 3137 3965 3138 3966
rect 3083 3967 3084 3968
rect 3104 3967 3105 3968
rect 3149 3967 3150 3968
rect 3164 3967 3165 3968
rect 3155 3969 3156 3970
rect 3259 3969 3260 3970
rect 3068 3971 3069 3972
rect 3259 3971 3260 3972
rect 3164 3973 3165 3974
rect 3262 3973 3263 3974
rect 3168 3975 3169 3976
rect 3256 3975 3257 3976
rect 3191 3977 3192 3978
rect 3197 3977 3198 3978
rect 3194 3979 3195 3980
rect 3224 3979 3225 3980
rect 3188 3981 3189 3982
rect 3194 3981 3195 3982
rect 3197 3981 3198 3982
rect 3315 3981 3316 3982
rect 3206 3983 3207 3984
rect 3218 3983 3219 3984
rect 3212 3985 3213 3986
rect 3218 3985 3219 3986
rect 3209 3987 3210 3988
rect 3212 3987 3213 3988
rect 3158 3989 3159 3990
rect 3209 3989 3210 3990
rect 2938 3991 2939 3992
rect 3158 3991 3159 3992
rect 2939 3993 2940 3994
rect 3022 3993 3023 3994
rect 2983 3995 2984 3996
rect 3023 3995 3024 3996
rect 2984 3997 2985 3998
rect 2992 3997 2993 3998
rect 3215 3997 3216 3998
rect 3252 3997 3253 3998
rect 3215 3999 3216 4000
rect 3266 3999 3267 4000
rect 3221 4001 3222 4002
rect 3287 4001 3288 4002
rect 3119 4003 3120 4004
rect 3287 4003 3288 4004
rect 3119 4005 3120 4006
rect 3152 4005 3153 4006
rect 3234 4005 3235 4006
rect 3302 4005 3303 4006
rect 3246 4007 3247 4008
rect 3253 4007 3254 4008
rect 3249 4009 3250 4010
rect 3319 4009 3320 4010
rect 3293 4011 3294 4012
rect 3306 4011 3307 4012
rect 3053 4013 3054 4014
rect 3306 4013 3307 4014
rect 3007 4015 3008 4016
rect 3053 4015 3054 4016
rect 3296 4015 3297 4016
rect 3322 4015 3323 4016
rect 2555 4024 2556 4025
rect 2570 4024 2571 4025
rect 2567 4026 2568 4027
rect 2634 4026 2635 4027
rect 2576 4028 2577 4029
rect 2851 4028 2852 4029
rect 2579 4030 2580 4031
rect 2586 4030 2587 4031
rect 2588 4030 2589 4031
rect 2595 4030 2596 4031
rect 2589 4032 2590 4033
rect 2690 4032 2691 4033
rect 2593 4034 2594 4035
rect 2891 4034 2892 4035
rect 2581 4036 2582 4037
rect 2890 4036 2891 4037
rect 2603 4038 2604 4039
rect 2801 4038 2802 4039
rect 2612 4040 2613 4041
rect 2672 4040 2673 4041
rect 2619 4042 2620 4043
rect 2944 4042 2945 4043
rect 2622 4044 2623 4045
rect 2831 4044 2832 4045
rect 2624 4046 2625 4047
rect 2741 4046 2742 4047
rect 2626 4048 2627 4049
rect 2734 4048 2735 4049
rect 2640 4050 2641 4051
rect 2912 4050 2913 4051
rect 2636 4052 2637 4053
rect 2911 4052 2912 4053
rect 2644 4054 2645 4055
rect 2984 4054 2985 4055
rect 2653 4056 2654 4057
rect 2708 4056 2709 4057
rect 2678 4058 2679 4059
rect 2830 4058 2831 4059
rect 2688 4060 2689 4061
rect 2791 4060 2792 4061
rect 2697 4062 2698 4063
rect 2705 4062 2706 4063
rect 2700 4064 2701 4065
rect 2711 4064 2712 4065
rect 2720 4064 2721 4065
rect 2959 4064 2960 4065
rect 2722 4066 2723 4067
rect 3007 4066 3008 4067
rect 2728 4068 2729 4069
rect 2738 4068 2739 4069
rect 2740 4068 2741 4069
rect 2750 4068 2751 4069
rect 2743 4070 2744 4071
rect 2753 4070 2754 4071
rect 2746 4072 2747 4073
rect 2762 4072 2763 4073
rect 2749 4074 2750 4075
rect 2867 4074 2868 4075
rect 2759 4076 2760 4077
rect 3293 4076 3294 4077
rect 2767 4078 2768 4079
rect 2954 4078 2955 4079
rect 2771 4080 2772 4081
rect 2981 4080 2982 4081
rect 2773 4082 2774 4083
rect 2783 4082 2784 4083
rect 2785 4082 2786 4083
rect 2795 4082 2796 4083
rect 2806 4082 2807 4083
rect 2816 4082 2817 4083
rect 2818 4082 2819 4083
rect 2828 4082 2829 4083
rect 2605 4084 2606 4085
rect 2827 4084 2828 4085
rect 2839 4084 2840 4085
rect 2855 4084 2856 4085
rect 2843 4086 2844 4087
rect 3184 4086 3185 4087
rect 2842 4088 2843 4089
rect 2858 4088 2859 4089
rect 2845 4090 2846 4091
rect 2861 4090 2862 4091
rect 2854 4092 2855 4093
rect 2939 4092 2940 4093
rect 2860 4094 2861 4095
rect 2918 4094 2919 4095
rect 2789 4096 2790 4097
rect 2917 4096 2918 4097
rect 2788 4098 2789 4099
rect 2798 4098 2799 4099
rect 2797 4100 2798 4101
rect 2813 4100 2814 4101
rect 2812 4102 2813 4103
rect 2837 4102 2838 4103
rect 2866 4102 2867 4103
rect 2879 4102 2880 4103
rect 2596 4104 2597 4105
rect 2878 4104 2879 4105
rect 2872 4106 2873 4107
rect 2885 4106 2886 4107
rect 2584 4108 2585 4109
rect 2884 4108 2885 4109
rect 2881 4110 2882 4111
rect 2894 4110 2895 4111
rect 2702 4112 2703 4113
rect 2893 4112 2894 4113
rect 2921 4112 2922 4113
rect 2938 4112 2939 4113
rect 2678 4114 2679 4115
rect 2920 4114 2921 4115
rect 2965 4114 2966 4115
rect 2992 4114 2993 4115
rect 2975 4116 2976 4117
rect 2980 4116 2981 4117
rect 2969 4118 2970 4119
rect 2974 4118 2975 4119
rect 2957 4120 2958 4121
rect 2968 4120 2969 4121
rect 2951 4122 2952 4123
rect 2956 4122 2957 4123
rect 2978 4122 2979 4123
rect 2983 4122 2984 4123
rect 2972 4124 2973 4125
rect 2977 4124 2978 4125
rect 2987 4124 2988 4125
rect 3032 4124 3033 4125
rect 2948 4126 2949 4127
rect 2986 4126 2987 4127
rect 2936 4128 2937 4129
rect 2947 4128 2948 4129
rect 2990 4128 2991 4129
rect 3029 4128 3030 4129
rect 2999 4130 3000 4131
rect 3001 4130 3002 4131
rect 3005 4130 3006 4131
rect 3040 4130 3041 4131
rect 3017 4132 3018 4133
rect 3019 4132 3020 4133
rect 3023 4132 3024 4133
rect 3058 4132 3059 4133
rect 3025 4134 3026 4135
rect 3181 4134 3182 4135
rect 3037 4136 3038 4137
rect 3125 4136 3126 4137
rect 3049 4138 3050 4139
rect 3098 4138 3099 4139
rect 3053 4140 3054 4141
rect 3130 4140 3131 4141
rect 3052 4142 3053 4143
rect 3157 4142 3158 4143
rect 3055 4144 3056 4145
rect 3119 4144 3120 4145
rect 3074 4146 3075 4147
rect 3332 4146 3333 4147
rect 3068 4148 3069 4149
rect 3073 4148 3074 4149
rect 3062 4150 3063 4151
rect 3067 4150 3068 4151
rect 3061 4152 3062 4153
rect 3083 4152 3084 4153
rect 3080 4154 3081 4155
rect 3103 4154 3104 4155
rect 3086 4156 3087 4157
rect 3109 4156 3110 4157
rect 3092 4158 3093 4159
rect 3227 4158 3228 4159
rect 3106 4160 3107 4161
rect 3167 4160 3168 4161
rect 3113 4162 3114 4163
rect 3203 4162 3204 4163
rect 3115 4164 3116 4165
rect 3152 4164 3153 4165
rect 3118 4166 3119 4167
rect 3188 4166 3189 4167
rect 3122 4168 3123 4169
rect 3241 4168 3242 4169
rect 3137 4170 3138 4171
rect 3302 4170 3303 4171
rect 3146 4172 3147 4173
rect 3166 4172 3167 4173
rect 3155 4174 3156 4175
rect 3260 4174 3261 4175
rect 3164 4176 3165 4177
rect 3320 4176 3321 4177
rect 3143 4178 3144 4179
rect 3163 4178 3164 4179
rect 3169 4178 3170 4179
rect 3285 4178 3286 4179
rect 3194 4180 3195 4181
rect 3200 4180 3201 4181
rect 3194 4182 3195 4183
rect 3276 4182 3277 4183
rect 3209 4184 3210 4185
rect 3236 4184 3237 4185
rect 2715 4186 2716 4187
rect 3209 4186 3210 4187
rect 3212 4186 3213 4187
rect 3248 4186 3249 4187
rect 3212 4188 3213 4189
rect 3215 4188 3216 4189
rect 3218 4188 3219 4189
rect 3251 4188 3252 4189
rect 3221 4190 3222 4191
rect 3269 4190 3270 4191
rect 3127 4192 3128 4193
rect 3221 4192 3222 4193
rect 3224 4192 3225 4193
rect 3230 4192 3231 4193
rect 3197 4194 3198 4195
rect 3224 4194 3225 4195
rect 3140 4196 3141 4197
rect 3197 4196 3198 4197
rect 3077 4198 3078 4199
rect 3139 4198 3140 4199
rect 3233 4198 3234 4199
rect 3309 4198 3310 4199
rect 3244 4200 3245 4201
rect 3253 4200 3254 4201
rect 3254 4202 3255 4203
rect 3316 4202 3317 4203
rect 3245 4204 3246 4205
rect 3316 4204 3317 4205
rect 3256 4206 3257 4207
rect 3306 4206 3307 4207
rect 3191 4208 3192 4209
rect 3257 4208 3258 4209
rect 3290 4208 3291 4209
rect 3313 4208 3314 4209
rect 3296 4210 3297 4211
rect 3299 4210 3300 4211
rect 2557 4219 2558 4220
rect 2570 4219 2571 4220
rect 2560 4221 2561 4222
rect 2564 4221 2565 4222
rect 2567 4221 2568 4222
rect 2576 4221 2577 4222
rect 2582 4221 2583 4222
rect 2730 4221 2731 4222
rect 2586 4223 2587 4224
rect 2706 4223 2707 4224
rect 2594 4225 2595 4226
rect 2881 4225 2882 4226
rect 2600 4227 2601 4228
rect 2917 4227 2918 4228
rect 2612 4229 2613 4230
rect 2682 4229 2683 4230
rect 2619 4231 2620 4232
rect 2890 4231 2891 4232
rect 2622 4233 2623 4234
rect 2851 4233 2852 4234
rect 2622 4235 2623 4236
rect 2860 4235 2861 4236
rect 2626 4237 2627 4238
rect 2715 4237 2716 4238
rect 2633 4239 2634 4240
rect 2920 4239 2921 4240
rect 2632 4241 2633 4242
rect 2947 4241 2948 4242
rect 2636 4243 2637 4244
rect 2734 4243 2735 4244
rect 2636 4245 2637 4246
rect 2740 4245 2741 4246
rect 2639 4247 2640 4248
rect 3013 4247 3014 4248
rect 2643 4249 2644 4250
rect 2971 4249 2972 4250
rect 2646 4251 2647 4252
rect 2821 4251 2822 4252
rect 2648 4253 2649 4254
rect 2845 4253 2846 4254
rect 2651 4255 2652 4256
rect 2667 4255 2668 4256
rect 2672 4255 2673 4256
rect 2688 4255 2689 4256
rect 2673 4257 2674 4258
rect 2718 4257 2719 4258
rect 2694 4259 2695 4260
rect 2851 4259 2852 4260
rect 2697 4261 2698 4262
rect 2848 4261 2849 4262
rect 2709 4263 2710 4264
rect 2743 4263 2744 4264
rect 2728 4265 2729 4266
rect 2764 4265 2765 4266
rect 2746 4267 2747 4268
rect 2800 4267 2801 4268
rect 2746 4269 2747 4270
rect 3118 4269 3119 4270
rect 2749 4271 2750 4272
rect 2995 4271 2996 4272
rect 2700 4273 2701 4274
rect 2749 4273 2750 4274
rect 2752 4273 2753 4274
rect 2992 4273 2993 4274
rect 2603 4275 2604 4276
rect 2992 4275 2993 4276
rect 2604 4277 2605 4278
rect 2608 4277 2609 4278
rect 2767 4277 2768 4278
rect 2776 4277 2777 4278
rect 2797 4277 2798 4278
rect 2857 4277 2858 4278
rect 2803 4279 2804 4280
rect 2806 4279 2807 4280
rect 2812 4279 2813 4280
rect 2860 4279 2861 4280
rect 2812 4281 2813 4282
rect 2905 4281 2906 4282
rect 2815 4283 2816 4284
rect 2854 4283 2855 4284
rect 2830 4285 2831 4286
rect 2869 4285 2870 4286
rect 2788 4287 2789 4288
rect 2830 4287 2831 4288
rect 2773 4289 2774 4290
rect 2788 4289 2789 4290
rect 2845 4289 2846 4290
rect 2965 4289 2966 4290
rect 2743 4291 2744 4292
rect 2965 4291 2966 4292
rect 2872 4293 2873 4294
rect 3016 4293 3017 4294
rect 2818 4295 2819 4296
rect 2872 4295 2873 4296
rect 2887 4295 2888 4296
rect 2902 4295 2903 4296
rect 2893 4297 2894 4298
rect 2962 4297 2963 4298
rect 2839 4299 2840 4300
rect 2893 4299 2894 4300
rect 2791 4301 2792 4302
rect 2839 4301 2840 4302
rect 2899 4301 2900 4302
rect 2917 4301 2918 4302
rect 2899 4303 2900 4304
rect 2938 4303 2939 4304
rect 2908 4305 2909 4306
rect 2947 4305 2948 4306
rect 2866 4307 2867 4308
rect 2908 4307 2909 4308
rect 2827 4309 2828 4310
rect 2866 4309 2867 4310
rect 2785 4311 2786 4312
rect 2827 4311 2828 4312
rect 2914 4311 2915 4312
rect 2989 4311 2990 4312
rect 2896 4313 2897 4314
rect 2914 4313 2915 4314
rect 2926 4313 2927 4314
rect 2953 4313 2954 4314
rect 2941 4315 2942 4316
rect 2968 4315 2969 4316
rect 2950 4317 2951 4318
rect 2998 4317 2999 4318
rect 2911 4319 2912 4320
rect 2950 4319 2951 4320
rect 2956 4319 2957 4320
rect 3300 4319 3301 4320
rect 2929 4321 2930 4322
rect 2956 4321 2957 4322
rect 2794 4323 2795 4324
rect 2929 4323 2930 4324
rect 2959 4323 2960 4324
rect 2986 4323 2987 4324
rect 2884 4325 2885 4326
rect 2959 4325 2960 4326
rect 2980 4325 2981 4326
rect 3031 4325 3032 4326
rect 2983 4327 2984 4328
rect 3034 4327 3035 4328
rect 2727 4329 2728 4330
rect 2983 4329 2984 4330
rect 3001 4329 3002 4330
rect 3076 4329 3077 4330
rect 2944 4331 2945 4332
rect 3001 4331 3002 4332
rect 3010 4331 3011 4332
rect 3022 4331 3023 4332
rect 3019 4333 3020 4334
rect 3082 4333 3083 4334
rect 3007 4335 3008 4336
rect 3019 4335 3020 4336
rect 3025 4335 3026 4336
rect 3088 4335 3089 4336
rect 3037 4337 3038 4338
rect 3079 4337 3080 4338
rect 3040 4339 3041 4340
rect 3139 4339 3140 4340
rect 3043 4341 3044 4342
rect 3157 4341 3158 4342
rect 3055 4343 3056 4344
rect 3091 4343 3092 4344
rect 3052 4345 3053 4346
rect 3055 4345 3056 4346
rect 2977 4347 2978 4348
rect 3052 4347 3053 4348
rect 2932 4349 2933 4350
rect 2977 4349 2978 4350
rect 2878 4351 2879 4352
rect 2932 4351 2933 4352
rect 3058 4351 3059 4352
rect 3184 4351 3185 4352
rect 3049 4353 3050 4354
rect 3058 4353 3059 4354
rect 2974 4355 2975 4356
rect 3049 4355 3050 4356
rect 2842 4357 2843 4358
rect 2974 4357 2975 4358
rect 3061 4357 3062 4358
rect 3094 4357 3095 4358
rect 3067 4359 3068 4360
rect 3139 4359 3140 4360
rect 3064 4361 3065 4362
rect 3067 4361 3068 4362
rect 3073 4361 3074 4362
rect 3278 4361 3279 4362
rect 3073 4363 3074 4364
rect 3115 4363 3116 4364
rect 3103 4365 3104 4366
rect 3121 4365 3122 4366
rect 3106 4367 3107 4368
rect 3124 4367 3125 4368
rect 3106 4369 3107 4370
rect 3206 4369 3207 4370
rect 3109 4371 3110 4372
rect 3157 4371 3158 4372
rect 3118 4373 3119 4374
rect 3257 4373 3258 4374
rect 3127 4375 3128 4376
rect 3184 4375 3185 4376
rect 3127 4377 3128 4378
rect 3267 4377 3268 4378
rect 3133 4379 3134 4380
rect 3281 4379 3282 4380
rect 3166 4381 3167 4382
rect 3205 4381 3206 4382
rect 3169 4383 3170 4384
rect 3326 4383 3327 4384
rect 3181 4385 3182 4386
rect 3221 4385 3222 4386
rect 3212 4387 3213 4388
rect 3218 4387 3219 4388
rect 2809 4389 2810 4390
rect 3217 4389 3218 4390
rect 3224 4389 3225 4390
rect 3260 4389 3261 4390
rect 3227 4391 3228 4392
rect 3263 4391 3264 4392
rect 3200 4393 3201 4394
rect 3226 4393 3227 4394
rect 3230 4393 3231 4394
rect 3266 4393 3267 4394
rect 3203 4395 3204 4396
rect 3229 4395 3230 4396
rect 3163 4397 3164 4398
rect 3202 4397 3203 4398
rect 3233 4397 3234 4398
rect 3269 4397 3270 4398
rect 3194 4399 3195 4400
rect 3232 4399 3233 4400
rect 3193 4401 3194 4402
rect 3370 4401 3371 4402
rect 3236 4403 3237 4404
rect 3291 4403 3292 4404
rect 3197 4405 3198 4406
rect 3235 4405 3236 4406
rect 3248 4405 3249 4406
rect 3315 4405 3316 4406
rect 3112 4407 3113 4408
rect 3248 4407 3249 4408
rect 3254 4407 3255 4408
rect 3306 4407 3307 4408
rect 3191 4409 3192 4410
rect 3254 4409 3255 4410
rect 3294 4409 3295 4410
rect 3329 4409 3330 4410
rect 3302 4411 3303 4412
rect 3319 4411 3320 4412
rect 3251 4413 3252 4414
rect 3303 4413 3304 4414
rect 3245 4415 3246 4416
rect 3251 4415 3252 4416
rect 3130 4417 3131 4418
rect 3245 4417 3246 4418
rect 3309 4417 3310 4418
rect 3347 4417 3348 4418
rect 3309 4419 3310 4420
rect 3343 4419 3344 4420
rect 3356 4419 3357 4420
rect 3367 4419 3368 4420
rect 2539 4428 2540 4429
rect 2749 4428 2750 4429
rect 2588 4430 2589 4431
rect 2899 4430 2900 4431
rect 2590 4432 2591 4433
rect 2959 4432 2960 4433
rect 2602 4434 2603 4435
rect 2778 4434 2779 4435
rect 2611 4436 2612 4437
rect 2615 4436 2616 4437
rect 2612 4438 2613 4439
rect 2947 4438 2948 4439
rect 2622 4440 2623 4441
rect 2682 4440 2683 4441
rect 2632 4442 2633 4443
rect 2908 4442 2909 4443
rect 2594 4444 2595 4445
rect 2907 4444 2908 4445
rect 2595 4446 2596 4447
rect 2706 4446 2707 4447
rect 2636 4448 2637 4449
rect 2925 4448 2926 4449
rect 2638 4450 2639 4451
rect 2953 4450 2954 4451
rect 2643 4452 2644 4453
rect 2860 4452 2861 4453
rect 2649 4454 2650 4455
rect 3052 4454 3053 4455
rect 2656 4456 2657 4457
rect 2835 4456 2836 4457
rect 2659 4458 2660 4459
rect 2848 4458 2849 4459
rect 2662 4460 2663 4461
rect 2667 4460 2668 4461
rect 2665 4462 2666 4463
rect 2709 4462 2710 4463
rect 2680 4464 2681 4465
rect 2983 4464 2984 4465
rect 2686 4466 2687 4467
rect 2950 4466 2951 4467
rect 2697 4468 2698 4469
rect 2821 4468 2822 4469
rect 2707 4470 2708 4471
rect 2730 4470 2731 4471
rect 2710 4472 2711 4473
rect 2962 4472 2963 4473
rect 2728 4474 2729 4475
rect 2735 4474 2736 4475
rect 2739 4474 2740 4475
rect 2941 4474 2942 4475
rect 2739 4476 2740 4477
rect 2998 4476 2999 4477
rect 2757 4478 2758 4479
rect 2800 4478 2801 4479
rect 2766 4480 2767 4481
rect 2776 4480 2777 4481
rect 2784 4480 2785 4481
rect 2827 4480 2828 4481
rect 2788 4482 2789 4483
rect 2790 4482 2791 4483
rect 2787 4484 2788 4485
rect 2830 4484 2831 4485
rect 2794 4486 2795 4487
rect 2805 4486 2806 4487
rect 2796 4488 2797 4489
rect 2857 4488 2858 4489
rect 2799 4490 2800 4491
rect 2992 4490 2993 4491
rect 2812 4492 2813 4493
rect 2889 4492 2890 4493
rect 2803 4494 2804 4495
rect 2811 4494 2812 4495
rect 2817 4494 2818 4495
rect 2872 4494 2873 4495
rect 2820 4496 2821 4497
rect 2839 4496 2840 4497
rect 2823 4498 2824 4499
rect 2956 4498 2957 4499
rect 2618 4500 2619 4501
rect 2955 4500 2956 4501
rect 2619 4502 2620 4503
rect 2764 4502 2765 4503
rect 2826 4502 2827 4503
rect 2866 4502 2867 4503
rect 2832 4504 2833 4505
rect 2845 4504 2846 4505
rect 2815 4506 2816 4507
rect 2844 4506 2845 4507
rect 2838 4508 2839 4509
rect 2851 4508 2852 4509
rect 2850 4510 2851 4511
rect 2893 4510 2894 4511
rect 2609 4512 2610 4513
rect 2892 4512 2893 4513
rect 2862 4514 2863 4515
rect 2887 4514 2888 4515
rect 2869 4516 2870 4517
rect 2895 4516 2896 4517
rect 2629 4518 2630 4519
rect 2868 4518 2869 4519
rect 2628 4520 2629 4521
rect 2688 4520 2689 4521
rect 2689 4522 2690 4523
rect 2914 4522 2915 4523
rect 2871 4524 2872 4525
rect 2917 4524 2918 4525
rect 2874 4526 2875 4527
rect 2932 4526 2933 4527
rect 2886 4528 2887 4529
rect 2905 4528 2906 4529
rect 2598 4530 2599 4531
rect 2904 4530 2905 4531
rect 2910 4530 2911 4531
rect 2977 4530 2978 4531
rect 2916 4532 2917 4533
rect 2971 4532 2972 4533
rect 2919 4534 2920 4535
rect 2974 4534 2975 4535
rect 2922 4536 2923 4537
rect 2989 4536 2990 4537
rect 2646 4538 2647 4539
rect 2988 4538 2989 4539
rect 2645 4540 2646 4541
rect 2934 4540 2935 4541
rect 2929 4542 2930 4543
rect 3129 4542 3130 4543
rect 2940 4544 2941 4545
rect 2995 4544 2996 4545
rect 2943 4546 2944 4547
rect 3001 4546 3002 4547
rect 2949 4548 2950 4549
rect 3013 4548 3014 4549
rect 2958 4550 2959 4551
rect 3016 4550 3017 4551
rect 2961 4552 2962 4553
rect 2965 4552 2966 4553
rect 2964 4554 2965 4555
rect 2986 4554 2987 4555
rect 2979 4556 2980 4557
rect 3031 4556 3032 4557
rect 2982 4558 2983 4559
rect 3034 4558 3035 4559
rect 2985 4560 2986 4561
rect 3049 4560 3050 4561
rect 2991 4562 2992 4563
rect 3019 4562 3020 4563
rect 2994 4564 2995 4565
rect 3022 4564 3023 4565
rect 3015 4566 3016 4567
rect 3076 4566 3077 4567
rect 3021 4568 3022 4569
rect 3067 4568 3068 4569
rect 3024 4570 3025 4571
rect 3079 4570 3080 4571
rect 3027 4572 3028 4573
rect 3055 4572 3056 4573
rect 3030 4574 3031 4575
rect 3043 4574 3044 4575
rect 3033 4576 3034 4577
rect 3082 4576 3083 4577
rect 3039 4578 3040 4579
rect 3088 4578 3089 4579
rect 3042 4580 3043 4581
rect 3091 4580 3092 4581
rect 3048 4582 3049 4583
rect 3121 4582 3122 4583
rect 3058 4584 3059 4585
rect 3241 4584 3242 4585
rect 3073 4586 3074 4587
rect 3141 4586 3142 4587
rect 3081 4588 3082 4589
rect 3214 4588 3215 4589
rect 3087 4590 3088 4591
rect 3124 4590 3125 4591
rect 3090 4592 3091 4593
rect 3094 4592 3095 4593
rect 3099 4592 3100 4593
rect 3127 4592 3128 4593
rect 3106 4594 3107 4595
rect 3245 4594 3246 4595
rect 3112 4596 3113 4597
rect 3150 4596 3151 4597
rect 3111 4598 3112 4599
rect 3282 4598 3283 4599
rect 3114 4600 3115 4601
rect 3244 4600 3245 4601
rect 3118 4602 3119 4603
rect 3120 4602 3121 4603
rect 3117 4604 3118 4605
rect 3254 4604 3255 4605
rect 3123 4606 3124 4607
rect 3263 4606 3264 4607
rect 3133 4608 3134 4609
rect 3256 4608 3257 4609
rect 3139 4610 3140 4611
rect 3271 4610 3272 4611
rect 3147 4612 3148 4613
rect 3181 4612 3182 4613
rect 3157 4614 3158 4615
rect 3241 4614 3242 4615
rect 3177 4616 3178 4617
rect 3235 4616 3236 4617
rect 3051 4618 3052 4619
rect 3235 4618 3236 4619
rect 3184 4620 3185 4621
rect 3187 4620 3188 4621
rect 3193 4620 3194 4621
rect 3363 4620 3364 4621
rect 3144 4622 3145 4623
rect 3192 4622 3193 4623
rect 3195 4622 3196 4623
rect 3202 4622 3203 4623
rect 3198 4624 3199 4625
rect 3205 4624 3206 4625
rect 3204 4626 3205 4627
rect 3238 4626 3239 4627
rect 3207 4628 3208 4629
rect 3269 4628 3270 4629
rect 3093 4630 3094 4631
rect 3268 4630 3269 4631
rect 3210 4632 3211 4633
rect 3226 4632 3227 4633
rect 3213 4634 3214 4635
rect 3229 4634 3230 4635
rect 3216 4636 3217 4637
rect 3232 4636 3233 4637
rect 3219 4638 3220 4639
rect 3321 4638 3322 4639
rect 3222 4640 3223 4641
rect 3329 4640 3330 4641
rect 3238 4642 3239 4643
rect 3312 4642 3313 4643
rect 3251 4644 3252 4645
rect 3315 4644 3316 4645
rect 3260 4646 3261 4647
rect 3262 4646 3263 4647
rect 3259 4648 3260 4649
rect 3340 4648 3341 4649
rect 3266 4650 3267 4651
rect 3314 4650 3315 4651
rect 3265 4652 3266 4653
rect 3291 4652 3292 4653
rect 3274 4654 3275 4655
rect 3303 4654 3304 4655
rect 3277 4656 3278 4657
rect 3347 4656 3348 4657
rect 3279 4658 3280 4659
rect 3283 4658 3284 4659
rect 3280 4660 3281 4661
rect 3309 4660 3310 4661
rect 3286 4662 3287 4663
rect 3306 4662 3307 4663
rect 3294 4664 3295 4665
rect 3337 4664 3338 4665
rect 2575 4673 2576 4674
rect 2784 4673 2785 4674
rect 2581 4675 2582 4676
rect 2707 4675 2708 4676
rect 2582 4677 2583 4678
rect 2778 4677 2779 4678
rect 2588 4679 2589 4680
rect 2874 4679 2875 4680
rect 2599 4681 2600 4682
rect 2750 4681 2751 4682
rect 2605 4683 2606 4684
rect 2925 4683 2926 4684
rect 2609 4685 2610 4686
rect 2799 4685 2800 4686
rect 2613 4687 2614 4688
rect 2686 4687 2687 4688
rect 2635 4689 2636 4690
rect 2873 4689 2874 4690
rect 2628 4691 2629 4692
rect 2635 4691 2636 4692
rect 2642 4691 2643 4692
rect 2868 4691 2869 4692
rect 2645 4693 2646 4694
rect 2783 4693 2784 4694
rect 2649 4695 2650 4696
rect 2820 4695 2821 4696
rect 2652 4697 2653 4698
rect 2949 4697 2950 4698
rect 2655 4699 2656 4700
rect 2662 4699 2663 4700
rect 2667 4699 2668 4700
rect 2895 4699 2896 4700
rect 2680 4701 2681 4702
rect 2961 4701 2962 4702
rect 2679 4703 2680 4704
rect 2683 4703 2684 4704
rect 2686 4703 2687 4704
rect 2698 4703 2699 4704
rect 2692 4705 2693 4706
rect 2985 4705 2986 4706
rect 2692 4707 2693 4708
rect 2710 4707 2711 4708
rect 2707 4709 2708 4710
rect 2787 4709 2788 4710
rect 2710 4711 2711 4712
rect 2757 4711 2758 4712
rect 2713 4713 2714 4714
rect 2982 4713 2983 4714
rect 2723 4715 2724 4716
rect 2940 4715 2941 4716
rect 2725 4717 2726 4718
rect 2979 4717 2980 4718
rect 2616 4719 2617 4720
rect 2726 4719 2727 4720
rect 2617 4721 2618 4722
rect 2892 4721 2893 4722
rect 2735 4723 2736 4724
rect 3125 4723 3126 4724
rect 2739 4725 2740 4726
rect 2898 4725 2899 4726
rect 2747 4727 2748 4728
rect 2817 4727 2818 4728
rect 2766 4729 2767 4730
rect 2768 4729 2769 4730
rect 2774 4729 2775 4730
rect 2790 4729 2791 4730
rect 2780 4731 2781 4732
rect 2826 4731 2827 4732
rect 2792 4733 2793 4734
rect 2832 4733 2833 4734
rect 2798 4735 2799 4736
rect 2838 4735 2839 4736
rect 2805 4737 2806 4738
rect 2819 4737 2820 4738
rect 2804 4739 2805 4740
rect 2850 4739 2851 4740
rect 2816 4741 2817 4742
rect 2844 4741 2845 4742
rect 2649 4743 2650 4744
rect 2843 4743 2844 4744
rect 2823 4745 2824 4746
rect 3310 4745 3311 4746
rect 2828 4747 2829 4748
rect 2904 4747 2905 4748
rect 2661 4749 2662 4750
rect 2903 4749 2904 4750
rect 2831 4751 2832 4752
rect 2907 4751 2908 4752
rect 2837 4753 2838 4754
rect 2964 4753 2965 4754
rect 2840 4755 2841 4756
rect 2922 4755 2923 4756
rect 2849 4757 2850 4758
rect 2916 4757 2917 4758
rect 2732 4759 2733 4760
rect 2915 4759 2916 4760
rect 2732 4761 2733 4762
rect 2796 4761 2797 4762
rect 2795 4763 2796 4764
rect 2835 4763 2836 4764
rect 2834 4765 2835 4766
rect 2862 4765 2863 4766
rect 2852 4767 2853 4768
rect 2919 4767 2920 4768
rect 2855 4769 2856 4770
rect 2910 4769 2911 4770
rect 2861 4771 2862 4772
rect 2934 4771 2935 4772
rect 2867 4773 2868 4774
rect 2943 4773 2944 4774
rect 2871 4775 2872 4776
rect 2876 4775 2877 4776
rect 2879 4775 2880 4776
rect 2955 4775 2956 4776
rect 2882 4777 2883 4778
rect 2958 4777 2959 4778
rect 2886 4779 2887 4780
rect 2891 4779 2892 4780
rect 2889 4781 2890 4782
rect 2918 4781 2919 4782
rect 2897 4783 2898 4784
rect 2951 4783 2952 4784
rect 2901 4785 2902 4786
rect 2966 4785 2967 4786
rect 2909 4787 2910 4788
rect 2988 4787 2989 4788
rect 2912 4789 2913 4790
rect 3068 4789 3069 4790
rect 2927 4791 2928 4792
rect 2994 4791 2995 4792
rect 2930 4793 2931 4794
rect 2991 4793 2992 4794
rect 2933 4795 2934 4796
rect 3015 4795 3016 4796
rect 2939 4797 2940 4798
rect 3021 4797 3022 4798
rect 2957 4799 2958 4800
rect 3033 4799 3034 4800
rect 2728 4801 2729 4802
rect 3032 4801 3033 4802
rect 2963 4803 2964 4804
rect 3024 4803 3025 4804
rect 2969 4805 2970 4806
rect 3039 4805 3040 4806
rect 2975 4807 2976 4808
rect 3120 4807 3121 4808
rect 2978 4809 2979 4810
rect 3045 4809 3046 4810
rect 2990 4811 2991 4812
rect 3027 4811 3028 4812
rect 2996 4813 2997 4814
rect 3081 4813 3082 4814
rect 3002 4815 3003 4816
rect 3165 4815 3166 4816
rect 3014 4817 3015 4818
rect 3099 4817 3100 4818
rect 3030 4819 3031 4820
rect 3035 4819 3036 4820
rect 3038 4819 3039 4820
rect 3111 4819 3112 4820
rect 3042 4821 3043 4822
rect 3080 4821 3081 4822
rect 3041 4823 3042 4824
rect 3123 4823 3124 4824
rect 3047 4825 3048 4826
rect 3051 4825 3052 4826
rect 3065 4825 3066 4826
rect 3087 4825 3088 4826
rect 3083 4827 3084 4828
rect 3131 4827 3132 4828
rect 3098 4829 3099 4830
rect 3147 4829 3148 4830
rect 3101 4831 3102 4832
rect 3150 4831 3151 4832
rect 3104 4833 3105 4834
rect 3195 4833 3196 4834
rect 3090 4835 3091 4836
rect 3194 4835 3195 4836
rect 3107 4837 3108 4838
rect 3198 4837 3199 4838
rect 3110 4839 3111 4840
rect 3192 4839 3193 4840
rect 3114 4841 3115 4842
rect 3253 4841 3254 4842
rect 3113 4843 3114 4844
rect 3144 4843 3145 4844
rect 3020 4845 3021 4846
rect 3143 4845 3144 4846
rect 3117 4847 3118 4848
rect 3235 4847 3236 4848
rect 3000 4849 3001 4850
rect 3116 4849 3117 4850
rect 3122 4849 3123 4850
rect 3207 4849 3208 4850
rect 3129 4851 3130 4852
rect 3156 4851 3157 4852
rect 3128 4853 3129 4854
rect 3216 4853 3217 4854
rect 3137 4855 3138 4856
rect 3222 4855 3223 4856
rect 3141 4857 3142 4858
rect 3189 4857 3190 4858
rect 3134 4859 3135 4860
rect 3140 4859 3141 4860
rect 3153 4859 3154 4860
rect 3210 4859 3211 4860
rect 3165 4861 3166 4862
rect 3201 4861 3202 4862
rect 3093 4863 3094 4864
rect 3200 4863 3201 4864
rect 3177 4865 3178 4866
rect 3293 4865 3294 4866
rect 3182 4867 3183 4868
rect 3213 4867 3214 4868
rect 3185 4869 3186 4870
rect 3259 4869 3260 4870
rect 3188 4871 3189 4872
rect 3262 4871 3263 4872
rect 3197 4873 3198 4874
rect 3274 4873 3275 4874
rect 3206 4875 3207 4876
rect 3280 4875 3281 4876
rect 3209 4877 3210 4878
rect 3283 4877 3284 4878
rect 3219 4879 3220 4880
rect 3296 4879 3297 4880
rect 3238 4881 3239 4882
rect 3256 4881 3257 4882
rect 3265 4881 3266 4882
rect 3334 4881 3335 4882
rect 3277 4883 3278 4884
rect 3328 4883 3329 4884
rect 3289 4885 3290 4886
rect 3300 4885 3301 4886
rect 3343 4885 3344 4886
rect 3350 4885 3351 4886
rect 2570 4894 2571 4895
rect 2703 4894 2704 4895
rect 2582 4896 2583 4897
rect 2831 4896 2832 4897
rect 2589 4898 2590 4899
rect 2804 4898 2805 4899
rect 2593 4900 2594 4901
rect 2846 4900 2847 4901
rect 2596 4902 2597 4903
rect 2664 4902 2665 4903
rect 2597 4904 2598 4905
rect 2620 4904 2621 4905
rect 2600 4906 2601 4907
rect 2840 4906 2841 4907
rect 2603 4908 2604 4909
rect 2667 4908 2668 4909
rect 2611 4910 2612 4911
rect 2780 4910 2781 4911
rect 2617 4912 2618 4913
rect 2783 4912 2784 4913
rect 2623 4914 2624 4915
rect 2864 4914 2865 4915
rect 2635 4916 2636 4917
rect 2642 4916 2643 4917
rect 2638 4918 2639 4919
rect 2658 4918 2659 4919
rect 2606 4920 2607 4921
rect 2638 4920 2639 4921
rect 2641 4920 2642 4921
rect 2655 4920 2656 4921
rect 2647 4922 2648 4923
rect 2879 4922 2880 4923
rect 2661 4924 2662 4925
rect 2861 4924 2862 4925
rect 2654 4926 2655 4927
rect 2861 4926 2862 4927
rect 2663 4928 2664 4929
rect 2894 4928 2895 4929
rect 2666 4930 2667 4931
rect 2789 4930 2790 4931
rect 2675 4932 2676 4933
rect 2692 4932 2693 4933
rect 2681 4934 2682 4935
rect 2798 4934 2799 4935
rect 2707 4936 2708 4937
rect 2735 4936 2736 4937
rect 2719 4938 2720 4939
rect 2732 4938 2733 4939
rect 2575 4940 2576 4941
rect 2732 4940 2733 4941
rect 2576 4942 2577 4943
rect 2583 4942 2584 4943
rect 2738 4942 2739 4943
rect 2747 4942 2748 4943
rect 2604 4944 2605 4945
rect 2747 4944 2748 4945
rect 2741 4946 2742 4947
rect 2750 4946 2751 4947
rect 2744 4948 2745 4949
rect 2915 4948 2916 4949
rect 2689 4950 2690 4951
rect 2915 4950 2916 4951
rect 2688 4952 2689 4953
rect 2912 4952 2913 4953
rect 2723 4954 2724 4955
rect 2912 4954 2913 4955
rect 2753 4956 2754 4957
rect 2876 4956 2877 4957
rect 2765 4958 2766 4959
rect 2768 4958 2769 4959
rect 2771 4958 2772 4959
rect 2774 4958 2775 4959
rect 2777 4958 2778 4959
rect 2792 4958 2793 4959
rect 2795 4958 2796 4959
rect 2897 4958 2898 4959
rect 2795 4960 2796 4961
rect 2810 4960 2811 4961
rect 2807 4962 2808 4963
rect 2816 4962 2817 4963
rect 2810 4964 2811 4965
rect 2819 4964 2820 4965
rect 2679 4966 2680 4967
rect 2819 4966 2820 4967
rect 2813 4968 2814 4969
rect 2834 4968 2835 4969
rect 2825 4970 2826 4971
rect 2843 4970 2844 4971
rect 2828 4972 2829 4973
rect 2843 4972 2844 4973
rect 2831 4974 2832 4975
rect 2855 4974 2856 4975
rect 2651 4976 2652 4977
rect 2855 4976 2856 4977
rect 2852 4978 2853 4979
rect 2858 4978 2859 4979
rect 2870 4978 2871 4979
rect 2891 4978 2892 4979
rect 2607 4980 2608 4981
rect 2891 4980 2892 4981
rect 2873 4982 2874 4983
rect 2888 4982 2889 4983
rect 2882 4984 2883 4985
rect 2885 4984 2886 4985
rect 2867 4986 2868 4987
rect 2882 4986 2883 4987
rect 2613 4988 2614 4989
rect 2867 4988 2868 4989
rect 2614 4990 2615 4991
rect 2726 4990 2727 4991
rect 2900 4990 2901 4991
rect 2903 4990 2904 4991
rect 2903 4992 2904 4993
rect 2909 4992 2910 4993
rect 2921 4992 2922 4993
rect 2927 4992 2928 4993
rect 2726 4994 2727 4995
rect 2927 4994 2928 4995
rect 2939 4994 2940 4995
rect 2945 4994 2946 4995
rect 2939 4996 2940 4997
rect 2966 4996 2967 4997
rect 2969 4996 2970 4997
rect 2981 4996 2982 4997
rect 2957 4998 2958 4999
rect 2969 4998 2970 4999
rect 2951 5000 2952 5001
rect 2957 5000 2958 5001
rect 2933 5002 2934 5003
rect 2951 5002 2952 5003
rect 2975 5002 2976 5003
rect 2993 5002 2994 5003
rect 2930 5004 2931 5005
rect 2975 5004 2976 5005
rect 2918 5006 2919 5007
rect 2930 5006 2931 5007
rect 2837 5008 2838 5009
rect 2918 5008 2919 5009
rect 2987 5008 2988 5009
rect 3116 5008 3117 5009
rect 2990 5010 2991 5011
rect 3026 5010 3027 5011
rect 2996 5012 2997 5013
rect 3008 5012 3009 5013
rect 2978 5014 2979 5015
rect 2996 5014 2997 5015
rect 2933 5016 2934 5017
rect 2978 5016 2979 5017
rect 3020 5016 3021 5017
rect 3071 5016 3072 5017
rect 3020 5018 3021 5019
rect 3194 5018 3195 5019
rect 2710 5020 2711 5021
rect 3195 5020 3196 5021
rect 3023 5022 3024 5023
rect 3032 5022 3033 5023
rect 3035 5022 3036 5023
rect 3140 5022 3141 5023
rect 3035 5024 3036 5025
rect 3125 5024 3126 5025
rect 3038 5026 3039 5027
rect 3177 5026 3178 5027
rect 3041 5028 3042 5029
rect 3183 5028 3184 5029
rect 3047 5030 3048 5031
rect 3056 5030 3057 5031
rect 3047 5032 3048 5033
rect 3065 5032 3066 5033
rect 3068 5032 3069 5033
rect 3107 5032 3108 5033
rect 3071 5034 3072 5035
rect 3203 5034 3204 5035
rect 3080 5036 3081 5037
rect 3089 5036 3090 5037
rect 2963 5038 2964 5039
rect 3080 5038 3081 5039
rect 2695 5040 2696 5041
rect 2963 5040 2964 5041
rect 3083 5040 3084 5041
rect 3092 5040 3093 5041
rect 3095 5040 3096 5041
rect 3098 5040 3099 5041
rect 3098 5042 3099 5043
rect 3101 5042 3102 5043
rect 3104 5042 3105 5043
rect 3214 5042 3215 5043
rect 3107 5044 3108 5045
rect 3110 5044 3111 5045
rect 3110 5046 3111 5047
rect 3113 5046 3114 5047
rect 3122 5046 3123 5047
rect 3134 5046 3135 5047
rect 3128 5048 3129 5049
rect 3212 5048 3213 5049
rect 3131 5050 3132 5051
rect 3233 5050 3234 5051
rect 3119 5052 3120 5053
rect 3232 5052 3233 5053
rect 3143 5054 3144 5055
rect 3239 5054 3240 5055
rect 3153 5056 3154 5057
rect 3161 5056 3162 5057
rect 3137 5058 3138 5059
rect 3152 5058 3153 5059
rect 3077 5060 3078 5061
rect 3137 5060 3138 5061
rect 3156 5060 3157 5061
rect 3164 5060 3165 5061
rect 2936 5062 2937 5063
rect 3155 5062 3156 5063
rect 3180 5062 3181 5063
rect 3185 5062 3186 5063
rect 3188 5062 3189 5063
rect 3256 5062 3257 5063
rect 3192 5064 3193 5065
rect 3197 5064 3198 5065
rect 3209 5064 3210 5065
rect 3253 5064 3254 5065
rect 3206 5066 3207 5067
rect 3208 5066 3209 5067
rect 3014 5068 3015 5069
rect 3205 5068 3206 5069
rect 3002 5070 3003 5071
rect 3014 5070 3015 5071
rect 2563 5079 2564 5080
rect 2774 5079 2775 5080
rect 2586 5081 2587 5082
rect 2590 5081 2591 5082
rect 2593 5081 2594 5082
rect 2741 5081 2742 5082
rect 2593 5083 2594 5084
rect 2951 5083 2952 5084
rect 2596 5085 2597 5086
rect 2867 5085 2868 5086
rect 2604 5087 2605 5088
rect 2852 5087 2853 5088
rect 2603 5089 2604 5090
rect 2843 5089 2844 5090
rect 2607 5091 2608 5092
rect 2638 5091 2639 5092
rect 2617 5093 2618 5094
rect 2620 5093 2621 5094
rect 2623 5093 2624 5094
rect 2915 5093 2916 5094
rect 2629 5095 2630 5096
rect 2641 5095 2642 5096
rect 2638 5097 2639 5098
rect 2891 5097 2892 5098
rect 2642 5099 2643 5100
rect 2882 5099 2883 5100
rect 2645 5101 2646 5102
rect 2647 5101 2648 5102
rect 2651 5101 2652 5102
rect 2897 5101 2898 5102
rect 2661 5103 2662 5104
rect 2675 5103 2676 5104
rect 2664 5105 2665 5106
rect 2894 5105 2895 5106
rect 2666 5107 2667 5108
rect 2837 5107 2838 5108
rect 2671 5109 2672 5110
rect 2771 5109 2772 5110
rect 2678 5111 2679 5112
rect 2819 5111 2820 5112
rect 2632 5113 2633 5114
rect 2819 5113 2820 5114
rect 2632 5115 2633 5116
rect 2846 5115 2847 5116
rect 2678 5117 2679 5118
rect 2714 5117 2715 5118
rect 2681 5119 2682 5120
rect 2870 5119 2871 5120
rect 2681 5121 2682 5122
rect 2900 5121 2901 5122
rect 2697 5123 2698 5124
rect 2703 5123 2704 5124
rect 2707 5123 2708 5124
rect 2726 5123 2727 5124
rect 2717 5125 2718 5126
rect 2891 5125 2892 5126
rect 2720 5127 2721 5128
rect 2732 5127 2733 5128
rect 2723 5129 2724 5130
rect 2735 5129 2736 5130
rect 2729 5131 2730 5132
rect 2930 5131 2931 5132
rect 2732 5133 2733 5134
rect 2738 5133 2739 5134
rect 2735 5135 2736 5136
rect 2753 5135 2754 5136
rect 2674 5137 2675 5138
rect 2753 5137 2754 5138
rect 2747 5139 2748 5140
rect 2876 5139 2877 5140
rect 2747 5141 2748 5142
rect 2765 5141 2766 5142
rect 2765 5143 2766 5144
rect 2795 5143 2796 5144
rect 2771 5145 2772 5146
rect 2777 5145 2778 5146
rect 2777 5147 2778 5148
rect 2789 5147 2790 5148
rect 2783 5149 2784 5150
rect 2807 5149 2808 5150
rect 2786 5151 2787 5152
rect 2810 5151 2811 5152
rect 2801 5153 2802 5154
rect 2825 5153 2826 5154
rect 2807 5155 2808 5156
rect 2831 5155 2832 5156
rect 2810 5157 2811 5158
rect 2885 5157 2886 5158
rect 2816 5159 2817 5160
rect 2918 5159 2919 5160
rect 2825 5161 2826 5162
rect 3077 5161 3078 5162
rect 2831 5163 2832 5164
rect 2849 5163 2850 5164
rect 2849 5165 2850 5166
rect 2864 5165 2865 5166
rect 2864 5167 2865 5168
rect 3080 5167 3081 5168
rect 2870 5169 2871 5170
rect 2903 5169 2904 5170
rect 2873 5171 2874 5172
rect 2888 5171 2889 5172
rect 2897 5171 2898 5172
rect 2933 5171 2934 5172
rect 2900 5173 2901 5174
rect 2936 5173 2937 5174
rect 2903 5175 2904 5176
rect 2984 5175 2985 5176
rect 2909 5177 2910 5178
rect 2927 5177 2928 5178
rect 2912 5179 2913 5180
rect 2915 5179 2916 5180
rect 2703 5181 2704 5182
rect 2912 5181 2913 5182
rect 2918 5181 2919 5182
rect 2939 5181 2940 5182
rect 2921 5183 2922 5184
rect 2978 5183 2979 5184
rect 2924 5185 2925 5186
rect 2957 5185 2958 5186
rect 2930 5187 2931 5188
rect 2945 5187 2946 5188
rect 2933 5189 2934 5190
rect 3116 5189 3117 5190
rect 2936 5191 2937 5192
rect 2987 5191 2988 5192
rect 2942 5193 2943 5194
rect 2969 5193 2970 5194
rect 2948 5195 2949 5196
rect 2981 5195 2982 5196
rect 2960 5197 2961 5198
rect 3023 5197 3024 5198
rect 2963 5199 2964 5200
rect 3137 5199 3138 5200
rect 2963 5201 2964 5202
rect 2996 5201 2997 5202
rect 2966 5203 2967 5204
rect 3177 5203 3178 5204
rect 2987 5205 2988 5206
rect 3056 5205 3057 5206
rect 2999 5207 3000 5208
rect 3092 5207 3093 5208
rect 3002 5209 3003 5210
rect 3014 5209 3015 5210
rect 3008 5211 3009 5212
rect 3014 5211 3015 5212
rect 3011 5213 3012 5214
rect 3164 5213 3165 5214
rect 3017 5215 3018 5216
rect 3068 5215 3069 5216
rect 3020 5217 3021 5218
rect 3205 5217 3206 5218
rect 3026 5219 3027 5220
rect 3158 5219 3159 5220
rect 3032 5221 3033 5222
rect 3107 5221 3108 5222
rect 3035 5223 3036 5224
rect 3067 5223 3068 5224
rect 3035 5225 3036 5226
rect 3071 5225 3072 5226
rect 3038 5227 3039 5228
rect 3095 5227 3096 5228
rect 3047 5229 3048 5230
rect 3174 5229 3175 5230
rect 2993 5231 2994 5232
rect 3048 5231 3049 5232
rect 3064 5231 3065 5232
rect 3119 5231 3120 5232
rect 3070 5233 3071 5234
rect 3086 5233 3087 5234
rect 3073 5235 3074 5236
rect 3083 5235 3084 5236
rect 3089 5235 3090 5236
rect 3146 5235 3147 5236
rect 3095 5237 3096 5238
rect 3161 5237 3162 5238
rect 3098 5239 3099 5240
rect 3202 5239 3203 5240
rect 3105 5241 3106 5242
rect 3262 5241 3263 5242
rect 3108 5243 3109 5244
rect 3180 5243 3181 5244
rect 3110 5245 3111 5246
rect 3170 5245 3171 5246
rect 3089 5247 3090 5248
rect 3170 5247 3171 5248
rect 3111 5249 3112 5250
rect 3183 5249 3184 5250
rect 3120 5251 3121 5252
rect 3192 5251 3193 5252
rect 3123 5253 3124 5254
rect 3152 5253 3153 5254
rect 3131 5255 3132 5256
rect 3235 5255 3236 5256
rect 3134 5257 3135 5258
rect 3232 5257 3233 5258
rect 3140 5259 3141 5260
rect 3246 5259 3247 5260
rect 3143 5261 3144 5262
rect 3253 5261 3254 5262
rect 3164 5263 3165 5264
rect 3208 5263 3209 5264
rect 2576 5272 2577 5273
rect 2720 5272 2721 5273
rect 2573 5274 2574 5275
rect 2576 5274 2577 5275
rect 2605 5274 2606 5275
rect 2629 5274 2630 5275
rect 2610 5276 2611 5277
rect 2849 5276 2850 5277
rect 2617 5278 2618 5279
rect 2620 5278 2621 5279
rect 2623 5278 2624 5279
rect 2664 5278 2665 5279
rect 2626 5280 2627 5281
rect 2831 5280 2832 5281
rect 2632 5282 2633 5283
rect 2635 5282 2636 5283
rect 2632 5284 2633 5285
rect 2876 5284 2877 5285
rect 2638 5286 2639 5287
rect 2810 5286 2811 5287
rect 2625 5288 2626 5289
rect 2811 5288 2812 5289
rect 2649 5290 2650 5291
rect 2753 5290 2754 5291
rect 2655 5292 2656 5293
rect 3120 5292 3121 5293
rect 2661 5294 2662 5295
rect 2688 5294 2689 5295
rect 2569 5296 2570 5297
rect 2689 5296 2690 5297
rect 2570 5298 2571 5299
rect 2774 5298 2775 5299
rect 2671 5300 2672 5301
rect 2747 5300 2748 5301
rect 2641 5302 2642 5303
rect 2748 5302 2749 5303
rect 2671 5304 2672 5305
rect 2692 5304 2693 5305
rect 2674 5306 2675 5307
rect 2816 5306 2817 5307
rect 2677 5308 2678 5309
rect 2723 5308 2724 5309
rect 2681 5310 2682 5311
rect 2870 5310 2871 5311
rect 2683 5312 2684 5313
rect 2765 5312 2766 5313
rect 2686 5314 2687 5315
rect 2697 5314 2698 5315
rect 2695 5316 2696 5317
rect 2732 5316 2733 5317
rect 2704 5318 2705 5319
rect 2735 5318 2736 5319
rect 2717 5320 2718 5321
rect 2900 5320 2901 5321
rect 2680 5322 2681 5323
rect 2717 5322 2718 5323
rect 2720 5322 2721 5323
rect 2835 5322 2836 5323
rect 2724 5324 2725 5325
rect 2871 5324 2872 5325
rect 2736 5326 2737 5327
rect 2783 5326 2784 5327
rect 2739 5328 2740 5329
rect 2786 5328 2787 5329
rect 2751 5330 2752 5331
rect 2771 5330 2772 5331
rect 2760 5332 2761 5333
rect 2777 5332 2778 5333
rect 2766 5334 2767 5335
rect 2868 5334 2869 5335
rect 2769 5336 2770 5337
rect 2918 5336 2919 5337
rect 2784 5338 2785 5339
rect 2807 5338 2808 5339
rect 2787 5340 2788 5341
rect 2801 5340 2802 5341
rect 2790 5342 2791 5343
rect 2819 5342 2820 5343
rect 2796 5344 2797 5345
rect 2837 5344 2838 5345
rect 2802 5346 2803 5347
rect 2855 5346 2856 5347
rect 2808 5348 2809 5349
rect 2852 5348 2853 5349
rect 2813 5350 2814 5351
rect 2817 5350 2818 5351
rect 2814 5352 2815 5353
rect 2858 5352 2859 5353
rect 2820 5354 2821 5355
rect 2861 5354 2862 5355
rect 2823 5356 2824 5357
rect 2873 5356 2874 5357
rect 2700 5358 2701 5359
rect 2874 5358 2875 5359
rect 2825 5360 2826 5361
rect 2984 5360 2985 5361
rect 2629 5362 2630 5363
rect 2826 5362 2827 5363
rect 2841 5362 2842 5363
rect 2891 5362 2892 5363
rect 2847 5364 2848 5365
rect 2915 5364 2916 5365
rect 2850 5366 2851 5367
rect 2903 5366 2904 5367
rect 2856 5368 2857 5369
rect 2897 5368 2898 5369
rect 2862 5370 2863 5371
rect 2909 5370 2910 5371
rect 2864 5372 2865 5373
rect 2981 5372 2982 5373
rect 2710 5374 2711 5375
rect 2865 5374 2866 5375
rect 2877 5374 2878 5375
rect 3009 5374 3010 5375
rect 2880 5376 2881 5377
rect 2930 5376 2931 5377
rect 2883 5378 2884 5379
rect 2933 5378 2934 5379
rect 2886 5380 2887 5381
rect 2924 5380 2925 5381
rect 2892 5382 2893 5383
rect 2942 5382 2943 5383
rect 2898 5384 2899 5385
rect 2936 5384 2937 5385
rect 2910 5386 2911 5387
rect 2960 5386 2961 5387
rect 2922 5388 2923 5389
rect 2999 5388 3000 5389
rect 2912 5390 2913 5391
rect 2999 5390 3000 5391
rect 2913 5392 2914 5393
rect 2963 5392 2964 5393
rect 2925 5394 2926 5395
rect 3002 5394 3003 5395
rect 2934 5396 2935 5397
rect 2987 5396 2988 5397
rect 2940 5398 2941 5399
rect 3035 5398 3036 5399
rect 2946 5400 2947 5401
rect 3037 5400 3038 5401
rect 2948 5402 2949 5403
rect 3002 5402 3003 5403
rect 2955 5404 2956 5405
rect 3067 5404 3068 5405
rect 2958 5406 2959 5407
rect 3011 5406 3012 5407
rect 2961 5408 2962 5409
rect 3014 5408 3015 5409
rect 2964 5410 2965 5411
rect 3017 5410 3018 5411
rect 2966 5412 2967 5413
rect 3048 5412 3049 5413
rect 2979 5414 2980 5415
rect 3032 5414 3033 5415
rect 2982 5416 2983 5417
rect 3045 5416 3046 5417
rect 3026 5418 3027 5419
rect 3154 5418 3155 5419
rect 3040 5420 3041 5421
rect 3147 5420 3148 5421
rect 3043 5422 3044 5423
rect 3089 5422 3090 5423
rect 3052 5424 3053 5425
rect 3108 5424 3109 5425
rect 3055 5426 3056 5427
rect 3076 5426 3077 5427
rect 3055 5428 3056 5429
rect 3111 5428 3112 5429
rect 3061 5430 3062 5431
rect 3143 5430 3144 5431
rect 3064 5432 3065 5433
rect 3140 5432 3141 5433
rect 3070 5434 3071 5435
rect 3102 5434 3103 5435
rect 3073 5436 3074 5437
rect 3079 5436 3080 5437
rect 3085 5436 3086 5437
rect 3123 5436 3124 5437
rect 3088 5438 3089 5439
rect 3170 5438 3171 5439
rect 3105 5440 3106 5441
rect 3167 5440 3168 5441
rect 2563 5449 2564 5450
rect 2576 5449 2577 5450
rect 2563 5451 2564 5452
rect 2566 5451 2567 5452
rect 2566 5453 2567 5454
rect 2605 5453 2606 5454
rect 2570 5455 2571 5456
rect 2686 5455 2687 5456
rect 2573 5457 2574 5458
rect 2689 5457 2690 5458
rect 2575 5459 2576 5460
rect 2582 5459 2583 5460
rect 2596 5459 2597 5460
rect 2635 5459 2636 5460
rect 2611 5461 2612 5462
rect 2638 5461 2639 5462
rect 2615 5463 2616 5464
rect 2823 5463 2824 5464
rect 2618 5465 2619 5466
rect 2702 5465 2703 5466
rect 2622 5467 2623 5468
rect 2802 5467 2803 5468
rect 2625 5469 2626 5470
rect 2796 5469 2797 5470
rect 2632 5471 2633 5472
rect 2650 5471 2651 5472
rect 2644 5473 2645 5474
rect 2677 5473 2678 5474
rect 2648 5475 2649 5476
rect 2820 5475 2821 5476
rect 2653 5477 2654 5478
rect 2695 5477 2696 5478
rect 2662 5479 2663 5480
rect 2771 5479 2772 5480
rect 2667 5481 2668 5482
rect 2692 5481 2693 5482
rect 2674 5483 2675 5484
rect 2710 5483 2711 5484
rect 2679 5485 2680 5486
rect 2736 5485 2737 5486
rect 2683 5487 2684 5488
rect 2739 5487 2740 5488
rect 2686 5489 2687 5490
rect 2795 5489 2796 5490
rect 2693 5491 2694 5492
rect 2883 5491 2884 5492
rect 2704 5493 2705 5494
rect 2720 5493 2721 5494
rect 2705 5495 2706 5496
rect 2748 5495 2749 5496
rect 2612 5497 2613 5498
rect 2747 5497 2748 5498
rect 2708 5499 2709 5500
rect 2751 5499 2752 5500
rect 2711 5501 2712 5502
rect 2865 5501 2866 5502
rect 2714 5503 2715 5504
rect 2760 5503 2761 5504
rect 2738 5505 2739 5506
rect 2808 5505 2809 5506
rect 2741 5507 2742 5508
rect 2784 5507 2785 5508
rect 2744 5509 2745 5510
rect 2787 5509 2788 5510
rect 2750 5511 2751 5512
rect 2811 5511 2812 5512
rect 2753 5513 2754 5514
rect 2814 5513 2815 5514
rect 2756 5515 2757 5516
rect 2790 5515 2791 5516
rect 2759 5517 2760 5518
rect 2826 5517 2827 5518
rect 2762 5519 2763 5520
rect 2862 5519 2863 5520
rect 2766 5521 2767 5522
rect 2847 5521 2848 5522
rect 2765 5523 2766 5524
rect 2880 5523 2881 5524
rect 2769 5525 2770 5526
rect 2856 5525 2857 5526
rect 2768 5527 2769 5528
rect 2817 5527 2818 5528
rect 2780 5529 2781 5530
rect 2835 5529 2836 5530
rect 2786 5531 2787 5532
rect 2841 5531 2842 5532
rect 2792 5533 2793 5534
rect 2850 5533 2851 5534
rect 2801 5535 2802 5536
rect 2910 5535 2911 5536
rect 2804 5537 2805 5538
rect 2868 5537 2869 5538
rect 2807 5539 2808 5540
rect 2871 5539 2872 5540
rect 2822 5541 2823 5542
rect 2967 5541 2968 5542
rect 2825 5543 2826 5544
rect 2886 5543 2887 5544
rect 2828 5545 2829 5546
rect 2992 5545 2993 5546
rect 2834 5547 2835 5548
rect 2925 5547 2926 5548
rect 2837 5549 2838 5550
rect 2922 5549 2923 5550
rect 2840 5551 2841 5552
rect 2892 5551 2893 5552
rect 2843 5553 2844 5554
rect 2913 5553 2914 5554
rect 2846 5555 2847 5556
rect 2919 5555 2920 5556
rect 2852 5557 2853 5558
rect 2891 5557 2892 5558
rect 2864 5559 2865 5560
rect 2934 5559 2935 5560
rect 2882 5561 2883 5562
rect 2982 5561 2983 5562
rect 2885 5563 2886 5564
rect 2940 5563 2941 5564
rect 2888 5565 2889 5566
rect 2964 5565 2965 5566
rect 2898 5567 2899 5568
rect 2995 5567 2996 5568
rect 2849 5569 2850 5570
rect 2898 5569 2899 5570
rect 2901 5569 2902 5570
rect 2985 5569 2986 5570
rect 2910 5571 2911 5572
rect 2923 5571 2924 5572
rect 2913 5573 2914 5574
rect 2933 5573 2934 5574
rect 2930 5575 2931 5576
rect 2961 5575 2962 5576
rect 2937 5577 2938 5578
rect 2946 5577 2947 5578
rect 2947 5579 2948 5580
rect 3040 5579 3041 5580
rect 2955 5581 2956 5582
rect 2960 5581 2961 5582
rect 2958 5583 2959 5584
rect 3013 5583 3014 5584
rect 2957 5585 2958 5586
rect 3058 5585 3059 5586
rect 2969 5587 2970 5588
rect 3094 5587 3095 5588
rect 2972 5589 2973 5590
rect 3052 5589 3053 5590
rect 2975 5591 2976 5592
rect 3055 5591 3056 5592
rect 2979 5593 2980 5594
rect 3002 5593 3003 5594
rect 3014 5593 3015 5594
rect 3018 5593 3019 5594
rect 3027 5593 3028 5594
rect 3085 5593 3086 5594
rect 3043 5595 3044 5596
rect 3108 5595 3109 5596
rect 3088 5597 3089 5598
rect 3098 5597 3099 5598
rect 2563 5606 2564 5607
rect 2578 5606 2579 5607
rect 2581 5606 2582 5607
rect 2653 5606 2654 5607
rect 2599 5608 2600 5609
rect 2702 5608 2703 5609
rect 2602 5610 2603 5611
rect 2768 5610 2769 5611
rect 2606 5612 2607 5613
rect 2684 5612 2685 5613
rect 2612 5614 2613 5615
rect 2759 5614 2760 5615
rect 2566 5616 2567 5617
rect 2760 5616 2761 5617
rect 2615 5618 2616 5619
rect 2756 5618 2757 5619
rect 2619 5620 2620 5621
rect 2714 5620 2715 5621
rect 2619 5622 2620 5623
rect 2644 5622 2645 5623
rect 2626 5624 2627 5625
rect 2741 5624 2742 5625
rect 2629 5626 2630 5627
rect 2744 5626 2745 5627
rect 2642 5628 2643 5629
rect 2705 5628 2706 5629
rect 2645 5630 2646 5631
rect 2708 5630 2709 5631
rect 2650 5632 2651 5633
rect 2717 5632 2718 5633
rect 2662 5634 2663 5635
rect 2705 5634 2706 5635
rect 2665 5636 2666 5637
rect 2714 5636 2715 5637
rect 2681 5638 2682 5639
rect 2738 5638 2739 5639
rect 2687 5640 2688 5641
rect 2792 5640 2793 5641
rect 2690 5642 2691 5643
rect 2795 5642 2796 5643
rect 2693 5644 2694 5645
rect 2837 5644 2838 5645
rect 2693 5646 2694 5647
rect 2747 5646 2748 5647
rect 2696 5648 2697 5649
rect 2750 5648 2751 5649
rect 2711 5650 2712 5651
rect 2798 5650 2799 5651
rect 2711 5652 2712 5653
rect 2771 5652 2772 5653
rect 2739 5654 2740 5655
rect 2780 5654 2781 5655
rect 2745 5656 2746 5657
rect 2786 5656 2787 5657
rect 2751 5658 2752 5659
rect 2804 5658 2805 5659
rect 2763 5660 2764 5661
rect 2825 5660 2826 5661
rect 2769 5662 2770 5663
rect 2840 5662 2841 5663
rect 2772 5664 2773 5665
rect 2828 5664 2829 5665
rect 2775 5666 2776 5667
rect 2852 5666 2853 5667
rect 2782 5668 2783 5669
rect 2882 5668 2883 5669
rect 2801 5670 2802 5671
rect 2822 5670 2823 5671
rect 2766 5672 2767 5673
rect 2800 5672 2801 5673
rect 2803 5672 2804 5673
rect 2849 5672 2850 5673
rect 2815 5674 2816 5675
rect 2846 5674 2847 5675
rect 2830 5676 2831 5677
rect 2888 5676 2889 5677
rect 2834 5678 2835 5679
rect 2916 5678 2917 5679
rect 2812 5680 2813 5681
rect 2833 5680 2834 5681
rect 2836 5680 2837 5681
rect 2913 5680 2914 5681
rect 2840 5682 2841 5683
rect 2937 5682 2938 5683
rect 2843 5684 2844 5685
rect 2947 5684 2948 5685
rect 2864 5686 2865 5687
rect 2891 5686 2892 5687
rect 2865 5688 2866 5689
rect 2957 5688 2958 5689
rect 2868 5690 2869 5691
rect 2960 5690 2961 5691
rect 2877 5692 2878 5693
rect 2972 5692 2973 5693
rect 2880 5694 2881 5695
rect 2975 5694 2976 5695
rect 2885 5696 2886 5697
rect 2894 5696 2895 5697
rect 2753 5698 2754 5699
rect 2893 5698 2894 5699
rect 2754 5700 2755 5701
rect 2807 5700 2808 5701
rect 2806 5702 2807 5703
rect 2818 5702 2819 5703
rect 2910 5702 2911 5703
rect 2919 5702 2920 5703
rect 2969 5702 2970 5703
rect 3021 5702 3022 5703
rect 3001 5704 3002 5705
rect 3008 5704 3009 5705
rect 2575 5713 2576 5714
rect 2619 5713 2620 5714
rect 2599 5715 2600 5716
rect 2606 5715 2607 5716
rect 2602 5717 2603 5718
rect 2684 5717 2685 5718
rect 2613 5719 2614 5720
rect 2693 5719 2694 5720
rect 2635 5721 2636 5722
rect 2696 5721 2697 5722
rect 2642 5723 2643 5724
rect 2675 5723 2676 5724
rect 2652 5725 2653 5726
rect 2714 5725 2715 5726
rect 2581 5727 2582 5728
rect 2713 5727 2714 5728
rect 2656 5729 2657 5730
rect 2681 5729 2682 5730
rect 2648 5731 2649 5732
rect 2655 5731 2656 5732
rect 2658 5731 2659 5732
rect 2685 5731 2686 5732
rect 2661 5733 2662 5734
rect 2711 5733 2712 5734
rect 2664 5735 2665 5736
rect 2717 5735 2718 5736
rect 2666 5737 2667 5738
rect 2705 5737 2706 5738
rect 2678 5739 2679 5740
rect 2694 5739 2695 5740
rect 2641 5741 2642 5742
rect 2679 5741 2680 5742
rect 2682 5741 2683 5742
rect 2697 5741 2698 5742
rect 2690 5743 2691 5744
rect 2754 5743 2755 5744
rect 2687 5745 2688 5746
rect 2691 5745 2692 5746
rect 2707 5745 2708 5746
rect 2739 5745 2740 5746
rect 2719 5747 2720 5748
rect 2734 5747 2735 5748
rect 2723 5749 2724 5750
rect 2745 5749 2746 5750
rect 2728 5751 2729 5752
rect 2772 5751 2773 5752
rect 2730 5753 2731 5754
rect 2751 5753 2752 5754
rect 2731 5755 2732 5756
rect 2775 5755 2776 5756
rect 2737 5757 2738 5758
rect 2755 5757 2756 5758
rect 2740 5759 2741 5760
rect 2800 5759 2801 5760
rect 2746 5761 2747 5762
rect 2815 5761 2816 5762
rect 2761 5763 2762 5764
rect 2806 5763 2807 5764
rect 2763 5765 2764 5766
rect 2769 5765 2770 5766
rect 2764 5767 2765 5768
rect 2847 5767 2848 5768
rect 2773 5769 2774 5770
rect 2830 5769 2831 5770
rect 2779 5771 2780 5772
rect 2812 5771 2813 5772
rect 2789 5773 2790 5774
rect 2877 5773 2878 5774
rect 2803 5775 2804 5776
rect 2833 5775 2834 5776
rect 2836 5775 2837 5776
rect 2843 5775 2844 5776
rect 2862 5775 2863 5776
rect 2865 5775 2866 5776
rect 2868 5775 2869 5776
rect 2874 5775 2875 5776
rect 2880 5775 2881 5776
rect 2883 5775 2884 5776
rect 2617 5784 2618 5785
rect 2761 5784 2762 5785
rect 2644 5786 2645 5787
rect 2664 5786 2665 5787
rect 2648 5788 2649 5789
rect 2789 5788 2790 5789
rect 2651 5790 2652 5791
rect 2661 5790 2662 5791
rect 2665 5792 2666 5793
rect 2685 5792 2686 5793
rect 2674 5794 2675 5795
rect 2691 5794 2692 5795
rect 2677 5796 2678 5797
rect 2697 5796 2698 5797
rect 2694 5798 2695 5799
rect 2703 5798 2704 5799
rect 2707 5798 2708 5799
rect 2728 5798 2729 5799
rect 2710 5800 2711 5801
rect 2731 5800 2732 5801
rect 2713 5802 2714 5803
rect 2719 5802 2720 5803
rect 2737 5802 2738 5803
rect 2773 5802 2774 5803
rect 2740 5804 2741 5805
rect 2767 5804 2768 5805
rect 2746 5806 2747 5807
rect 2786 5806 2787 5807
rect 2764 5808 2765 5809
rect 2770 5808 2771 5809
rect 2623 5817 2624 5818
rect 2737 5817 2738 5818
rect 2653 5819 2654 5820
rect 2677 5819 2678 5820
rect 2656 5821 2657 5822
rect 2668 5821 2669 5822
rect 2665 5823 2666 5824
rect 2674 5823 2675 5824
rect 2707 5823 2708 5824
rect 2716 5823 2717 5824
rect 2710 5825 2711 5826
rect 2713 5825 2714 5826
<< end >>
