magic
tech scmos
timestamp 1395743115
<< m1p >>
use CELL  1
transform -1 0 1498 0 1 10092
box 0 0 6 6
use CELL  2
transform -1 0 1443 0 1 3126
box 0 0 6 6
use CELL  3
transform -1 0 1502 0 1 2557
box 0 0 6 6
use CELL  4
transform -1 0 3006 0 1 8585
box 0 0 6 6
use CELL  5
transform -1 0 1456 0 1 9631
box 0 0 6 6
use CELL  6
transform -1 0 1478 0 1 1571
box 0 0 6 6
use CELL  7
transform -1 0 2698 0 1 1571
box 0 0 6 6
use CELL  8
transform -1 0 1501 0 1 11105
box 0 0 6 6
use CELL  9
transform -1 0 3222 0 1 6808
box 0 0 6 6
use CELL  10
transform -1 0 2231 0 1 10850
box 0 0 6 6
use CELL  11
transform -1 0 2419 0 1 1182
box 0 0 6 6
use CELL  12
transform -1 0 3393 0 1 4917
box 0 0 6 6
use CELL  13
transform -1 0 3439 0 1 6171
box 0 0 6 6
use CELL  14
transform -1 0 3156 0 1 8006
box 0 0 6 6
use CELL  15
transform -1 0 1537 0 1 6171
box 0 0 6 6
use CELL  16
transform -1 0 2630 0 1 1571
box 0 0 6 6
use CELL  17
transform -1 0 2412 0 1 1182
box 0 0 6 6
use CELL  18
transform -1 0 2951 0 1 8585
box 0 0 6 6
use CELL  19
transform -1 0 1464 0 1 2028
box 0 0 6 6
use CELL  20
transform -1 0 1512 0 1 3699
box 0 0 6 6
use CELL  21
transform -1 0 1435 0 1 8585
box 0 0 6 6
use CELL  22
transform -1 0 1597 0 1 1182
box 0 0 6 6
use CELL  23
transform -1 0 1480 0 1 3699
box 0 0 6 6
use CELL  24
transform -1 0 1454 0 1 8006
box 0 0 6 6
use CELL  25
transform -1 0 2410 0 1 10509
box 0 0 6 6
use CELL  26
transform -1 0 3248 0 1 6808
box 0 0 6 6
use CELL  27
transform -1 0 1482 0 1 11321
box 0 0 6 6
use CELL  28
transform -1 0 3235 0 1 4917
box 0 0 6 6
use CELL  29
transform -1 0 1590 0 1 9128
box 0 0 6 6
use CELL  30
transform -1 0 1512 0 1 4294
box 0 0 6 6
use CELL  31
transform -1 0 1447 0 1 8006
box 0 0 6 6
use CELL  32
transform -1 0 1428 0 1 5572
box 0 0 6 6
use CELL  33
transform -1 0 2622 0 1 9128
box 0 0 6 6
use CELL  34
transform -1 0 1530 0 1 3699
box 0 0 6 6
use CELL  35
transform -1 0 1435 0 1 5572
box 0 0 6 6
use CELL  36
transform -1 0 1429 0 1 1571
box 0 0 6 6
use CELL  37
transform -1 0 2835 0 1 2028
box 0 0 6 6
use CELL  38
transform -1 0 1531 0 1 4294
box 0 0 6 6
use CELL  39
transform -1 0 1429 0 1 6808
box 0 0 6 6
use CELL  40
transform -1 0 1436 0 1 4294
box 0 0 6 6
use CELL  41
transform -1 0 1603 0 1 4294
box 0 0 6 6
use CELL  42
transform -1 0 3083 0 1 8006
box 0 0 6 6
use CELL  43
transform -1 0 1485 0 1 1571
box 0 0 6 6
use CELL  44
transform -1 0 1505 0 1 6808
box 0 0 6 6
use CELL  45
transform -1 0 1436 0 1 3126
box 0 0 6 6
use CELL  46
transform -1 0 2573 0 1 10092
box 0 0 6 6
use CELL  47
transform -1 0 1486 0 1 5572
box 0 0 6 6
use CELL  48
transform -1 0 3229 0 1 4294
box 0 0 6 6
use CELL  49
transform -1 0 2443 0 1 10509
box 0 0 6 6
use CELL  50
transform -1 0 2357 0 1 1182
box 0 0 6 6
use CELL  51
transform -1 0 3032 0 1 8585
box 0 0 6 6
use CELL  52
transform -1 0 3169 0 1 3126
box 0 0 6 6
use CELL  53
transform -1 0 1507 0 1 1182
box 0 0 6 6
use CELL  54
transform -1 0 3284 0 1 6171
box 0 0 6 6
use CELL  55
transform -1 0 1924 0 1 901
box 0 0 6 6
use CELL  56
transform -1 0 3432 0 1 6171
box 0 0 6 6
use CELL  57
transform -1 0 2916 0 1 2028
box 0 0 6 6
use CELL  58
transform -1 0 2588 0 1 1571
box 0 0 6 6
use CELL  59
transform -1 0 1479 0 1 901
box 0 0 6 6
use CELL  60
transform -1 0 2642 0 1 10092
box 0 0 6 6
use CELL  61
transform -1 0 1577 0 1 10092
box 0 0 6 6
use CELL  62
transform -1 0 3316 0 1 4917
box 0 0 6 6
use CELL  63
transform -1 0 3241 0 1 6808
box 0 0 6 6
use CELL  64
transform -1 0 3131 0 1 8006
box 0 0 6 6
use CELL  65
transform -1 0 2747 0 1 8585
box 0 0 6 6
use CELL  66
transform -1 0 3424 0 1 5572
box 0 0 6 6
use CELL  67
transform -1 0 1486 0 1 901
box 0 0 6 6
use CELL  68
transform -1 0 1934 0 1 11105
box 0 0 6 6
use CELL  69
transform -1 0 2436 0 1 10509
box 0 0 6 6
use CELL  70
transform -1 0 2585 0 1 10092
box 0 0 6 6
use CELL  71
transform -1 0 2725 0 1 1571
box 0 0 6 6
use CELL  72
transform -1 0 3102 0 1 2557
box 0 0 6 6
use CELL  73
transform -1 0 1505 0 1 4917
box 0 0 6 6
use CELL  74
transform -1 0 3070 0 1 8585
box 0 0 6 6
use CELL  75
transform -1 0 1578 0 1 9631
box 0 0 6 6
use CELL  76
transform -1 0 3198 0 1 7369
box 0 0 6 6
use CELL  77
transform -1 0 1449 0 1 11105
box 0 0 6 6
use CELL  78
transform -1 0 1457 0 1 1182
box 0 0 6 6
use CELL  79
transform -1 0 1443 0 1 1182
box 0 0 6 6
use CELL  80
transform -1 0 3217 0 1 4294
box 0 0 6 6
use CELL  81
transform -1 0 3297 0 1 7369
box 0 0 6 6
use CELL  82
transform -1 0 1548 0 1 732
box 0 0 6 6
use CELL  83
transform -1 0 1961 0 1 11105
box 0 0 6 6
use CELL  84
transform -1 0 1506 0 1 11264
box 0 0 6 6
use CELL  85
transform -1 0 2850 0 1 9128
box 0 0 6 6
use CELL  86
transform -1 0 1517 0 1 5572
box 0 0 6 6
use CELL  87
transform -1 0 2970 0 1 9128
box 0 0 6 6
use CELL  88
transform -1 0 2169 0 1 10850
box 0 0 6 6
use CELL  89
transform -1 0 1523 0 1 10092
box 0 0 6 6
use CELL  90
transform -1 0 1468 0 1 10092
box 0 0 6 6
use CELL  91
transform -1 0 1711 0 1 4294
box 0 0 6 6
use CELL  92
transform -1 0 1429 0 1 3699
box 0 0 6 6
use CELL  93
transform -1 0 1443 0 1 6808
box 0 0 6 6
use CELL  94
transform -1 0 2648 0 1 10092
box 0 0 6 6
use CELL  95
transform -1 0 3398 0 1 5572
box 0 0 6 6
use CELL  96
transform -1 0 1543 0 1 4917
box 0 0 6 6
use CELL  97
transform -1 0 1422 0 1 1182
box 0 0 6 6
use CELL  98
transform -1 0 1600 0 1 8006
box 0 0 6 6
use CELL  99
transform -1 0 1436 0 1 6171
box 0 0 6 6
use CELL  100
transform -1 0 3379 0 1 4917
box 0 0 6 6
use CELL  101
transform -1 0 3157 0 1 3699
box 0 0 6 6
use CELL  102
transform -1 0 2320 0 1 10509
box 0 0 6 6
use CELL  103
transform -1 0 1552 0 1 901
box 0 0 6 6
use CELL  104
transform -1 0 1455 0 1 2557
box 0 0 6 6
use CELL  105
transform -1 0 1498 0 1 901
box 0 0 6 6
use CELL  106
transform -1 0 2637 0 1 1571
box 0 0 6 6
use CELL  107
transform -1 0 2433 0 1 1182
box 0 0 6 6
use CELL  108
transform -1 0 2930 0 1 2028
box 0 0 6 6
use CELL  109
transform -1 0 1473 0 1 8006
box 0 0 6 6
use CELL  110
transform -1 0 3242 0 1 4917
box 0 0 6 6
use CELL  111
transform -1 0 1436 0 1 6808
box 0 0 6 6
use CELL  112
transform -1 0 2609 0 1 10092
box 0 0 6 6
use CELL  113
transform -1 0 1529 0 1 8585
box 0 0 6 6
use CELL  114
transform -1 0 1466 0 1 8006
box 0 0 6 6
use CELL  115
transform -1 0 1531 0 1 4917
box 0 0 6 6
use CELL  116
transform -1 0 1589 0 1 6808
box 0 0 6 6
use CELL  117
transform -1 0 2008 0 1 901
box 0 0 6 6
use CELL  118
transform -1 0 2674 0 1 1571
box 0 0 6 6
use CELL  119
transform -1 0 1448 0 1 901
box 0 0 6 6
use CELL  120
transform -1 0 1628 0 1 11264
box 0 0 6 6
use CELL  121
transform -1 0 2939 0 1 9128
box 0 0 6 6
use CELL  122
transform -1 0 1442 0 1 10092
box 0 0 6 6
use CELL  123
transform -1 0 1442 0 1 9631
box 0 0 6 6
use CELL  124
transform -1 0 1464 0 1 1571
box 0 0 6 6
use CELL  125
transform -1 0 3029 0 1 2557
box 0 0 6 6
use CELL  126
transform -1 0 1504 0 1 2028
box 0 0 6 6
use CELL  127
transform -1 0 1460 0 1 10509
box 0 0 6 6
use CELL  128
transform -1 0 3279 0 1 4294
box 0 0 6 6
use CELL  129
transform -1 0 1543 0 1 5572
box 0 0 6 6
use CELL  130
transform -1 0 2457 0 1 10509
box 0 0 6 6
use CELL  131
transform -1 0 3405 0 1 5572
box 0 0 6 6
use CELL  132
transform -1 0 1523 0 1 7369
box 0 0 6 6
use CELL  133
transform -1 0 3175 0 1 8006
box 0 0 6 6
use CELL  134
transform -1 0 1512 0 1 732
box 0 0 6 6
use CELL  135
transform -1 0 1620 0 1 732
box 0 0 6 6
use CELL  136
transform -1 0 3017 0 1 2557
box 0 0 6 6
use CELL  137
transform -1 0 3120 0 1 3699
box 0 0 6 6
use CELL  138
transform -1 0 1468 0 1 8585
box 0 0 6 6
use CELL  139
transform -1 0 1456 0 1 8585
box 0 0 6 6
use CELL  140
transform -1 0 1948 0 1 11105
box 0 0 6 6
use CELL  141
transform -1 0 1566 0 1 9631
box 0 0 6 6
use CELL  142
transform -1 0 1457 0 1 1571
box 0 0 6 6
use CELL  143
transform -1 0 1428 0 1 7369
box 0 0 6 6
use CELL  144
transform -1 0 2932 0 1 9128
box 0 0 6 6
use CELL  145
transform -1 0 1529 0 1 9631
box 0 0 6 6
use CELL  146
transform -1 0 1554 0 1 9128
box 0 0 6 6
use CELL  147
transform -1 0 3449 0 1 5572
box 0 0 6 6
use CELL  148
transform -1 0 1456 0 1 9128
box 0 0 6 6
use CELL  149
transform -1 0 3161 0 1 6808
box 0 0 6 6
use CELL  150
transform -1 0 3370 0 1 6171
box 0 0 6 6
use CELL  151
transform -1 0 3266 0 1 6808
box 0 0 6 6
use CELL  152
transform -1 0 2429 0 1 10509
box 0 0 6 6
use CELL  153
transform -1 0 1491 0 1 10850
box 0 0 6 6
use CELL  154
transform -1 0 3193 0 1 3699
box 0 0 6 6
use CELL  155
transform -1 0 3322 0 1 7369
box 0 0 6 6
use CELL  156
transform -1 0 1492 0 1 1571
box 0 0 6 6
use CELL  157
transform -1 0 1467 0 1 10509
box 0 0 6 6
use CELL  158
transform -1 0 3298 0 1 6808
box 0 0 6 6
use CELL  159
transform -1 0 1435 0 1 7369
box 0 0 6 6
use CELL  160
transform -1 0 2739 0 1 9631
box 0 0 6 6
use CELL  161
transform -1 0 3286 0 1 4294
box 0 0 6 6
use CELL  162
transform -1 0 3175 0 1 3699
box 0 0 6 6
use CELL  163
transform -1 0 2720 0 1 9631
box 0 0 6 6
use CELL  164
transform -1 0 2464 0 1 10509
box 0 0 6 6
use CELL  165
transform -1 0 3168 0 1 6808
box 0 0 6 6
use CELL  166
transform -1 0 2440 0 1 1182
box 0 0 6 6
use CELL  167
transform -1 0 1614 0 1 11264
box 0 0 6 6
use CELL  168
transform -1 0 2581 0 1 1571
box 0 0 6 6
use CELL  169
transform -1 0 1455 0 1 901
box 0 0 6 6
use CELL  170
transform -1 0 1464 0 1 1182
box 0 0 6 6
use CELL  171
transform -1 0 1464 0 1 11105
box 0 0 6 6
use CELL  172
transform -1 0 1751 0 1 7369
box 0 0 6 6
use CELL  173
transform -1 0 1448 0 1 11264
box 0 0 6 6
use CELL  174
transform -1 0 1429 0 1 2028
box 0 0 6 6
use CELL  175
transform -1 0 3304 0 1 7369
box 0 0 6 6
use CELL  176
transform -1 0 3277 0 1 6171
box 0 0 6 6
use CELL  177
transform -1 0 2925 0 1 9128
box 0 0 6 6
use CELL  178
transform -1 0 2918 0 1 9128
box 0 0 6 6
use CELL  179
transform -1 0 1626 0 1 3699
box 0 0 6 6
use CELL  180
transform -1 0 3252 0 1 3126
box 0 0 6 6
use CELL  181
transform -1 0 2902 0 1 2028
box 0 0 6 6
use CELL  182
transform -1 0 3290 0 1 7369
box 0 0 6 6
use CELL  183
transform -1 0 1442 0 1 732
box 0 0 6 6
use CELL  184
transform -1 0 2545 0 1 1571
box 0 0 6 6
use CELL  185
transform -1 0 1480 0 1 4917
box 0 0 6 6
use CELL  186
transform -1 0 2732 0 1 9631
box 0 0 6 6
use CELL  187
transform -1 0 1436 0 1 2028
box 0 0 6 6
use CELL  188
transform -1 0 1460 0 1 10850
box 0 0 6 6
use CELL  189
transform -1 0 1429 0 1 3126
box 0 0 6 6
use CELL  190
transform -1 0 3214 0 1 3699
box 0 0 6 6
use CELL  191
transform -1 0 1450 0 1 2028
box 0 0 6 6
use CELL  192
transform -1 0 3013 0 1 8585
box 0 0 6 6
use CELL  193
transform -1 0 3157 0 1 3126
box 0 0 6 6
use CELL  194
transform -1 0 3412 0 1 5572
box 0 0 6 6
use CELL  195
transform -1 0 1915 0 1 11105
box 0 0 6 6
use CELL  196
transform -1 0 3307 0 1 4294
box 0 0 6 6
use CELL  197
transform -1 0 3084 0 1 8585
box 0 0 6 6
use CELL  198
transform -1 0 1516 0 1 10092
box 0 0 6 6
use CELL  199
transform -1 0 1457 0 1 732
box 0 0 6 6
use CELL  200
transform -1 0 3231 0 1 3126
box 0 0 6 6
use CELL  201
transform -1 0 1453 0 1 10850
box 0 0 6 6
use CELL  202
transform -1 0 2628 0 1 9631
box 0 0 6 6
use CELL  203
transform -1 0 3066 0 1 2557
box 0 0 6 6
use CELL  204
transform -1 0 3335 0 1 4917
box 0 0 6 6
use CELL  205
transform -1 0 1436 0 1 4917
box 0 0 6 6
use CELL  206
transform -1 0 1428 0 1 8006
box 0 0 6 6
use CELL  207
transform -1 0 3054 0 1 3699
box 0 0 6 6
use CELL  208
transform -1 0 3109 0 1 2557
box 0 0 6 6
use CELL  209
transform -1 0 1955 0 1 11105
box 0 0 6 6
use CELL  210
transform -1 0 1466 0 1 732
box 0 0 6 6
use CELL  211
transform -1 0 1428 0 1 9128
box 0 0 6 6
use CELL  212
transform -1 0 1428 0 1 11105
box 0 0 6 6
use CELL  213
transform -1 0 1442 0 1 5572
box 0 0 6 6
use CELL  214
transform -1 0 1994 0 1 901
box 0 0 6 6
use CELL  215
transform -1 0 3325 0 1 5572
box 0 0 6 6
use CELL  216
transform -1 0 1500 0 1 3126
box 0 0 6 6
use CELL  217
transform -1 0 2872 0 1 2028
box 0 0 6 6
use CELL  218
transform -1 0 1507 0 1 3126
box 0 0 6 6
use CELL  219
transform -1 0 1488 0 1 2557
box 0 0 6 6
use CELL  220
transform -1 0 3116 0 1 2557
box 0 0 6 6
use CELL  221
transform -1 0 1495 0 1 2557
box 0 0 6 6
use CELL  222
transform -1 0 1558 0 1 10509
box 0 0 6 6
use CELL  223
transform -1 0 3400 0 1 6171
box 0 0 6 6
use CELL  224
transform -1 0 1475 0 1 3126
box 0 0 6 6
use CELL  225
transform -1 0 1613 0 1 6808
box 0 0 6 6
use CELL  226
transform -1 0 1476 0 1 2557
box 0 0 6 6
use CELL  227
transform -1 0 3168 0 1 8006
box 0 0 6 6
use CELL  228
transform -1 0 1446 0 1 10850
box 0 0 6 6
use CELL  229
transform -1 0 1475 0 1 9631
box 0 0 6 6
use CELL  230
transform -1 0 1505 0 1 4294
box 0 0 6 6
use CELL  231
transform -1 0 2394 0 1 1182
box 0 0 6 6
use CELL  232
transform -1 0 2969 0 1 2557
box 0 0 6 6
use CELL  233
transform -1 0 3059 0 1 2557
box 0 0 6 6
use CELL  234
transform -1 0 3077 0 1 8585
box 0 0 6 6
use CELL  235
transform -1 0 2712 0 1 1571
box 0 0 6 6
use CELL  236
transform -1 0 1484 0 1 10850
box 0 0 6 6
use CELL  237
transform -1 0 1478 0 1 2028
box 0 0 6 6
use CELL  238
transform -1 0 1512 0 1 4917
box 0 0 6 6
use CELL  239
transform -1 0 3365 0 1 4917
box 0 0 6 6
use CELL  240
transform -1 0 1434 0 1 11264
box 0 0 6 6
use CELL  241
transform -1 0 3071 0 1 8006
box 0 0 6 6
use CELL  242
transform -1 0 1627 0 1 732
box 0 0 6 6
use CELL  243
transform -1 0 2906 0 1 9128
box 0 0 6 6
use CELL  244
transform -1 0 1487 0 1 6171
box 0 0 6 6
use CELL  245
transform -1 0 1422 0 1 2028
box 0 0 6 6
use CELL  246
transform -1 0 2635 0 1 10092
box 0 0 6 6
use CELL  247
transform -1 0 3194 0 1 3126
box 0 0 6 6
use CELL  248
transform -1 0 1582 0 1 8006
box 0 0 6 6
use CELL  249
transform -1 0 1469 0 1 2557
box 0 0 6 6
use CELL  250
transform -1 0 1480 0 1 6171
box 0 0 6 6
use CELL  251
transform -1 0 1922 0 1 11105
box 0 0 6 6
use CELL  252
transform -1 0 3254 0 1 4294
box 0 0 6 6
use CELL  253
transform -1 0 3221 0 1 3699
box 0 0 6 6
use CELL  254
transform -1 0 3245 0 1 3126
box 0 0 6 6
use CELL  255
transform -1 0 2746 0 1 9631
box 0 0 6 6
use CELL  256
transform -1 0 1488 0 1 1182
box 0 0 6 6
use CELL  257
transform -1 0 3039 0 1 8585
box 0 0 6 6
use CELL  258
transform -1 0 2034 0 1 901
box 0 0 6 6
use CELL  259
transform -1 0 1436 0 1 3699
box 0 0 6 6
use CELL  260
transform -1 0 1614 0 1 3699
box 0 0 6 6
use CELL  261
transform -1 0 1641 0 1 732
box 0 0 6 6
use CELL  262
transform -1 0 3431 0 1 5572
box 0 0 6 6
use CELL  263
transform -1 0 1442 0 1 11105
box 0 0 6 6
use CELL  264
transform -1 0 1603 0 1 3126
box 0 0 6 6
use CELL  265
transform -1 0 3273 0 1 6808
box 0 0 6 6
use CELL  266
transform -1 0 1621 0 1 11264
box 0 0 6 6
use CELL  267
transform -1 0 3224 0 1 3126
box 0 0 6 6
use CELL  268
transform -1 0 2555 0 1 10092
box 0 0 6 6
use CELL  269
transform -1 0 2899 0 1 9128
box 0 0 6 6
use CELL  270
transform -1 0 1479 0 1 5572
box 0 0 6 6
use CELL  271
transform -1 0 1487 0 1 4294
box 0 0 6 6
use CELL  272
transform -1 0 3356 0 1 6171
box 0 0 6 6
use CELL  273
transform -1 0 1549 0 1 6171
box 0 0 6 6
use CELL  274
transform -1 0 1829 0 1 6808
box 0 0 6 6
use CELL  275
transform -1 0 3302 0 1 4917
box 0 0 6 6
use CELL  276
transform -1 0 3214 0 1 8006
box 0 0 6 6
use CELL  277
transform -1 0 3372 0 1 4917
box 0 0 6 6
use CELL  278
transform -1 0 1607 0 1 8006
box 0 0 6 6
use CELL  279
transform -1 0 2041 0 1 901
box 0 0 6 6
use CELL  280
transform -1 0 3079 0 1 3126
box 0 0 6 6
use CELL  281
transform -1 0 3305 0 1 6808
box 0 0 6 6
use CELL  282
transform -1 0 2719 0 1 1571
box 0 0 6 6
use CELL  283
transform -1 0 1442 0 1 9128
box 0 0 6 6
use CELL  284
transform -1 0 3446 0 1 6171
box 0 0 6 6
use CELL  285
transform -1 0 2035 0 1 6171
box 0 0 6 6
use CELL  286
transform -1 0 1480 0 1 7369
box 0 0 6 6
use CELL  287
transform -1 0 1462 0 1 2557
box 0 0 6 6
use CELL  288
transform -1 0 2828 0 1 2028
box 0 0 6 6
use CELL  289
transform -1 0 1429 0 1 4917
box 0 0 6 6
use CELL  290
transform -1 0 3123 0 1 2557
box 0 0 6 6
use CELL  291
transform -1 0 1463 0 1 9631
box 0 0 6 6
use CELL  292
transform -1 0 3332 0 1 5572
box 0 0 6 6
use CELL  293
transform -1 0 1536 0 1 9631
box 0 0 6 6
use CELL  294
transform -1 0 3271 0 1 7369
box 0 0 6 6
use CELL  295
transform -1 0 1577 0 1 8585
box 0 0 6 6
use CELL  296
transform -1 0 1487 0 1 4917
box 0 0 6 6
use CELL  297
transform -1 0 1517 0 1 8585
box 0 0 6 6
use CELL  298
transform -1 0 1481 0 1 6808
box 0 0 6 6
use CELL  299
transform -1 0 2664 0 1 3699
box 0 0 6 6
use CELL  300
transform -1 0 1635 0 1 10850
box 0 0 6 6
use CELL  301
transform -1 0 2195 0 1 10850
box 0 0 6 6
use CELL  302
transform -1 0 3293 0 1 4294
box 0 0 6 6
use CELL  303
transform -1 0 2753 0 1 9631
box 0 0 6 6
use CELL  304
transform -1 0 1471 0 1 2028
box 0 0 6 6
use CELL  305
transform -1 0 3145 0 1 4294
box 0 0 6 6
use CELL  306
transform -1 0 1605 0 1 732
box 0 0 6 6
use CELL  307
transform -1 0 1422 0 1 1571
box 0 0 6 6
use CELL  308
transform -1 0 2447 0 1 1182
box 0 0 6 6
use CELL  309
transform -1 0 1449 0 1 5572
box 0 0 6 6
use CELL  310
transform -1 0 1524 0 1 5572
box 0 0 6 6
use CELL  311
transform -1 0 3336 0 1 7369
box 0 0 6 6
use CELL  312
transform -1 0 1455 0 1 11105
box 0 0 6 6
use CELL  313
transform -1 0 1563 0 1 10850
box 0 0 6 6
use CELL  314
transform -1 0 1487 0 1 3699
box 0 0 6 6
use CELL  315
transform -1 0 3025 0 1 8585
box 0 0 6 6
use CELL  316
transform -1 0 3138 0 1 3699
box 0 0 6 6
use CELL  317
transform -1 0 2899 0 1 3126
box 0 0 6 6
use CELL  318
transform -1 0 3182 0 1 8006
box 0 0 6 6
use CELL  319
transform -1 0 1515 0 1 8006
box 0 0 6 6
use CELL  320
transform -1 0 3109 0 1 3126
box 0 0 6 6
use CELL  321
transform -1 0 3272 0 1 4294
box 0 0 6 6
use CELL  322
transform -1 0 1428 0 1 8585
box 0 0 6 6
use CELL  323
transform -1 0 1443 0 1 6171
box 0 0 6 6
use CELL  324
transform -1 0 1461 0 1 3126
box 0 0 6 6
use CELL  325
transform -1 0 1976 0 1 901
box 0 0 6 6
use CELL  326
transform -1 0 1467 0 1 901
box 0 0 6 6
use CELL  327
transform -1 0 3200 0 1 3699
box 0 0 6 6
use CELL  328
transform -1 0 1442 0 1 8585
box 0 0 6 6
use CELL  329
transform -1 0 1517 0 1 6808
box 0 0 6 6
use CELL  330
transform -1 0 1457 0 1 2028
box 0 0 6 6
use CELL  331
transform -1 0 1473 0 1 4294
box 0 0 6 6
use CELL  332
transform -1 0 1473 0 1 4917
box 0 0 6 6
use CELL  333
transform -1 0 1503 0 1 10509
box 0 0 6 6
use CELL  334
transform -1 0 2392 0 1 10509
box 0 0 6 6
use CELL  335
transform -1 0 3207 0 1 8006
box 0 0 6 6
use CELL  336
transform -1 0 3163 0 1 4294
box 0 0 6 6
use CELL  337
transform -1 0 2644 0 1 1571
box 0 0 6 6
use CELL  338
transform -1 0 1429 0 1 6171
box 0 0 6 6
use CELL  339
transform -1 0 3386 0 1 4917
box 0 0 6 6
use CELL  340
transform -1 0 1530 0 1 6171
box 0 0 6 6
use CELL  341
transform -1 0 1435 0 1 9631
box 0 0 6 6
use CELL  342
transform -1 0 1443 0 1 3699
box 0 0 6 6
use CELL  343
transform -1 0 1601 0 1 7369
box 0 0 6 6
use CELL  344
transform -1 0 1473 0 1 732
box 0 0 6 6
use CELL  345
transform -1 0 2369 0 1 1182
box 0 0 6 6
use CELL  346
transform -1 0 1435 0 1 732
box 0 0 6 6
use CELL  347
transform -1 0 1441 0 1 901
box 0 0 6 6
use CELL  348
transform -1 0 3150 0 1 3699
box 0 0 6 6
use CELL  349
transform -1 0 1529 0 1 9128
box 0 0 6 6
use CELL  350
transform -1 0 1625 0 1 7369
box 0 0 6 6
use CELL  351
transform -1 0 1663 0 1 4917
box 0 0 6 6
use CELL  352
transform -1 0 1570 0 1 10509
box 0 0 6 6
use CELL  353
transform -1 0 2921 0 1 2557
box 0 0 6 6
use CELL  354
transform -1 0 1472 0 1 10850
box 0 0 6 6
use CELL  355
transform -1 0 1440 0 1 8006
box 0 0 6 6
use CELL  356
transform -1 0 2350 0 1 1182
box 0 0 6 6
use CELL  357
transform -1 0 1595 0 1 8585
box 0 0 6 6
use CELL  358
transform -1 0 1969 0 1 901
box 0 0 6 6
use CELL  359
transform -1 0 3204 0 1 6808
box 0 0 6 6
use CELL  360
transform -1 0 1443 0 1 4917
box 0 0 6 6
use CELL  361
transform -1 0 1450 0 1 6808
box 0 0 6 6
use CELL  362
transform -1 0 3130 0 1 2557
box 0 0 6 6
use CELL  363
transform -1 0 1441 0 1 2557
box 0 0 6 6
use CELL  364
transform -1 0 2020 0 1 901
box 0 0 6 6
use CELL  365
transform -1 0 1435 0 1 901
box 0 0 6 6
use CELL  366
transform -1 0 1541 0 1 6808
box 0 0 6 6
use CELL  367
transform -1 0 1443 0 1 2028
box 0 0 6 6
use CELL  368
transform -1 0 1497 0 1 2028
box 0 0 6 6
use CELL  369
transform -1 0 2783 0 1 9631
box 0 0 6 6
use CELL  370
transform -1 0 2705 0 1 1571
box 0 0 6 6
use CELL  371
transform -1 0 2923 0 1 2028
box 0 0 6 6
use CELL  372
transform -1 0 1436 0 1 1182
box 0 0 6 6
use CELL  373
transform -1 0 3238 0 1 3126
box 0 0 6 6
use CELL  374
transform -1 0 2677 0 1 9631
box 0 0 6 6
use CELL  375
transform -1 0 1493 0 1 5572
box 0 0 6 6
use CELL  376
transform -1 0 1436 0 1 1571
box 0 0 6 6
use CELL  377
transform -1 0 2958 0 1 8585
box 0 0 6 6
use CELL  378
transform -1 0 1450 0 1 1571
box 0 0 6 6
use CELL  379
transform -1 0 1435 0 1 9128
box 0 0 6 6
use CELL  380
transform -1 0 1694 0 1 2557
box 0 0 6 6
use CELL  381
transform -1 0 3425 0 1 6171
box 0 0 6 6
use CELL  382
transform -1 0 1442 0 1 7369
box 0 0 6 6
use CELL  383
transform -1 0 1480 0 1 4294
box 0 0 6 6
use CELL  384
transform -1 0 3456 0 1 5572
box 0 0 6 6
use CELL  385
transform -1 0 2670 0 1 9631
box 0 0 6 6
use CELL  386
transform -1 0 2628 0 1 10092
box 0 0 6 6
use CELL  387
transform -1 0 1534 0 1 1571
box 0 0 6 6
use CELL  388
transform -1 0 1422 0 1 4294
box 0 0 6 6
use CELL  389
transform -1 0 1468 0 1 3126
box 0 0 6 6
use CELL  390
transform -1 0 1449 0 1 9631
box 0 0 6 6
use CELL  391
transform -1 0 1941 0 1 11105
box 0 0 6 6
use CELL  392
transform -1 0 2201 0 1 10850
box 0 0 6 6
use CELL  393
transform -1 0 2001 0 1 901
box 0 0 6 6
use CELL  394
transform -1 0 1441 0 1 11264
box 0 0 6 6
use CELL  395
transform -1 0 2655 0 1 10092
box 0 0 6 6
use CELL  396
transform -1 0 3291 0 1 6808
box 0 0 6 6
use CELL  397
transform -1 0 1553 0 1 7369
box 0 0 6 6
use CELL  398
transform -1 0 3229 0 1 6808
box 0 0 6 6
use CELL  399
transform -1 0 3149 0 1 8006
box 0 0 6 6
use CELL  400
transform -1 0 3046 0 1 8585
box 0 0 6 6
use CELL  401
transform -1 0 2713 0 1 9631
box 0 0 6 6
use CELL  402
transform -1 0 1448 0 1 732
box 0 0 6 6
use CELL  403
transform -1 0 1441 0 1 10509
box 0 0 6 6
use CELL  404
transform -1 0 1591 0 1 3126
box 0 0 6 6
use CELL  405
transform -1 0 1608 0 1 11264
box 0 0 6 6
use CELL  406
transform -1 0 2450 0 1 10509
box 0 0 6 6
use CELL  407
transform -1 0 1510 0 1 10509
box 0 0 6 6
use CELL  408
transform -1 0 1494 0 1 6171
box 0 0 6 6
use CELL  409
transform -1 0 1449 0 1 7369
box 0 0 6 6
use CELL  410
transform -1 0 2027 0 1 901
box 0 0 6 6
use CELL  411
transform -1 0 1428 0 1 9631
box 0 0 6 6
use CELL  412
transform -1 0 1536 0 1 9128
box 0 0 6 6
use CELL  413
transform -1 0 1490 0 1 2028
box 0 0 6 6
use CELL  414
transform -1 0 1450 0 1 6171
box 0 0 6 6
use CELL  415
transform -1 0 1519 0 1 4294
box 0 0 6 6
use CELL  416
transform -1 0 1448 0 1 10509
box 0 0 6 6
use CELL  417
transform -1 0 1891 0 1 5572
box 0 0 6 6
use CELL  418
transform -1 0 1494 0 1 11105
box 0 0 6 6
use CELL  419
transform -1 0 1450 0 1 1182
box 0 0 6 6
use CELL  420
transform -1 0 1493 0 1 3126
box 0 0 6 6
use CELL  421
transform -1 0 1428 0 1 10092
box 0 0 6 6
use CELL  422
transform -1 0 1443 0 1 4294
box 0 0 6 6
use CELL  423
transform -1 0 1449 0 1 9128
box 0 0 6 6
use CELL  424
transform -1 0 1531 0 1 5572
box 0 0 6 6
use CELL  425
transform -1 0 3329 0 1 7369
box 0 0 6 6
use CELL  426
transform -1 0 1634 0 1 732
box 0 0 6 6
use CELL  427
transform -1 0 2842 0 1 2028
box 0 0 6 6
use CELL  428
transform -1 0 1429 0 1 1182
box 0 0 6 6
use CELL  429
transform -1 0 1461 0 1 10092
box 0 0 6 6
use CELL  430
transform -1 0 1422 0 1 4917
box 0 0 6 6
use CELL  431
transform -1 0 1422 0 1 6171
box 0 0 6 6
use CELL  432
transform -1 0 1474 0 1 6808
box 0 0 6 6
use CELL  433
transform -1 0 1443 0 1 1571
box 0 0 6 6
use CELL  434
transform -1 0 1463 0 1 9128
box 0 0 6 6
use CELL  435
transform -1 0 1428 0 1 901
box 0 0 6 6
use CELL  436
transform -1 0 1539 0 1 10850
box 0 0 6 6
use CELL  437
transform -1 0 3328 0 1 4917
box 0 0 6 6
use CELL  438
transform -1 0 1456 0 1 7369
box 0 0 6 6
use CELL  439
transform -1 0 3187 0 1 3126
box 0 0 6 6
use CELL  440
transform -1 0 2181 0 1 10850
box 0 0 6 6
use CELL  441
transform -1 0 1505 0 1 3699
box 0 0 6 6
use CELL  442
transform -1 0 2422 0 1 10509
box 0 0 6 6
use CELL  443
transform -1 0 1487 0 1 7369
box 0 0 6 6
use CELL  444
transform -1 0 1476 0 1 1182
box 0 0 6 6
use CELL  445
transform -1 0 1422 0 1 3126
box 0 0 6 6
use CELL  446
transform -1 0 1613 0 1 10092
box 0 0 6 6
use CELL  447
transform -1 0 3407 0 1 6171
box 0 0 6 6
use CELL  448
transform -1 0 3300 0 1 4294
box 0 0 6 6
use CELL  449
transform -1 0 1522 0 1 8006
box 0 0 6 6
use CELL  450
transform -1 0 3264 0 1 7369
box 0 0 6 6
use CELL  451
transform -1 0 1473 0 1 3699
box 0 0 6 6
use CELL  452
transform -1 0 1519 0 1 4917
box 0 0 6 6
use CELL  453
transform -1 0 1434 0 1 10509
box 0 0 6 6
use CELL  454
transform -1 0 3400 0 1 4917
box 0 0 6 6
use CELL  455
transform -1 0 2780 0 1 2028
box 0 0 6 6
use CELL  456
transform -1 0 1494 0 1 11264
box 0 0 6 6
use CELL  457
transform -1 0 1422 0 1 3699
box 0 0 6 6
use CELL  458
transform -1 0 1449 0 1 8585
box 0 0 6 6
use CELL  459
transform -1 0 2224 0 1 10509
box 0 0 6 6
use CELL  460
transform -1 0 2426 0 1 1182
box 0 0 6 6
use CELL  461
transform -1 0 1495 0 1 1182
box 0 0 6 6
use CELL  462
transform -1 0 1435 0 1 10092
box 0 0 6 6
use CELL  463
transform -1 0 1455 0 1 11264
box 0 0 6 6
use CELL  464
transform -1 0 2621 0 1 10092
box 0 0 6 6
use CELL  465
transform -1 0 2857 0 1 9128
box 0 0 6 6
use CELL  466
transform -1 0 2713 0 1 2028
box 0 0 6 6
use CELL  467
transform -1 0 2145 0 1 10850
box 0 0 6 6
use CELL  468
transform -1 0 3207 0 1 3699
box 0 0 6 6
use CELL  469
transform -1 0 1422 0 1 6808
box 0 0 6 6
use CELL  470
transform -1 0 3363 0 1 6171
box 0 0 6 6
use CELL  471
transform -1 0 2103 0 1 10850
box 0 0 6 6
use CELL  472
transform -1 0 1429 0 1 4294
box 0 0 6 6
use CELL  473
transform -1 0 1475 0 1 9128
box 0 0 6 6
use CELL  474
transform -1 0 1867 0 1 11105
box 0 0 6 6
use CELL  475
transform -1 0 3309 0 1 4917
box 0 0 6 6
use CELL  476
transform -1 0 2376 0 1 1182
box 0 0 6 6
use CELL  477
transform -1 0 3470 0 1 5572
box 0 0 6 6
use CELL  478
transform -1 0 3191 0 1 7369
box 0 0 6 6
use CELL  479
transform -1 0 1449 0 1 10092
box 0 0 6 6
use CELL  480
transform -1 0 2909 0 1 2028
box 0 0 6 6
use CELL  481
transform -1 0 3189 0 1 8006
box 0 0 6 6
use CELL  482
transform -1 0 1634 0 1 11264
box 0 0 6 6
use CELL  483
transform -1 0 1471 0 1 1571
box 0 0 6 6
use CELL  484
transform -1 0 1475 0 1 8585
box 0 0 6 6
use CELL  485
transform -1 0 2977 0 1 9128
box 0 0 6 6
use CELL  486
transform -1 0 1435 0 1 11105
box 0 0 6 6
use CELL  487
transform -1 0 1491 0 1 10509
box 0 0 6 6
use CELL  488
transform -1 0 2963 0 1 9128
box 0 0 6 6
use CELL  489
transform -1 0 3278 0 1 7369
box 0 0 6 6
use CELL  490
transform -1 0 1434 0 1 2557
box 0 0 6 6
use CELL  491
transform -1 0 3453 0 1 6171
box 0 0 6 6
use CELL  492
transform -1 0 3463 0 1 5572
box 0 0 6 6
use CELL  493
transform -1 0 3078 0 1 3699
box 0 0 6 6
use CELL  494
transform -1 0 1428 0 1 732
box 0 0 6 6
use CELL  495
transform -1 0 1448 0 1 2557
box 0 0 6 6
use CELL  496
transform -1 0 3236 0 1 4294
box 0 0 6 6
use CELL  497
transform -1 0 2773 0 1 2028
box 0 0 6 6
use CELL  498
transform -1 0 2188 0 1 10850
box 0 0 6 6
use CELL  499
transform -1 0 1518 0 1 6171
box 0 0 6 6
use CELL  500
transform -1 0 2207 0 1 10850
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 1922 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 1887 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 2343 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 2366 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 2354 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 2234 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 2065 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 1941 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 1771 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 1505 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 1505 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 1511 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 1511 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 1505 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 1503 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 1511 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 2222 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 2590 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 2878 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 2301 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 2026 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 2230 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 1936 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 1924 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 2018 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 2000 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 2276 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 2270 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 2253 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 1845 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 1862 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 1981 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 1449 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 1449 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 1449 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 1455 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 1456 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 2176 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 1455 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 1455 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 1455 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 1461 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 1462 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 1456 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 1462 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 1449 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 1461 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 1461 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 1461 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 1467 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 1468 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 1462 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 1468 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 2399 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 2491 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 2377 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 2320 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 1906 0 1 901
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 1605 0 1 732
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 1592 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 1594 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 1558 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 1610 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 2440 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 2445 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 2926 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 2920 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 3106 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 3112 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 1606 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 1576 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 2323 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 2982 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 2881 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 2695 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 2591 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 2398 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 2157 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 1903 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 3119 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 3234 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 3192 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 3320 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 3368 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 3272 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 3193 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 2985 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 2884 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 2698 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 2163 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 2313 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 2330 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 2312 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 2024 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 2306 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 2332 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 2356 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 2278 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 2080 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 2373 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 2362 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 2333 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 2203 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 1898 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 1499 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 1493 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 1479 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 1499 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-109
transform 1 0 1493 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-110
transform 1 0 1500 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-111
transform 1 0 1499 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-112
transform 1 0 1493 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-113
transform 1 0 1493 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-114
transform 1 0 1493 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-115
transform 1 0 1481 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-116
transform 1 0 1499 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-117
transform 1 0 1486 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-118
transform 1 0 2041 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-119
transform 1 0 1734 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-120
transform 1 0 1455 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-121
transform 1 0 1455 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-122
transform 1 0 2245 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-123
transform 1 0 2375 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-124
transform 1 0 2386 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-125
transform 1 0 1546 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-126
transform 1 0 1520 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-127
transform 1 0 2155 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-128
transform 1 0 1570 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-129
transform 1 0 1556 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-130
transform 1 0 1549 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-131
transform 1 0 2403 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-132
transform 1 0 2104 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-133
transform 1 0 2326 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-134
transform 1 0 2686 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-135
transform 1 0 2890 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-136
transform 1 0 3090 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-137
transform 1 0 3200 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-138
transform 1 0 3163 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-139
transform 1 0 3242 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-140
transform 1 0 2689 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-141
transform 1 0 2893 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-142
transform 1 0 3093 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-143
transform 1 0 3203 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-144
transform 1 0 3166 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-145
transform 1 0 3245 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-146
transform 1 0 3316 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-147
transform 1 0 3412 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-148
transform 1 0 3370 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-149
transform 1 0 3229 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-150
transform 1 0 3278 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-151
transform 1 0 3156 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-152
transform 1 0 3013 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-153
transform 1 0 2906 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-154
transform 1 0 2720 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-155
transform 1 0 2674 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-156
transform 1 0 2872 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-157
transform 1 0 3078 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-158
transform 1 0 1510 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-159
transform 1 0 1905 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-160
transform 1 0 1507 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-161
transform 1 0 1497 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-162
transform 1 0 1951 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-163
transform 1 0 2132 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-164
transform 1 0 2415 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-165
transform 1 0 2031 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-166
transform 1 0 2360 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-167
transform 1 0 2360 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-168
transform 1 0 2768 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-169
transform 1 0 2336 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-170
transform 1 0 2800 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-171
transform 1 0 3022 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-172
transform 1 0 2428 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-173
transform 1 0 2842 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-174
transform 1 0 1503 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-175
transform 1 0 1540 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-176
transform 1 0 1553 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-177
transform 1 0 1554 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-178
transform 1 0 1542 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-179
transform 1 0 1565 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-180
transform 1 0 1570 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-181
transform 1 0 1509 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-182
transform 1 0 3240 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-183
transform 1 0 3344 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-184
transform 1 0 3386 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-185
transform 1 0 3290 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-186
transform 1 0 3347 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-187
transform 1 0 3389 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-188
transform 1 0 3293 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-189
transform 1 0 3199 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-190
transform 1 0 3120 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-191
transform 1 0 3157 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-192
transform 1 0 3017 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-193
transform 1 0 2219 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-194
transform 1 0 2488 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-195
transform 1 0 2679 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-196
transform 1 0 2771 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-197
transform 1 0 2222 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-198
transform 1 0 2491 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-199
transform 1 0 2682 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-200
transform 1 0 2476 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-201
transform 1 0 2667 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-202
transform 1 0 2774 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-203
transform 1 0 2951 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-204
transform 1 0 3058 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-205
transform 1 0 2470 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-206
transform 1 0 2661 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-207
transform 1 0 2759 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-208
transform 1 0 2954 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-209
transform 1 0 3061 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-210
transform 1 0 3195 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-211
transform 1 0 3310 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-212
transform 1 0 2662 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-213
transform 1 0 2860 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-214
transform 1 0 3047 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-215
transform 1 0 2665 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-216
transform 1 0 2863 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-217
transform 1 0 3050 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-218
transform 1 0 3175 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-219
transform 1 0 2400 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-220
transform 1 0 2650 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-221
transform 1 0 2848 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-222
transform 1 0 3035 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-223
transform 1 0 3178 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-224
transform 1 0 3138 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-225
transform 1 0 3217 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-226
transform 1 0 2403 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-227
transform 1 0 2644 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-228
transform 1 0 2842 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-229
transform 1 0 3029 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-230
transform 1 0 3353 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-231
transform 1 0 3260 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-232
transform 1 0 3181 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-233
transform 1 0 3212 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-234
transform 1 0 3072 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-235
transform 1 0 3356 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-236
transform 1 0 3263 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-237
transform 1 0 3184 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-238
transform 1 0 3215 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-239
transform 1 0 3075 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-240
transform 1 0 2878 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-241
transform 1 0 3341 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-242
transform 1 0 3437 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-243
transform 1 0 3413 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-244
transform 1 0 3279 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-245
transform 1 0 3335 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-246
transform 1 0 3440 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-247
transform 1 0 3416 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-248
transform 1 0 3282 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-249
transform 1 0 3313 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-250
transform 1 0 3198 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-251
transform 1 0 3046 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-252
transform 1 0 2939 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-253
transform 1 0 2753 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-254
transform 1 0 2655 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-255
transform 1 0 2464 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-256
transform 1 0 2207 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-257
transform 1 0 3388 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-258
transform 1 0 3391 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-259
transform 1 0 3254 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-260
transform 1 0 3376 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-261
transform 1 0 3257 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-262
transform 1 0 3137 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-263
transform 1 0 3252 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-264
transform 1 0 3210 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-265
transform 1 0 3338 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-266
transform 1 0 2994 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-267
transform 1 0 2887 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-268
transform 1 0 2701 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-269
transform 1 0 2609 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-270
transform 1 0 2410 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-271
transform 1 0 3255 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-272
transform 1 0 3213 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-273
transform 1 0 3341 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-274
transform 1 0 3380 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-275
transform 1 0 3284 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-276
transform 1 0 3205 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-277
transform 1 0 3126 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-278
transform 1 0 3140 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-279
transform 1 0 2997 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-280
transform 1 0 2912 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-281
transform 1 0 2894 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-282
transform 1 0 3010 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-283
transform 1 0 3034 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-284
transform 1 0 2356 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-285
transform 1 0 2896 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-286
transform 1 0 1651 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-287
transform 1 0 1657 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-288
transform 1 0 1603 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-289
transform 1 0 2816 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-290
transform 1 0 3005 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-291
transform 1 0 3145 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-292
transform 1 0 3108 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-293
transform 1 0 3196 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-294
transform 1 0 3275 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-295
transform 1 0 3371 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-296
transform 1 0 3323 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-297
transform 1 0 3195 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-298
transform 1 0 3237 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-299
transform 1 0 3122 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-300
transform 1 0 2970 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-301
transform 1 0 2869 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-302
transform 1 0 2677 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-303
transform 1 0 2594 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-304
transform 1 0 2401 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-305
transform 1 0 2600 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-306
transform 1 0 2819 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-307
transform 1 0 3008 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-308
transform 1 0 3148 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-309
transform 1 0 3111 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-310
transform 1 0 2603 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-311
transform 1 0 2780 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-312
transform 1 0 2969 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-313
transform 1 0 3109 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-314
transform 1 0 3078 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-315
transform 1 0 3163 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-316
transform 1 0 3242 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-317
transform 1 0 3332 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-318
transform 1 0 3284 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-319
transform 1 0 3168 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-320
transform 1 0 3198 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-321
transform 1 0 3083 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-322
transform 1 0 2958 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-323
transform 1 0 2857 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-324
transform 1 0 2618 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-325
transform 1 0 2810 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-326
transform 1 0 2999 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-327
transform 1 0 3139 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-328
transform 1 0 3129 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-329
transform 1 0 3208 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-330
transform 1 0 3287 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-331
transform 1 0 3383 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-332
transform 1 0 3314 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-333
transform 1 0 3186 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-334
transform 1 0 3228 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-335
transform 1 0 3113 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-336
transform 1 0 2621 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-337
transform 1 0 2813 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-338
transform 1 0 3002 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-339
transform 1 0 3142 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-340
transform 1 0 3096 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-341
transform 1 0 3181 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-342
transform 1 0 3260 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-343
transform 1 0 3356 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-344
transform 1 0 3308 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-345
transform 1 0 3180 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-346
transform 1 0 3222 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-347
transform 1 0 3107 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-348
transform 1 0 2382 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-349
transform 1 0 2385 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-350
transform 1 0 2606 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-351
transform 1 0 2798 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-352
transform 1 0 2987 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-353
transform 1 0 3127 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-354
transform 1 0 2832 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-355
transform 1 0 2652 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-356
transform 1 0 2933 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-357
transform 1 0 3062 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-358
transform 1 0 3173 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-359
transform 1 0 3143 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-360
transform 1 0 3259 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-361
transform 1 0 3307 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-362
transform 1 0 3211 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-363
transform 1 0 2936 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-364
transform 1 0 2835 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-365
transform 1 0 2655 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-366
transform 1 0 2555 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-367
transform 1 0 2308 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-368
transform 1 0 1971 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-369
transform 1 0 1882 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-370
transform 1 0 3059 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-371
transform 1 0 3176 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-372
transform 1 0 3146 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-373
transform 1 0 3262 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-374
transform 1 0 3310 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-375
transform 1 0 3214 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-376
transform 1 0 3103 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-377
transform 1 0 3018 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-378
transform 1 0 3055 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-379
transform 1 0 2879 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-380
transform 1 0 2743 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-381
transform 1 0 2545 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-382
transform 1 0 2338 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-383
transform 1 0 1951 0 1 901
box 0 0 3 6
use FEEDTHRU  F-384
transform 1 0 2249 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-385
transform 1 0 2284 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-386
transform 1 0 2193 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-387
transform 1 0 2023 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-388
transform 1 0 2011 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-389
transform 1 0 1633 0 1 901
box 0 0 3 6
use FEEDTHRU  F-390
transform 1 0 2125 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-391
transform 1 0 1514 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-392
transform 1 0 1513 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-393
transform 1 0 1518 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-394
transform 1 0 1573 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-395
transform 1 0 1555 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-396
transform 1 0 2824 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-397
transform 1 0 2806 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-398
transform 1 0 1596 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-399
transform 1 0 1591 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-400
transform 1 0 1561 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-401
transform 1 0 1597 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-402
transform 1 0 1627 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-403
transform 1 0 1567 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-404
transform 1 0 1574 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-405
transform 1 0 1576 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-406
transform 1 0 1546 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-407
transform 1 0 1921 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-408
transform 1 0 1735 0 1 901
box 0 0 3 6
use FEEDTHRU  F-409
transform 1 0 2228 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-410
transform 1 0 2234 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-411
transform 1 0 1970 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-412
transform 1 0 1904 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-413
transform 1 0 1918 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-414
transform 1 0 2187 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-415
transform 1 0 1851 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-416
transform 1 0 1886 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-417
transform 1 0 1491 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-418
transform 1 0 1487 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-419
transform 1 0 1493 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-420
transform 1 0 1493 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-421
transform 1 0 1480 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-422
transform 1 0 2029 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-423
transform 1 0 2374 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-424
transform 1 0 2488 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-425
transform 1 0 2281 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-426
transform 1 0 2275 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-427
transform 1 0 1594 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-428
transform 1 0 1636 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-429
transform 1 0 1652 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-430
transform 1 0 1663 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-431
transform 1 0 1662 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-432
transform 1 0 1627 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-433
transform 1 0 1651 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-434
transform 1 0 1669 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-435
transform 1 0 1747 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-436
transform 1 0 3014 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-437
transform 1 0 3008 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-438
transform 1 0 2834 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-439
transform 1 0 2732 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-440
transform 1 0 1530 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-441
transform 1 0 1525 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-442
transform 1 0 1544 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-443
transform 1 0 1564 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-444
transform 1 0 2077 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-445
transform 1 0 1554 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-446
transform 1 0 1555 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-447
transform 1 0 1543 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-448
transform 1 0 1543 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-449
transform 1 0 1549 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-450
transform 1 0 1517 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-451
transform 1 0 1523 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-452
transform 1 0 1572 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-453
transform 1 0 1522 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-454
transform 1 0 1517 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-455
transform 1 0 1517 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-456
transform 1 0 1517 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-457
transform 1 0 1529 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-458
transform 1 0 1535 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-459
transform 1 0 1523 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-460
transform 1 0 1555 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-461
transform 1 0 1561 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-462
transform 1 0 1549 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-463
transform 1 0 2374 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-464
transform 1 0 2368 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-465
transform 1 0 2573 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-466
transform 1 0 2658 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-467
transform 1 0 2838 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-468
transform 1 0 2939 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-469
transform 1 0 3071 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-470
transform 1 0 3179 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-471
transform 1 0 3149 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-472
transform 1 0 3265 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-473
transform 1 0 3313 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-474
transform 1 0 3217 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-475
transform 1 0 3145 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-476
transform 1 0 3054 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-477
transform 1 0 3085 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-478
transform 1 0 2945 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-479
transform 1 0 2755 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-480
transform 1 0 2563 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-481
transform 1 0 2326 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-482
transform 1 0 2344 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-483
transform 1 0 2320 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-484
transform 1 0 2160 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-485
transform 1 0 3281 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-486
transform 1 0 3159 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-487
transform 1 0 3016 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-488
transform 1 0 2909 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-489
transform 1 0 2723 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-490
transform 1 0 2597 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-491
transform 1 0 2380 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-492
transform 1 0 2169 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-493
transform 1 0 1922 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-494
transform 1 0 3204 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-495
transform 1 0 3095 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-496
transform 1 0 3373 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-497
transform 1 0 3415 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-498
transform 1 0 3290 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-499
transform 1 0 3338 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-500
transform 1 0 3319 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-501
transform 1 0 3175 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-502
transform 1 0 3090 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-503
transform 1 0 3121 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-504
transform 1 0 2981 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-505
transform 1 0 2786 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-506
transform 1 0 2594 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-507
transform 1 0 2357 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-508
transform 1 0 2008 0 1 901
box 0 0 3 6
use FEEDTHRU  F-509
transform 1 0 1641 0 1 732
box 0 0 3 6
use FEEDTHRU  F-510
transform 1 0 1488 0 1 11321
box 0 0 3 6
use FEEDTHRU  F-511
transform 1 0 1584 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-512
transform 1 0 1573 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-513
transform 1 0 1491 0 1 11321
box 0 0 3 6
use FEEDTHRU  F-514
transform 1 0 1587 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-515
transform 1 0 1576 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-516
transform 1 0 1953 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-517
transform 1 0 2077 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-518
transform 1 0 2426 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-519
transform 1 0 2469 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-520
transform 1 0 2355 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-521
transform 1 0 2318 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-522
transform 1 0 1533 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-523
transform 1 0 1518 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-524
transform 1 0 1513 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-525
transform 1 0 1551 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-526
transform 1 0 3289 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-527
transform 1 0 3247 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-528
transform 1 0 3131 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-529
transform 1 0 3161 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-530
transform 1 0 3053 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-531
transform 1 0 3283 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-532
transform 1 0 3241 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-533
transform 1 0 3169 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-534
transform 1 0 3277 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-535
transform 1 0 3235 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-536
transform 1 0 3125 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-537
transform 1 0 2331 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-538
transform 1 0 2547 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-539
transform 1 0 2453 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-540
transform 1 0 1626 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-541
transform 1 0 2520 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-542
transform 1 0 1650 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-543
transform 1 0 2544 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-544
transform 1 0 1621 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-545
transform 1 0 1633 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-546
transform 1 0 1639 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-547
transform 1 0 2426 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-548
transform 1 0 2390 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-549
transform 1 0 2336 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-550
transform 1 0 2348 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-551
transform 1 0 2325 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-552
transform 1 0 2211 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-553
transform 1 0 1627 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-554
transform 1 0 1639 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-555
transform 1 0 1609 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-556
transform 1 0 1633 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-557
transform 1 0 1645 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-558
transform 1 0 1645 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-559
transform 1 0 1595 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-560
transform 1 0 1607 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-561
transform 1 0 1588 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-562
transform 1 0 1583 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-563
transform 1 0 1596 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-564
transform 1 0 1614 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-565
transform 1 0 1591 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-566
transform 1 0 1586 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-567
transform 1 0 2288 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-568
transform 1 0 2042 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-569
transform 1 0 2090 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-570
transform 1 0 1966 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-571
transform 1 0 2276 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-572
transform 1 0 2259 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-573
transform 1 0 1571 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-574
transform 1 0 1559 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-575
transform 1 0 1609 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-576
transform 1 0 1552 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-577
transform 1 0 1547 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-578
transform 1 0 1572 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-579
transform 1 0 1888 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-580
transform 1 0 1876 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-581
transform 1 0 1567 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-582
transform 1 0 1886 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-583
transform 1 0 1958 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-584
transform 1 0 2282 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-585
transform 1 0 2288 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-586
transform 1 0 1555 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-587
transform 1 0 2796 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-588
transform 1 0 2891 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-589
transform 1 0 2891 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-590
transform 1 0 3155 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-591
transform 1 0 3077 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-592
transform 1 0 3205 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-593
transform 1 0 3217 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-594
transform 1 0 2995 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-595
transform 1 0 2941 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-596
transform 1 0 2894 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-597
transform 1 0 2894 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-598
transform 1 0 3158 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-599
transform 1 0 2799 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-600
transform 1 0 2610 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-601
transform 1 0 2525 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-602
transform 1 0 2500 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-603
transform 1 0 2459 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-604
transform 1 0 2323 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-605
transform 1 0 2197 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-606
transform 1 0 2215 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-607
transform 1 0 1819 0 1 901
box 0 0 3 6
use FEEDTHRU  F-608
transform 1 0 1593 0 1 732
box 0 0 3 6
use FEEDTHRU  F-609
transform 1 0 1615 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-610
transform 1 0 1906 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-611
transform 1 0 2290 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-612
transform 1 0 2062 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-613
transform 1 0 2409 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-614
transform 1 0 2374 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-615
transform 1 0 2339 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-616
transform 1 0 1591 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-617
transform 1 0 2173 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-618
transform 1 0 1516 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-619
transform 1 0 2315 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-620
transform 1 0 2350 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-621
transform 1 0 2205 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-622
transform 1 0 1960 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-623
transform 1 0 2146 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-624
transform 1 0 1579 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-625
transform 1 0 2059 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-626
transform 1 0 1522 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-627
transform 1 0 1498 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-628
transform 1 0 1528 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-629
transform 1 0 1532 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-630
transform 1 0 1537 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-631
transform 1 0 1542 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-632
transform 1 0 1543 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-633
transform 1 0 1573 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-634
transform 1 0 1585 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-635
transform 1 0 1579 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-636
transform 1 0 1541 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-637
transform 1 0 1553 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-638
transform 1 0 3020 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-639
transform 1 0 3160 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-640
transform 1 0 3123 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-641
transform 1 0 2761 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-642
transform 1 0 2951 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-643
transform 1 0 3091 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-644
transform 1 0 3060 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-645
transform 1 0 3202 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-646
transform 1 0 3223 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-647
transform 1 0 3295 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-648
transform 1 0 2569 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-649
transform 1 0 2332 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-650
transform 1 0 1976 0 1 901
box 0 0 3 6
use FEEDTHRU  F-651
transform 1 0 1663 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-652
transform 1 0 1735 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-653
transform 1 0 1795 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-654
transform 1 0 1715 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-655
transform 1 0 1709 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-656
transform 1 0 2366 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-657
transform 1 0 1679 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-658
transform 1 0 1651 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-659
transform 1 0 2433 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-660
transform 1 0 2494 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-661
transform 1 0 2435 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-662
transform 1 0 1693 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-663
transform 1 0 1687 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-664
transform 1 0 1753 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-665
transform 1 0 1656 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-666
transform 1 0 1651 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-667
transform 1 0 1622 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-668
transform 1 0 2317 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-669
transform 1 0 1553 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-670
transform 1 0 1591 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-671
transform 1 0 1603 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-672
transform 1 0 1591 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-673
transform 1 0 1561 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-674
transform 1 0 1560 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-675
transform 1 0 1555 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-676
transform 1 0 1565 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-677
transform 1 0 1546 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-678
transform 1 0 1597 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-679
transform 1 0 1609 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-680
transform 1 0 1597 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-681
transform 1 0 1567 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-682
transform 1 0 1566 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-683
transform 1 0 1561 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-684
transform 1 0 1550 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-685
transform 1 0 1540 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-686
transform 1 0 1504 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-687
transform 1 0 1603 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-688
transform 1 0 1609 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-689
transform 1 0 1621 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-690
transform 1 0 1615 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-691
transform 1 0 1565 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-692
transform 1 0 1577 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-693
transform 1 0 1558 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-694
transform 1 0 1553 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-695
transform 1 0 1560 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-696
transform 1 0 1536 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-697
transform 1 0 1579 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-698
transform 1 0 1578 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-699
transform 1 0 1573 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-700
transform 1 0 1562 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-701
transform 1 0 2161 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-702
transform 1 0 2065 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-703
transform 1 0 1584 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-704
transform 1 0 1579 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-705
transform 1 0 1568 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-706
transform 1 0 1558 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-707
transform 1 0 1522 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-708
transform 1 0 1675 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-709
transform 1 0 1681 0 1 901
box 0 0 3 6
use FEEDTHRU  F-710
transform 1 0 1585 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-711
transform 1 0 1615 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-712
transform 1 0 1627 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-713
transform 1 0 1621 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-714
transform 1 0 1571 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-715
transform 1 0 1583 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-716
transform 1 0 1564 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-717
transform 1 0 1559 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-718
transform 1 0 1566 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-719
transform 1 0 1542 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-720
transform 1 0 1498 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-721
transform 1 0 1479 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-722
transform 1 0 1699 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-723
transform 1 0 3103 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-724
transform 1 0 3109 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-725
transform 1 0 3011 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-726
transform 1 0 3005 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-727
transform 1 0 1649 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-728
transform 1 0 2923 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-729
transform 1 0 1819 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-730
transform 1 0 3049 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-731
transform 1 0 3037 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-732
transform 1 0 2957 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-733
transform 1 0 2999 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-734
transform 1 0 1643 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-735
transform 1 0 2729 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-736
transform 1 0 1728 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-737
transform 1 0 2538 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-738
transform 1 0 2456 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-739
transform 1 0 1764 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-740
transform 1 0 1765 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-741
transform 1 0 1676 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-742
transform 1 0 1774 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-743
transform 1 0 1600 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-744
transform 1 0 3005 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-745
transform 1 0 3149 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-746
transform 1 0 3119 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-747
transform 1 0 3229 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-748
transform 1 0 3271 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-749
transform 1 0 3152 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-750
transform 1 0 3122 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-751
transform 1 0 3232 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-752
transform 1 0 3274 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-753
transform 1 0 3193 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-754
transform 1 0 3109 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-755
transform 1 0 3036 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-756
transform 1 0 1582 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-757
transform 1 0 1513 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-758
transform 1 0 1504 0 1 901
box 0 0 3 6
use FEEDTHRU  F-759
transform 1 0 1596 0 1 732
box 0 0 3 6
use FEEDTHRU  F-760
transform 1 0 1624 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-761
transform 1 0 1640 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-762
transform 1 0 1588 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-763
transform 1 0 1630 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-764
transform 1 0 1646 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-765
transform 1 0 1657 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-766
transform 1 0 1519 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-767
transform 1 0 1522 0 1 901
box 0 0 3 6
use FEEDTHRU  F-768
transform 1 0 1581 0 1 732
box 0 0 3 6
use FEEDTHRU  F-769
transform 1 0 1613 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-770
transform 1 0 1663 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-771
transform 1 0 1675 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-772
transform 1 0 1625 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-773
transform 1 0 1613 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-774
transform 1 0 1601 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-775
transform 1 0 1608 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-776
transform 1 0 1632 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-777
transform 1 0 1699 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-778
transform 1 0 1729 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-779
transform 1 0 2320 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-780
transform 1 0 2098 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-781
transform 1 0 2439 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-782
transform 1 0 2404 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-783
transform 1 0 2369 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-784
transform 1 0 1643 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-785
transform 1 0 1661 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-786
transform 1 0 1625 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-787
transform 1 0 1602 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-788
transform 1 0 1603 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-789
transform 1 0 1639 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-790
transform 1 0 1651 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-791
transform 1 0 1603 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-792
transform 1 0 1598 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-793
transform 1 0 1582 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-794
transform 1 0 2558 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-795
transform 1 0 2604 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-796
transform 1 0 2724 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-797
transform 1 0 2861 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-798
transform 1 0 2873 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-799
transform 1 0 3095 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-800
transform 1 0 3065 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-801
transform 1 0 3169 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-802
transform 1 0 3211 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-803
transform 1 0 3163 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-804
transform 1 0 3106 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-805
transform 1 0 3021 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-806
transform 1 0 3058 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-807
transform 1 0 2882 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-808
transform 1 0 2746 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-809
transform 1 0 2548 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-810
transform 1 0 2507 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-811
transform 1 0 2311 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-812
transform 1 0 1935 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-813
transform 1 0 1885 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-814
transform 1 0 1578 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-815
transform 1 0 2501 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-816
transform 1 0 2230 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-817
transform 1 0 1653 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-818
transform 1 0 2566 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-819
transform 1 0 2180 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-820
transform 1 0 2192 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-821
transform 1 0 2294 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-822
transform 1 0 2336 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-823
transform 1 0 2307 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-824
transform 1 0 2199 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-825
transform 1 0 1850 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-826
transform 1 0 1957 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-827
transform 1 0 2572 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-828
transform 1 0 2158 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-829
transform 1 0 2002 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-830
transform 1 0 1632 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-831
transform 1 0 1633 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-832
transform 1 0 1628 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-833
transform 1 0 1612 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-834
transform 1 0 1570 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-835
transform 1 0 1675 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-836
transform 1 0 1639 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-837
transform 1 0 1638 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-838
transform 1 0 1639 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-839
transform 1 0 1687 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-840
transform 1 0 1675 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-841
transform 1 0 3133 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-842
transform 1 0 3042 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-843
transform 1 0 3079 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-844
transform 1 0 2921 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-845
transform 1 0 2764 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-846
transform 1 0 3127 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-847
transform 1 0 3121 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-848
transform 1 0 3205 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-849
transform 1 0 3265 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-850
transform 1 0 3223 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-851
transform 1 0 3113 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-852
transform 1 0 3243 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-853
transform 1 0 3011 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-854
transform 1 0 2897 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-855
transform 1 0 2383 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-856
transform 1 0 2600 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-857
transform 1 0 2356 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-858
transform 1 0 2172 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-859
transform 1 0 2350 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-860
transform 1 0 2145 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-861
transform 1 0 1925 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-862
transform 1 0 2524 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-863
transform 1 0 2341 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-864
transform 1 0 2518 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-865
transform 1 0 2674 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-866
transform 1 0 2834 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-867
transform 1 0 3025 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-868
transform 1 0 3000 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-869
transform 1 0 3067 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-870
transform 1 0 3151 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-871
transform 1 0 3199 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-872
transform 1 0 3163 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-873
transform 1 0 3059 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-874
transform 1 0 3089 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-875
transform 1 0 1715 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-876
transform 1 0 2777 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-877
transform 1 0 2706 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-878
transform 1 0 2598 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-879
transform 1 0 2495 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-880
transform 1 0 2296 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-881
transform 1 0 2512 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-882
transform 1 0 2668 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-883
transform 1 0 1760 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-884
transform 1 0 2989 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-885
transform 1 0 2952 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-886
transform 1 0 3013 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-887
transform 1 0 3031 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-888
transform 1 0 3145 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-889
transform 1 0 3151 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-890
transform 1 0 3053 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-891
transform 1 0 3059 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-892
transform 1 0 2814 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-893
transform 1 0 2634 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-894
transform 1 0 2531 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-895
transform 1 0 2332 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-896
transform 1 0 2127 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-897
transform 1 0 1888 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-898
transform 1 0 2915 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-899
transform 1 0 3032 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-900
transform 1 0 3029 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-901
transform 1 0 3137 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-902
transform 1 0 3107 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-903
transform 1 0 3217 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-904
transform 1 0 3259 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-905
transform 1 0 3199 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-906
transform 1 0 3220 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-907
transform 1 0 3049 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-908
transform 1 0 2873 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-909
transform 1 0 2701 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-910
transform 1 0 3012 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-911
transform 1 0 3079 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-912
transform 1 0 3043 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-913
transform 1 0 1885 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-914
transform 1 0 1642 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-915
transform 1 0 1658 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-916
transform 1 0 1669 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-917
transform 1 0 1668 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-918
transform 1 0 1717 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-919
transform 1 0 1705 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-920
transform 1 0 2947 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-921
transform 1 0 2236 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-922
transform 1 0 1630 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-923
transform 1 0 1660 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-924
transform 1 0 1664 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-925
transform 1 0 1681 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-926
transform 1 0 1680 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-927
transform 1 0 1831 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-928
transform 1 0 1711 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-929
transform 1 0 3001 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-930
transform 1 0 3007 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-931
transform 1 0 2909 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-932
transform 1 0 2891 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-933
transform 1 0 1679 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-934
transform 1 0 1709 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-935
transform 1 0 1698 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-936
transform 1 0 2239 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-937
transform 1 0 1612 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-938
transform 1 0 1648 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-939
transform 1 0 1670 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-940
transform 1 0 1759 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-941
transform 1 0 1758 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-942
transform 1 0 2893 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-943
transform 1 0 1795 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-944
transform 1 0 3031 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-945
transform 1 0 2965 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-946
transform 1 0 2867 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-947
transform 1 0 2267 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-948
transform 1 0 1655 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-949
transform 1 0 1691 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-950
transform 1 0 3145 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-951
transform 1 0 3193 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-952
transform 1 0 3196 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-953
transform 1 0 3112 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-954
transform 1 0 3039 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-955
transform 1 0 3001 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-956
transform 1 0 2507 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-957
transform 1 0 2662 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-958
transform 1 0 2494 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-959
transform 1 0 2287 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-960
transform 1 0 3139 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-961
transform 1 0 3187 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-962
transform 1 0 3127 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-963
transform 1 0 3049 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-964
transform 1 0 2964 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-965
transform 1 0 3163 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-966
transform 1 0 3121 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-967
transform 1 0 3019 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-968
transform 1 0 3115 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-969
transform 1 0 3017 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-970
transform 1 0 3053 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-971
transform 1 0 3008 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-972
transform 1 0 2251 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-973
transform 1 0 2254 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-974
transform 1 0 2203 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-975
transform 1 0 2269 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-976
transform 1 0 2363 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-977
transform 1 0 2875 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-978
transform 1 0 2469 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-979
transform 1 0 2944 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-980
transform 1 0 2998 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-981
transform 1 0 3220 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-982
transform 1 0 3208 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-983
transform 1 0 3080 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-984
transform 1 0 2993 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-985
transform 1 0 1912 0 1 901
box 0 0 3 6
use FEEDTHRU  F-986
transform 1 0 3199 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-987
transform 1 0 3247 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-988
transform 1 0 3187 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-989
transform 1 0 3097 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-990
transform 1 0 3202 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-991
transform 1 0 3250 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-992
transform 1 0 3187 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-993
transform 1 0 3101 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-994
transform 1 0 3131 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-995
transform 1 0 3047 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-996
transform 1 0 2927 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-997
transform 1 0 3235 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-998
transform 1 0 2939 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-999
transform 1 0 3067 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1000
transform 1 0 3030 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1001
transform 1 0 3100 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1002
transform 1 0 3190 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1003
transform 1 0 3229 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1004
transform 1 0 3181 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1005
transform 1 0 3104 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1006
transform 1 0 3134 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1007
transform 1 0 3050 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1008
transform 1 0 2942 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1009
transform 1 0 2737 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1010
transform 1 0 2927 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1011
transform 1 0 3070 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1012
transform 1 0 3033 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1013
transform 1 0 3085 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1014
transform 1 0 3175 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1015
transform 1 0 3223 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1016
transform 1 0 3175 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1017
transform 1 0 3089 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1018
transform 1 0 3119 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1019
transform 1 0 3035 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1020
transform 1 0 2665 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1021
transform 1 0 1790 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1022
transform 1 0 3004 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1023
transform 1 0 2922 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1024
transform 1 0 2497 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1025
transform 1 0 2290 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1026
transform 1 0 1924 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1027
transform 1 0 2488 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1028
transform 1 0 2638 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1029
transform 1 0 2060 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1030
transform 1 0 2929 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1031
transform 1 0 2886 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1032
transform 1 0 2995 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1033
transform 1 0 1510 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1034
transform 1 0 1512 0 1 732
box 0 0 3 6
use FEEDTHRU  F-1035
transform 1 0 1525 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1036
transform 1 0 1618 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1037
transform 1 0 1516 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1038
transform 1 0 1531 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1039
transform 1 0 1624 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1040
transform 1 0 1654 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1041
transform 1 0 1682 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1042
transform 1 0 1675 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1043
transform 1 0 1674 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1044
transform 1 0 2338 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1045
transform 1 0 2133 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1046
transform 1 0 2543 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1047
transform 1 0 2646 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1048
transform 1 0 2826 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1049
transform 1 0 2909 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1050
transform 1 0 3017 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1051
transform 1 0 3101 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1052
transform 1 0 3232 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1053
transform 1 0 3157 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1054
transform 1 0 3205 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1055
transform 1 0 3157 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1056
transform 1 0 3061 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1057
transform 1 0 2994 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1058
transform 1 0 3031 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1059
transform 1 0 2885 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1060
transform 1 0 2695 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1061
transform 1 0 2530 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1062
transform 1 0 2360 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1063
transform 1 0 2011 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1064
transform 1 0 2537 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1065
transform 1 0 2640 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1066
transform 1 0 2820 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1067
transform 1 0 2903 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1068
transform 1 0 2423 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1069
transform 1 0 2466 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1070
transform 1 0 1704 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1071
transform 1 0 1697 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1072
transform 1 0 1661 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1073
transform 1 0 2561 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1074
transform 1 0 2465 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1075
transform 1 0 2857 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1076
transform 1 0 3025 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1077
transform 1 0 1777 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1078
transform 1 0 2863 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1079
transform 1 0 1746 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1080
transform 1 0 1735 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1081
transform 1 0 1742 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1082
transform 1 0 1744 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1083
transform 1 0 1714 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1084
transform 1 0 2218 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1085
transform 1 0 2357 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1086
transform 1 0 2430 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1087
transform 1 0 1625 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1088
transform 1 0 3181 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1089
transform 1 0 3133 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1090
transform 1 0 3047 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1091
transform 1 0 3083 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1092
transform 1 0 2999 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1093
transform 1 0 2873 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1094
transform 1 0 3169 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1095
transform 1 0 3121 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1096
transform 1 0 3023 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1097
transform 1 0 3065 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1098
transform 1 0 2981 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1099
transform 1 0 3110 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1100
transform 1 0 3220 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1101
transform 1 0 3262 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1102
transform 1 0 3202 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1103
transform 1 0 3043 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1104
transform 1 0 3141 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1105
transform 1 0 2995 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1106
transform 1 0 3035 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1107
transform 1 0 3140 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1108
transform 1 0 2993 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1109
transform 1 0 2918 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1110
transform 1 0 2817 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1111
transform 1 0 2637 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1112
transform 1 0 2534 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1113
transform 1 0 2335 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1114
transform 1 0 3029 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1115
transform 1 0 3071 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1116
transform 1 0 2987 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1117
transform 1 0 2879 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1118
transform 1 0 2801 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1119
transform 1 0 2784 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1120
transform 1 0 2885 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1121
transform 1 0 2783 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1122
transform 1 0 2742 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1123
transform 1 0 2592 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1124
transform 1 0 2489 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1125
transform 1 0 3047 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1126
transform 1 0 2975 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1127
transform 1 0 3061 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1128
transform 1 0 3109 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1129
transform 1 0 3007 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1130
transform 1 0 2953 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1131
transform 1 0 2832 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1132
transform 1 0 2911 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1133
transform 1 0 1796 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1134
transform 1 0 2632 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1135
transform 1 0 2464 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1136
transform 1 0 2329 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1137
transform 1 0 1936 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1138
transform 1 0 1611 0 1 732
box 0 0 3 6
use FEEDTHRU  F-1139
transform 1 0 2682 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1140
transform 1 0 2613 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1141
transform 1 0 2528 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1142
transform 1 0 2023 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1143
transform 1 0 1923 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1144
transform 1 0 2670 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1145
transform 1 0 2484 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1146
transform 1 0 2369 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1147
transform 1 0 1831 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1148
transform 1 0 1575 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1149
transform 1 0 1762 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1150
transform 1 0 1721 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1151
transform 1 0 2939 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1152
transform 1 0 2897 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1153
transform 1 0 2995 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1154
transform 1 0 3043 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1155
transform 1 0 1801 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1156
transform 1 0 2899 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1157
transform 1 0 1745 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1158
transform 1 0 2915 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1159
transform 1 0 3151 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1160
transform 1 0 3109 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1161
transform 1 0 3007 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1162
transform 1 0 3115 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1163
transform 1 0 3001 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1164
transform 1 0 2946 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1165
transform 1 0 2983 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1166
transform 1 0 2212 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1167
transform 1 0 1684 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1168
transform 1 0 1708 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1169
transform 1 0 1694 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1170
transform 1 0 1711 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1171
transform 1 0 2062 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1172
transform 1 0 1534 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1173
transform 1 0 2110 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1174
transform 1 0 1702 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1175
transform 1 0 1720 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1176
transform 1 0 1700 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1177
transform 1 0 1723 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1178
transform 1 0 2421 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1179
transform 1 0 2611 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1180
transform 1 0 1783 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1181
transform 1 0 3019 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1182
transform 1 0 1540 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1183
transform 1 0 2128 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1184
transform 1 0 1708 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1185
transform 1 0 1738 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1186
transform 1 0 1706 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1187
transform 1 0 1729 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1188
transform 1 0 1740 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1189
transform 1 0 2839 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1190
transform 1 0 1876 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1191
transform 1 0 2091 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1192
transform 1 0 2413 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1193
transform 1 0 2612 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1194
transform 1 0 2704 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1195
transform 1 0 2890 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1196
transform 1 0 2855 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1197
transform 1 0 2975 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1198
transform 1 0 3041 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1199
transform 1 0 3005 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1200
transform 1 0 3103 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1201
transform 1 0 3139 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1202
transform 1 0 3097 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1203
transform 1 0 2977 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1204
transform 1 0 2910 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1205
transform 1 0 2941 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1206
transform 1 0 2810 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1207
transform 1 0 1879 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1208
transform 1 0 2094 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1209
transform 1 0 2296 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1210
transform 1 0 2477 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1211
transform 1 0 2580 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1212
transform 1 0 2772 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1213
transform 1 0 2849 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1214
transform 1 0 2073 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1215
transform 1 0 2272 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1216
transform 1 0 2471 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1217
transform 1 0 2085 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1218
transform 1 0 2242 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1219
transform 1 0 2459 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1220
transform 1 0 2568 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1221
transform 1 0 2748 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1222
transform 1 0 2813 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1223
transform 1 0 2927 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1224
transform 1 0 3017 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1225
transform 1 0 2987 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1226
transform 1 0 3085 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1227
transform 1 0 3127 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1228
transform 1 0 3037 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1229
transform 1 0 2971 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1230
transform 1 0 2892 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1231
transform 1 0 2935 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1232
transform 1 0 2804 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1233
transform 1 0 2260 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1234
transform 1 0 2254 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1235
transform 1 0 2465 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1236
transform 1 0 2574 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1237
transform 1 0 2766 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1238
transform 1 0 2831 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1239
transform 1 0 2969 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1240
transform 1 0 3035 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1241
transform 1 0 2999 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1242
transform 1 0 3097 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1243
transform 1 0 3133 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1244
transform 1 0 3043 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1245
transform 1 0 2417 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1246
transform 1 0 2514 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1247
transform 1 0 2700 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1248
transform 1 0 2771 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1249
transform 1 0 2843 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1250
transform 1 0 2975 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1251
transform 1 0 2921 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1252
transform 1 0 3025 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1253
transform 1 0 3067 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1254
transform 1 0 2420 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1255
transform 1 0 2517 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1256
transform 1 0 2703 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1257
transform 1 0 2774 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1258
transform 1 0 2837 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1259
transform 1 0 2945 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1260
transform 1 0 2915 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1261
transform 1 0 3019 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1262
transform 1 0 3061 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1263
transform 1 0 2399 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1264
transform 1 0 2200 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1265
transform 1 0 1779 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1266
transform 1 0 1672 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1267
transform 1 0 2387 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1268
transform 1 0 2881 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1269
transform 1 0 2909 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1270
transform 1 0 2725 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1271
transform 1 0 2903 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1272
transform 1 0 3019 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1273
transform 1 0 2982 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1274
transform 1 0 3037 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1275
transform 1 0 2557 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1276
transform 1 0 2719 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1277
transform 1 0 2897 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1278
transform 1 0 3013 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1279
transform 1 0 2976 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1280
transform 1 0 3031 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1281
transform 1 0 2560 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1282
transform 1 0 2713 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1283
transform 1 0 2891 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1284
transform 1 0 3007 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1285
transform 1 0 2970 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1286
transform 1 0 3025 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1287
transform 1 0 3133 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1288
transform 1 0 3157 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1289
transform 1 0 2971 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1290
transform 1 0 2916 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1291
transform 1 0 2989 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1292
transform 1 0 3079 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1293
transform 1 0 3121 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1294
transform 1 0 3079 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1295
transform 1 0 2981 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1296
transform 1 0 3011 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1297
transform 1 0 2897 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1298
transform 1 0 2840 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1299
transform 1 0 2846 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1300
transform 1 0 2953 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1301
transform 1 0 2852 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1302
transform 1 0 2947 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1303
transform 1 0 1747 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1304
transform 1 0 1783 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1305
transform 1 0 1716 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1306
transform 1 0 1717 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1307
transform 1 0 1748 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1308
transform 1 0 2221 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1309
transform 1 0 2107 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1310
transform 1 0 2044 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1311
transform 1 0 1723 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1312
transform 1 0 2875 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1313
transform 1 0 1753 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1314
transform 1 0 1709 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1315
transform 1 0 1715 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1316
transform 1 0 1667 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1317
transform 1 0 1661 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1318
transform 1 0 1668 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1319
transform 1 0 1650 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1320
transform 1 0 1577 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1321
transform 1 0 1534 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1322
transform 1 0 1759 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1323
transform 1 0 2593 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1324
transform 1 0 1777 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1325
transform 1 0 1722 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1326
transform 1 0 2930 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1327
transform 1 0 2963 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1328
transform 1 0 2837 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1329
transform 1 0 2945 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1330
transform 1 0 3029 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1331
transform 1 0 2951 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1332
transform 1 0 2957 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1333
transform 1 0 3023 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1334
transform 1 0 2993 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1335
transform 1 0 3091 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1336
transform 1 0 3115 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1337
transform 1 0 3103 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1338
transform 1 0 2983 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1339
transform 1 0 2934 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1340
transform 1 0 2965 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1341
transform 1 0 2867 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1342
transform 1 0 2740 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1343
transform 1 0 2327 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1344
transform 1 0 2448 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1345
transform 1 0 1896 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1346
transform 1 0 2675 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1347
transform 1 0 1769 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1348
transform 1 0 2873 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1349
transform 1 0 2843 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1350
transform 1 0 2442 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1351
transform 1 0 2309 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1352
transform 1 0 2059 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1353
transform 1 0 2933 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1354
transform 1 0 2903 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1355
transform 1 0 3013 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1356
transform 1 0 3037 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1357
transform 1 0 2927 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1358
transform 1 0 2867 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1359
transform 1 0 2753 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1360
transform 1 0 2676 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1361
transform 1 0 2478 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1362
transform 1 0 2363 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1363
transform 1 0 2921 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1364
transform 1 0 2855 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1365
transform 1 0 1594 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1366
transform 1 0 1875 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1367
transform 1 0 2011 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1368
transform 1 0 1868 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1369
transform 1 0 1857 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1370
transform 1 0 1620 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1371
transform 1 0 1613 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1372
transform 1 0 1673 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1373
transform 1 0 1476 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1374
transform 1 0 1521 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1375
transform 1 0 1527 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1376
transform 1 0 1522 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1377
transform 1 0 2035 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1378
transform 1 0 1636 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1379
transform 1 0 1696 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1380
transform 1 0 1718 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1381
transform 1 0 1687 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1382
transform 1 0 1573 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1383
transform 1 0 1672 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1384
transform 1 0 1702 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1385
transform 1 0 1724 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1386
transform 1 0 1693 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1387
transform 1 0 1698 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1388
transform 1 0 1711 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1389
transform 1 0 1741 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1390
transform 1 0 1765 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1391
transform 1 0 1717 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1392
transform 1 0 1697 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1393
transform 1 0 1703 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1394
transform 1 0 1697 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1395
transform 1 0 1637 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1396
transform 1 0 1644 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1397
transform 1 0 1614 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1398
transform 1 0 1579 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1399
transform 1 0 1678 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1400
transform 1 0 2053 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1401
transform 1 0 2167 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1402
transform 1 0 1735 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1403
transform 1 0 1648 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1404
transform 1 0 1672 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1405
transform 1 0 1567 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1406
transform 1 0 1666 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1407
transform 1 0 1678 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1408
transform 1 0 2321 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1409
transform 1 0 2917 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1410
transform 1 0 3013 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1411
transform 1 0 2905 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1412
transform 1 0 2915 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1413
transform 1 0 2963 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1414
transform 1 0 2945 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1415
transform 1 0 3055 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1416
transform 1 0 3079 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1417
transform 1 0 3073 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1418
transform 1 0 2939 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1419
transform 1 0 3043 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1420
transform 1 0 3073 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1421
transform 1 0 3061 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1422
transform 1 0 2935 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1423
transform 1 0 2957 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1424
transform 1 0 2903 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1425
transform 1 0 2789 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1426
transform 1 0 1831 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1427
transform 1 0 2164 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1428
transform 1 0 1720 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1429
transform 1 0 1750 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1430
transform 1 0 1784 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1431
transform 1 0 1753 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1432
transform 1 0 1752 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1433
transform 1 0 2635 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1434
transform 1 0 1813 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1435
transform 1 0 2995 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1436
transform 1 0 1548 0 1 732
box 0 0 3 6
use FEEDTHRU  F-1437
transform 1 0 1567 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1438
transform 1 0 1894 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1439
transform 1 0 2121 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1440
transform 1 0 2290 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1441
transform 1 0 2441 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1442
transform 1 0 2562 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1443
transform 1 0 2760 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1444
transform 1 0 2825 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1445
transform 1 0 2939 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1446
transform 1 0 2987 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1447
transform 1 0 2969 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1448
transform 1 0 3073 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1449
transform 1 0 3091 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1450
transform 1 0 3091 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1451
transform 1 0 2965 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1452
transform 1 0 2124 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1453
transform 1 0 2293 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1454
transform 1 0 2444 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1455
transform 1 0 2565 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1456
transform 1 0 2763 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1457
transform 1 0 2828 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1458
transform 1 0 2942 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1459
transform 1 0 2990 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1460
transform 1 0 2963 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1461
transform 1 0 3067 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1462
transform 1 0 3094 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1463
transform 1 0 3094 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1464
transform 1 0 2968 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1465
transform 1 0 2940 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1466
transform 1 0 2109 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1467
transform 1 0 2278 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1468
transform 1 0 2429 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1469
transform 1 0 2550 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1470
transform 1 0 1512 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-1471
transform 1 0 1549 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1472
transform 1 0 1581 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1473
transform 1 0 1570 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1474
transform 1 0 1506 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-1475
transform 1 0 1519 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1476
transform 1 0 1587 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1477
transform 1 0 1582 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1478
transform 1 0 1727 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1479
transform 1 0 1525 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1480
transform 1 0 1593 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1481
transform 1 0 1588 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1482
transform 1 0 2261 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1483
transform 1 0 2436 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1484
transform 1 0 1734 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1485
transform 1 0 1715 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1486
transform 1 0 1775 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1487
transform 1 0 2783 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1488
transform 1 0 2579 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1489
transform 1 0 2941 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1490
transform 1 0 2971 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1491
transform 1 0 1807 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1492
transform 1 0 1543 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1493
transform 1 0 1623 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1494
transform 1 0 1606 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1495
transform 1 0 2460 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1496
transform 1 0 2351 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1497
transform 1 0 2664 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1498
transform 1 0 2735 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1499
transform 1 0 2849 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1500
transform 1 0 2897 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1501
transform 1 0 2891 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1502
transform 1 0 3001 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1503
transform 1 0 3007 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1504
transform 1 0 2977 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1505
transform 1 0 2887 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1506
transform 1 0 1914 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1507
transform 1 0 2791 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1508
transform 1 0 2018 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1509
transform 1 0 2658 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1510
transform 1 0 2454 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1511
transform 1 0 2345 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1512
transform 1 0 1792 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1513
transform 1 0 1659 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1514
transform 1 0 1567 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1515
transform 1 0 2803 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1516
transform 1 0 2821 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1517
transform 1 0 2767 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1518
transform 1 0 2779 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1519
transform 1 0 2736 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1520
transform 1 0 2807 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1521
transform 1 0 2921 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1522
transform 1 0 2969 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1523
transform 1 0 2951 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1524
transform 1 0 3049 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1525
transform 1 0 3055 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1526
transform 1 0 3067 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1527
transform 1 0 2947 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1528
transform 1 0 2943 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1529
transform 1 0 2959 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1530
transform 1 0 2864 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1531
transform 1 0 2692 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1532
transform 1 0 2536 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1533
transform 1 0 2293 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1534
transform 1 0 2532 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1535
transform 1 0 2411 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1536
transform 1 0 2266 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1537
transform 1 0 2730 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1538
transform 1 0 2526 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1539
transform 1 0 1906 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1540
transform 1 0 1545 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-1541
transform 1 0 1594 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1542
transform 1 0 1605 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1543
transform 1 0 1655 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1544
transform 1 0 1600 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1545
transform 1 0 2412 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1546
transform 1 0 1644 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1547
transform 1 0 1686 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1548
transform 1 0 1685 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1549
transform 1 0 1727 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1550
transform 1 0 1638 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1551
transform 1 0 1692 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1552
transform 1 0 2857 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1553
transform 1 0 2079 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1554
transform 1 0 2878 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1555
transform 1 0 1802 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1556
transform 1 0 2971 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1557
transform 1 0 2965 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1558
transform 1 0 2959 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1559
transform 1 0 2861 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1560
transform 1 0 2845 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1561
transform 1 0 1831 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1562
transform 1 0 2953 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1563
transform 1 0 2947 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1564
transform 1 0 2849 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1565
transform 1 0 2879 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1566
transform 1 0 1878 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1567
transform 1 0 1891 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1568
transform 1 0 1904 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1569
transform 1 0 1984 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1570
transform 1 0 1657 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1571
transform 1 0 1717 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1572
transform 1 0 1693 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1573
transform 1 0 1663 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1574
transform 1 0 1723 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1575
transform 1 0 1699 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1576
transform 1 0 1681 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1577
transform 1 0 1619 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1578
transform 1 0 1637 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1579
transform 1 0 1686 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1580
transform 1 0 1669 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1581
transform 1 0 1729 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1582
transform 1 0 1705 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1583
transform 1 0 1687 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1584
transform 1 0 1625 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1585
transform 1 0 1643 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1586
transform 1 0 1692 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1587
transform 1 0 1687 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1588
transform 1 0 1735 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1589
transform 1 0 1711 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1590
transform 1 0 1693 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1591
transform 1 0 1631 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1592
transform 1 0 1649 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1593
transform 1 0 1685 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1594
transform 1 0 1619 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1595
transform 1 0 2265 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1596
transform 1 0 1797 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1597
transform 1 0 1826 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1598
transform 1 0 1939 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1599
transform 1 0 1851 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1600
transform 1 0 1696 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1601
transform 1 0 1661 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1602
transform 1 0 1723 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1603
transform 1 0 1667 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1604
transform 1 0 1741 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1605
transform 1 0 1747 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1606
transform 1 0 1753 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1607
transform 1 0 1685 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1608
transform 1 0 1685 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1609
transform 1 0 1709 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1610
transform 1 0 1643 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1611
transform 1 0 1656 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1612
transform 1 0 1602 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1613
transform 1 0 2393 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1614
transform 1 0 2496 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1615
transform 1 0 2718 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1616
transform 1 0 2795 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1617
transform 1 0 2909 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1618
transform 1 0 2951 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1619
transform 1 0 2927 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1620
transform 1 0 2499 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1621
transform 1 0 2721 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1622
transform 1 0 2989 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1623
transform 1 0 2885 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1624
transform 1 0 2989 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1625
transform 1 0 2989 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1626
transform 1 0 2983 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1627
transform 1 0 1837 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1628
transform 1 0 1885 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1629
transform 1 0 2833 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1630
transform 1 0 1788 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1631
transform 1 0 1807 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1632
transform 1 0 1820 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1633
transform 1 0 2827 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1634
transform 1 0 1872 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1635
transform 1 0 1879 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1636
transform 1 0 1892 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1637
transform 1 0 1972 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1638
transform 1 0 1792 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1639
transform 1 0 2188 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1640
transform 1 0 1963 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1641
transform 1 0 2941 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1642
transform 1 0 2935 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1643
transform 1 0 2837 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1644
transform 1 0 2867 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1645
transform 1 0 1781 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1646
transform 1 0 1739 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1647
transform 1 0 1800 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1648
transform 1 0 2316 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1649
transform 1 0 2189 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1650
transform 1 0 1663 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1651
transform 1 0 1588 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1652
transform 1 0 1549 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1653
transform 1 0 1969 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1654
transform 1 0 2071 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1655
transform 1 0 2195 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1656
transform 1 0 2230 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1657
transform 1 0 2175 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1658
transform 1 0 1870 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1659
transform 1 0 2044 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1660
transform 1 0 1828 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1661
transform 1 0 1828 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1662
transform 1 0 1850 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1663
transform 1 0 1555 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1664
transform 1 0 1660 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1665
transform 1 0 1690 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1666
transform 1 0 1736 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1667
transform 1 0 1705 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1668
transform 1 0 1710 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1669
transform 1 0 1681 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1670
transform 1 0 1771 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1671
transform 1 0 1723 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1672
transform 1 0 1711 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1673
transform 1 0 1655 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1674
transform 1 0 1904 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1675
transform 1 0 2114 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1676
transform 1 0 2054 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1677
transform 1 0 2013 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1678
transform 1 0 1725 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1679
transform 1 0 1742 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1680
transform 1 0 1793 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1681
transform 1 0 2861 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1682
transform 1 0 2831 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1683
transform 1 0 2929 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1684
transform 1 0 2935 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1685
transform 1 0 1799 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1686
transform 1 0 2855 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1687
transform 1 0 2825 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1688
transform 1 0 2923 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1689
transform 1 0 2929 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1690
transform 1 0 1897 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1691
transform 1 0 2821 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1692
transform 1 0 1794 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1693
transform 1 0 1849 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1694
transform 1 0 1880 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1695
transform 1 0 1834 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1696
transform 1 0 1835 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1697
transform 1 0 1907 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1698
transform 1 0 1830 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1699
transform 1 0 2358 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1700
transform 1 0 2255 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1701
transform 1 0 1648 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1702
transform 1 0 2831 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1703
transform 1 0 1729 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1704
transform 1 0 1741 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1705
transform 1 0 1789 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1706
transform 1 0 1699 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1707
transform 1 0 1728 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1708
transform 1 0 1673 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1709
transform 1 0 1673 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1710
transform 1 0 1733 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1711
transform 1 0 1649 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1712
transform 1 0 1662 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1713
transform 1 0 1608 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1714
transform 1 0 1735 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1715
transform 1 0 1679 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1716
transform 1 0 1679 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1717
transform 1 0 1739 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1718
transform 1 0 1655 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1719
transform 1 0 3049 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1720
transform 1 0 2911 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1721
transform 1 0 3055 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1722
transform 1 0 3013 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1723
transform 1 0 2874 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1724
transform 1 0 2923 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1725
transform 1 0 2917 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1726
transform 1 0 2828 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1727
transform 1 0 2656 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1728
transform 1 0 2506 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1729
transform 1 0 2257 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1730
transform 1 0 1957 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1731
transform 1 0 2868 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1732
transform 1 0 2881 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1733
transform 1 0 3025 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1734
transform 1 0 2983 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1735
transform 1 0 2977 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1736
transform 1 0 2879 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1737
transform 1 0 2909 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1738
transform 1 0 1665 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1739
transform 1 0 1756 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1740
transform 1 0 1768 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1741
transform 1 0 2182 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1742
transform 1 0 1774 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1743
transform 1 0 1816 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1744
transform 1 0 1874 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1745
transform 1 0 1837 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1746
transform 1 0 1806 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1747
transform 1 0 2815 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1748
transform 1 0 2917 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1749
transform 1 0 2923 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1750
transform 1 0 2917 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1751
transform 1 0 2819 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1752
transform 1 0 2849 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1753
transform 1 0 1979 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1754
transform 1 0 1853 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1755
transform 1 0 1824 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1756
transform 1 0 2340 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1757
transform 1 0 2219 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1758
transform 1 0 1678 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1759
transform 1 0 1947 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1760
transform 1 0 1909 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1761
transform 1 0 1608 0 1 732
box 0 0 3 6
use FEEDTHRU  F-1762
transform 1 0 1738 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1763
transform 1 0 2176 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1764
transform 1 0 1762 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1765
transform 1 0 1786 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1766
transform 1 0 1850 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1767
transform 1 0 1831 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1768
transform 1 0 1824 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1769
transform 1 0 2779 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1770
transform 1 0 2749 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1771
transform 1 0 2887 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1772
transform 1 0 2869 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1773
transform 1 0 2717 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1774
transform 1 0 2825 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1775
transform 1 0 1943 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1776
transform 1 0 1829 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1777
transform 1 0 1818 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1778
transform 1 0 2322 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1779
transform 1 0 2207 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1780
transform 1 0 1672 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1781
transform 1 0 1650 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1782
transform 1 0 1888 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1783
transform 1 0 2170 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1784
transform 1 0 1744 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1785
transform 1 0 1780 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1786
transform 1 0 1826 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1787
transform 1 0 1819 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1788
transform 1 0 1860 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1789
transform 1 0 2725 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1790
transform 1 0 2695 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1791
transform 1 0 2881 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1792
transform 1 0 2863 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1793
transform 1 0 2711 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1794
transform 1 0 2789 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1795
transform 1 0 1937 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1796
transform 1 0 1769 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1797
transform 1 0 1741 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1798
transform 1 0 1770 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1799
transform 1 0 1735 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1800
transform 1 0 1825 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1801
transform 1 0 1795 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1802
transform 1 0 1765 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1803
transform 1 0 1772 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1804
transform 1 0 1726 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1805
transform 1 0 1696 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1806
transform 1 0 1778 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1807
transform 1 0 1747 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1808
transform 1 0 1776 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1809
transform 1 0 1741 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1810
transform 1 0 1732 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1811
transform 1 0 2158 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1812
transform 1 0 1732 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1813
transform 1 0 1768 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1814
transform 1 0 1814 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1815
transform 1 0 1801 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1816
transform 1 0 1842 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1817
transform 1 0 1828 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1818
transform 1 0 2152 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1819
transform 1 0 1726 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1820
transform 1 0 1762 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1821
transform 1 0 1808 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1822
transform 1 0 1789 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1823
transform 1 0 1848 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1824
transform 1 0 2617 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1825
transform 1 0 1915 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1826
transform 1 0 2839 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1827
transform 1 0 2821 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1828
transform 1 0 2543 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1829
transform 1 0 2717 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1830
transform 1 0 1805 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1831
transform 1 0 1721 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1832
transform 1 0 1746 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1833
transform 1 0 2256 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1834
transform 1 0 1840 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1835
transform 1 0 1886 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1836
transform 1 0 2572 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1837
transform 1 0 1990 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1838
transform 1 0 2290 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1839
transform 1 0 1930 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1840
transform 1 0 2485 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1841
transform 1 0 2629 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1842
transform 1 0 2795 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1843
transform 1 0 2887 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1844
transform 1 0 2482 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1845
transform 1 0 2626 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1846
transform 1 0 2792 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1847
transform 1 0 2230 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1848
transform 1 0 2476 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1849
transform 1 0 2620 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1850
transform 1 0 2714 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1851
transform 1 0 2890 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1852
transform 1 0 2880 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1853
transform 1 0 2851 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1854
transform 1 0 3001 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1855
transform 1 0 2959 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1856
transform 1 0 2953 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1857
transform 1 0 2855 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1858
transform 1 0 2885 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1859
transform 1 0 2861 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1860
transform 1 0 2747 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1861
transform 1 0 2825 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1862
transform 1 0 2905 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1863
transform 1 0 2904 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1864
transform 1 0 2875 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1865
transform 1 0 2653 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1866
transform 1 0 2500 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1867
transform 1 0 2248 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1868
transform 1 0 1985 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1869
transform 1 0 2650 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1870
transform 1 0 2822 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1871
transform 1 0 2908 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1872
transform 1 0 2907 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1873
transform 1 0 2878 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1874
transform 1 0 3019 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1875
transform 1 0 2977 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1876
transform 1 0 2971 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1877
transform 1 0 2873 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1878
transform 1 0 2903 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1879
transform 1 0 2879 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1880
transform 1 0 2765 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1881
transform 1 0 2694 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1882
transform 1 0 2472 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1883
transform 1 0 2381 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1884
transform 1 0 2248 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1885
transform 1 0 1787 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1886
transform 1 0 1703 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1887
transform 1 0 1710 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1888
transform 1 0 1692 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1889
transform 1 0 1751 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1890
transform 1 0 1793 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1891
transform 1 0 2587 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1892
transform 1 0 2731 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1893
transform 1 0 1849 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1894
transform 1 0 2923 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1895
transform 1 0 2785 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1896
transform 1 0 1920 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1897
transform 1 0 1843 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1898
transform 1 0 1970 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1899
transform 1 0 2116 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1900
transform 1 0 2392 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1901
transform 1 0 2917 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1902
transform 1 0 2911 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1903
transform 1 0 2789 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1904
transform 1 0 2965 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1905
transform 1 0 2911 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1906
transform 1 0 2899 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1907
transform 1 0 2777 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1908
transform 1 0 2831 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1909
transform 1 0 1973 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1910
transform 1 0 1847 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1911
transform 1 0 1691 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1912
transform 1 0 1751 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1913
transform 1 0 1667 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1914
transform 1 0 1674 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1915
transform 1 0 1620 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1916
transform 1 0 1559 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1917
transform 1 0 1691 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1918
transform 1 0 1697 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1919
transform 1 0 1757 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1920
transform 1 0 1673 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1921
transform 1 0 1680 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1922
transform 1 0 1626 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1923
transform 1 0 1565 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1924
transform 1 0 1576 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1925
transform 1 0 1776 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1926
transform 1 0 2285 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1927
transform 1 0 2394 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1928
transform 1 0 1842 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1929
transform 1 0 1859 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1930
transform 1 0 2009 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1931
transform 1 0 2837 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1932
transform 1 0 2273 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1933
transform 1 0 1786 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-1934
transform 1 0 1737 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-1935
transform 1 0 1660 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-1936
transform 1 0 2388 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1937
transform 1 0 1848 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1938
transform 1 0 1865 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1939
transform 1 0 2783 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1940
transform 1 0 2843 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1941
transform 1 0 2783 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1942
transform 1 0 2905 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1943
transform 1 0 1752 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1944
transform 1 0 2220 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1945
transform 1 0 1745 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1946
transform 1 0 1871 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1947
transform 1 0 2765 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1948
transform 1 0 1859 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1949
transform 1 0 2797 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1950
transform 1 0 2815 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1951
transform 1 0 1945 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1952
transform 1 0 1913 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1953
transform 1 0 2741 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1954
transform 1 0 1763 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1955
transform 1 0 1770 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1956
transform 1 0 2250 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1957
transform 1 0 2129 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-1958
transform 1 0 1811 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1959
transform 1 0 1877 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1960
transform 1 0 1727 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1961
transform 1 0 2563 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1962
transform 1 0 2569 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1963
transform 1 0 1879 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1964
transform 1 0 1771 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1965
transform 1 0 1829 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1966
transform 1 0 1871 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1967
transform 1 0 1739 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1968
transform 1 0 2473 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1969
transform 1 0 2491 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1970
transform 1 0 1867 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1971
transform 1 0 1753 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1972
transform 1 0 1805 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1973
transform 1 0 1787 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-1974
transform 1 0 2461 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1975
transform 1 0 2479 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-1976
transform 1 0 1855 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1977
transform 1 0 1903 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-1978
transform 1 0 1807 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-1979
transform 1 0 1866 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1980
transform 1 0 1813 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1981
transform 1 0 2555 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1982
transform 1 0 1925 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1983
transform 1 0 2501 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-1984
transform 1 0 1919 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-1985
transform 1 0 1823 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-1986
transform 1 0 1806 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-1987
transform 1 0 2274 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-1988
transform 1 0 2725 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-1989
transform 1 0 2206 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1990
transform 1 0 2446 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1991
transform 1 0 2554 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1992
transform 1 0 2200 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-1993
transform 1 0 2440 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-1994
transform 1 0 1942 0 1 901
box 0 0 3 6
use FEEDTHRU  F-1995
transform 1 0 2590 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1996
transform 1 0 2768 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-1997
transform 1 0 2851 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-1998
transform 1 0 2862 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-1999
transform 1 0 2809 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2000
transform 1 0 2953 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2001
transform 1 0 2899 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2002
transform 1 0 2881 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2003
transform 1 0 2801 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2004
transform 1 0 2819 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2005
transform 1 0 2813 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2006
transform 1 0 2711 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2007
transform 1 0 2458 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2008
transform 1 0 2614 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2009
transform 1 0 2786 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2010
transform 1 0 2032 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2011
transform 1 0 1750 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2012
transform 1 0 1798 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2013
transform 1 0 1838 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2014
transform 1 0 1900 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2015
transform 1 0 1705 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2016
transform 1 0 2020 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2017
transform 1 0 1756 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2018
transform 1 0 1810 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2019
transform 1 0 1844 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2020
transform 1 0 1783 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2021
transform 1 0 1812 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2022
transform 1 0 1596 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-2023
transform 1 0 1891 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2024
transform 1 0 2130 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2025
transform 1 0 1894 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2026
transform 1 0 2315 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2027
transform 1 0 2424 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2028
transform 1 0 2640 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2029
transform 1 0 2705 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2030
transform 1 0 2807 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2031
transform 1 0 2801 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2032
transform 1 0 2795 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2033
transform 1 0 2875 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2034
transform 1 0 2893 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2035
transform 1 0 2947 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2036
transform 1 0 2803 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2037
transform 1 0 2856 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2038
transform 1 0 2839 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2039
transform 1 0 2774 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2040
transform 1 0 2602 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2041
transform 1 0 2452 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2042
transform 1 0 2194 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2043
transform 1 0 1960 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2044
transform 1 0 1599 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-2045
transform 1 0 1675 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2046
transform 1 0 1681 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2047
transform 1 0 1687 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2048
transform 1 0 1830 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2049
transform 1 0 2167 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2050
transform 1 0 2321 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2051
transform 1 0 2418 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2052
transform 1 0 2622 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2053
transform 1 0 2687 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2054
transform 1 0 2789 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2055
transform 1 0 2795 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2056
transform 1 0 2652 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2057
transform 1 0 2750 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2058
transform 1 0 2864 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2059
transform 1 0 2888 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2060
transform 1 0 2858 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2061
transform 1 0 2956 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2062
transform 1 0 2655 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2063
transform 1 0 2723 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2064
transform 1 0 2825 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2065
transform 1 0 2807 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2066
transform 1 0 2807 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2067
transform 1 0 2887 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2068
transform 1 0 2962 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2069
transform 1 0 3004 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2070
transform 1 0 1589 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2071
transform 1 0 1656 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2072
transform 1 0 1716 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2073
transform 1 0 1727 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2074
transform 1 0 1817 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2075
transform 1 0 1595 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2076
transform 1 0 1680 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2077
transform 1 0 1722 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2078
transform 1 0 1733 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2079
transform 1 0 1823 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2080
transform 1 0 1721 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2081
transform 1 0 1721 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2082
transform 1 0 1789 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2083
transform 1 0 1789 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2084
transform 1 0 1843 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2085
transform 1 0 1723 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2086
transform 1 0 1800 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2087
transform 1 0 1771 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2088
transform 1 0 1832 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2089
transform 1 0 1792 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2090
transform 1 0 1601 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2091
transform 1 0 1662 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2092
transform 1 0 1822 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2093
transform 1 0 1856 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2094
transform 1 0 1795 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2095
transform 1 0 1830 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2096
transform 1 0 1759 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2097
transform 1 0 1873 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2098
transform 1 0 2473 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2099
transform 1 0 2455 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2100
transform 1 0 1751 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2101
transform 1 0 1781 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2102
transform 1 0 1847 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2103
transform 1 0 1757 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2104
transform 1 0 1768 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2105
transform 1 0 1828 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2106
transform 1 0 1862 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2107
transform 1 0 1939 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2108
transform 1 0 2826 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2109
transform 1 0 2773 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2110
transform 1 0 2911 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2111
transform 1 0 2869 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2112
transform 1 0 2851 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2113
transform 1 0 3116 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2114
transform 1 0 2759 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2115
transform 1 0 1963 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2116
transform 1 0 2814 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2117
transform 1 0 2761 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2118
transform 1 0 2893 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2119
transform 1 0 2851 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2120
transform 1 0 2833 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2121
transform 1 0 2753 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2122
transform 1 0 2753 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2123
transform 1 0 3014 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2124
transform 1 0 2900 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2125
transform 1 0 2535 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2126
transform 1 0 2382 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2127
transform 1 0 2297 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2128
transform 1 0 2726 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2129
transform 1 0 2779 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2130
transform 1 0 2808 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2131
transform 1 0 2755 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2132
transform 1 0 2887 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2133
transform 1 0 2845 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2134
transform 1 0 2827 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2135
transform 1 0 2747 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2136
transform 1 0 2747 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2137
transform 1 0 2771 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2138
transform 1 0 1913 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2139
transform 1 0 1893 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2140
transform 1 0 2385 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2141
transform 1 0 1976 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2142
transform 1 0 1861 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2143
transform 1 0 2012 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2144
transform 1 0 1867 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2145
transform 1 0 1890 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2146
transform 1 0 1897 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2147
transform 1 0 1921 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2148
transform 1 0 2719 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2149
transform 1 0 2707 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2150
transform 1 0 2459 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2151
transform 1 0 2399 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2152
transform 1 0 1931 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2153
transform 1 0 1835 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2154
transform 1 0 2368 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2155
transform 1 0 2140 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2156
transform 1 0 1834 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2157
transform 1 0 1566 0 1 732
box 0 0 3 6
use FEEDTHRU  F-2158
transform 1 0 1612 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2159
transform 1 0 1631 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2160
transform 1 0 1618 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2161
transform 1 0 1637 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2162
transform 1 0 1686 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2163
transform 1 0 1740 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2164
transform 1 0 1751 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2165
transform 1 0 1841 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2166
transform 1 0 1757 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2167
transform 1 0 1745 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2168
transform 1 0 1624 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2169
transform 1 0 1599 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2170
transform 1 0 2941 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2171
transform 1 0 2883 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2172
transform 1 0 2869 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2173
transform 1 0 2838 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2174
transform 1 0 2857 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2175
transform 1 0 2671 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2176
transform 1 0 1939 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2177
transform 1 0 2659 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2178
transform 1 0 2357 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2179
transform 1 0 2665 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2180
transform 1 0 2647 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2181
transform 1 0 2079 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2182
transform 1 0 2396 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2183
transform 1 0 2406 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2184
transform 1 0 2634 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2185
transform 1 0 2699 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2186
transform 1 0 2801 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2187
transform 1 0 2777 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2188
transform 1 0 2771 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2189
transform 1 0 2845 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2190
transform 1 0 2863 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2191
transform 1 0 2935 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2192
transform 1 0 2797 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2193
transform 1 0 2333 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2194
transform 1 0 2400 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2195
transform 1 0 2628 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2196
transform 1 0 2693 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2197
transform 1 0 2795 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2198
transform 1 0 2771 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2199
transform 1 0 2765 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2200
transform 1 0 2839 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2201
transform 1 0 2857 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2202
transform 1 0 2929 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2203
transform 1 0 2791 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2204
transform 1 0 2844 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2205
transform 1 0 2863 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2206
transform 1 0 2798 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2207
transform 1 0 2773 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2208
transform 1 0 2705 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2209
transform 1 0 2723 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2210
transform 1 0 2003 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2211
transform 1 0 1901 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2212
transform 1 0 1878 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2213
transform 1 0 2352 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2214
transform 1 0 2300 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2215
transform 1 0 2809 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2216
transform 1 0 2809 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2217
transform 1 0 2731 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2218
transform 1 0 2802 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2219
transform 1 0 2857 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2220
transform 1 0 1829 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2221
transform 1 0 1901 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2222
transform 1 0 1793 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2223
transform 1 0 1776 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2224
transform 1 0 2208 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2225
transform 1 0 2072 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2226
transform 1 0 2053 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2227
transform 1 0 1929 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2228
transform 1 0 1777 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2229
transform 1 0 1494 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-2230
transform 1 0 1817 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2231
transform 1 0 1877 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2232
transform 1 0 1817 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2233
transform 1 0 1794 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2234
transform 1 0 2027 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2235
transform 1 0 2735 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2236
transform 1 0 2741 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2237
transform 1 0 2815 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2238
transform 1 0 2833 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2239
transform 1 0 2905 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2240
transform 1 0 2729 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2241
transform 1 0 2735 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2242
transform 1 0 2809 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2243
transform 1 0 2827 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2244
transform 1 0 2899 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2245
transform 1 0 2767 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2246
transform 1 0 2820 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2247
transform 1 0 2845 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2248
transform 1 0 2780 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2249
transform 1 0 2608 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2250
transform 1 0 2033 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2251
transform 1 0 1925 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2252
transform 1 0 1902 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2253
transform 1 0 1744 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2254
transform 1 0 2092 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2255
transform 1 0 1864 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2256
transform 1 0 1816 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2257
transform 1 0 2086 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2258
transform 1 0 1828 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2259
transform 1 0 1912 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2260
transform 1 0 1922 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2261
transform 1 0 1518 0 1 732
box 0 0 3 6
use FEEDTHRU  F-2262
transform 1 0 1792 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2263
transform 1 0 2068 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2264
transform 1 0 1804 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2265
transform 1 0 1882 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2266
transform 1 0 1910 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2267
transform 1 0 1915 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2268
transform 1 0 2104 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2269
transform 1 0 1930 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2270
transform 1 0 1551 0 1 732
box 0 0 3 6
use FEEDTHRU  F-2271
transform 1 0 1876 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2272
transform 1 0 2098 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2273
transform 1 0 1888 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2274
transform 1 0 1969 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2275
transform 1 0 2736 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2276
transform 1 0 2011 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2277
transform 1 0 2494 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2278
transform 1 0 2350 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2279
transform 1 0 2122 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2280
transform 1 0 1939 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2281
transform 1 0 2132 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2282
transform 1 0 2731 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2283
transform 1 0 2730 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2284
transform 1 0 2671 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2285
transform 1 0 2803 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2286
transform 1 0 2773 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2287
transform 1 0 2761 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2288
transform 1 0 2549 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2289
transform 1 0 2507 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2290
transform 1 0 2665 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2291
transform 1 0 2755 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2292
transform 1 0 2767 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2293
transform 1 0 2694 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2294
transform 1 0 2125 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2295
transform 1 0 2664 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2296
transform 1 0 2683 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2297
transform 1 0 2210 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2298
transform 1 0 1799 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2299
transform 1 0 1883 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2300
transform 1 0 1799 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2301
transform 1 0 1788 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2302
transform 1 0 2196 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2303
transform 1 0 1649 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2304
transform 1 0 1654 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2305
transform 1 0 1811 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2306
transform 1 0 1895 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2307
transform 1 0 1787 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2308
transform 1 0 1775 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2309
transform 1 0 2359 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2310
transform 1 0 2383 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2311
transform 1 0 1889 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2312
transform 1 0 1763 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2313
transform 1 0 1769 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2314
transform 1 0 1805 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2315
transform 1 0 1782 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2316
transform 1 0 1780 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2317
transform 1 0 1846 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2318
transform 1 0 2055 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2319
transform 1 0 1852 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2320
transform 1 0 2061 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2321
transform 1 0 2206 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2322
transform 1 0 2303 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2323
transform 1 0 2376 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2324
transform 1 0 1908 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2325
transform 1 0 1931 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2326
transform 1 0 2183 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2327
transform 1 0 1696 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2328
transform 1 0 1725 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2329
transform 1 0 2165 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2330
transform 1 0 1732 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2331
transform 1 0 2238 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2332
transform 1 0 2147 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2333
transform 1 0 1702 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2334
transform 1 0 1683 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2335
transform 1 0 1780 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2336
transform 1 0 2014 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2337
transform 1 0 1786 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2338
transform 1 0 1906 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2339
transform 1 0 1570 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2340
transform 1 0 1853 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2341
transform 1 0 1775 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2342
transform 1 0 1727 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2343
transform 1 0 1733 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2344
transform 1 0 1759 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2345
transform 1 0 1759 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2346
transform 1 0 1861 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2347
transform 1 0 1729 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2348
transform 1 0 1818 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2349
transform 1 0 1825 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2350
transform 1 0 1868 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2351
transform 1 0 1804 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2352
transform 1 0 1733 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2353
transform 1 0 1859 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2354
transform 1 0 1781 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2355
transform 1 0 1758 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2356
transform 1 0 1668 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2357
transform 1 0 1613 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2358
transform 1 0 1636 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2359
transform 1 0 1611 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2360
transform 1 0 1531 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2361
transform 1 0 1739 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2362
transform 1 0 1865 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2363
transform 1 0 1787 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2364
transform 1 0 1764 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2365
transform 1 0 1674 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2366
transform 1 0 1619 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2367
transform 1 0 1642 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2368
transform 1 0 1617 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2369
transform 1 0 1537 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2370
transform 1 0 1926 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2371
transform 1 0 1955 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2372
transform 1 0 2717 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2373
transform 1 0 2699 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2374
transform 1 0 2729 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2375
transform 1 0 2791 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2376
transform 1 0 2803 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2377
transform 1 0 2881 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2378
transform 1 0 2749 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2379
transform 1 0 2796 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2380
transform 1 0 2833 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2381
transform 1 0 2756 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2382
transform 1 0 1932 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2383
transform 1 0 1973 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2384
transform 1 0 2759 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2385
transform 1 0 2705 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2386
transform 1 0 2586 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2387
transform 1 0 2370 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2388
transform 1 0 2279 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2389
transform 1 0 1985 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2390
transform 1 0 2765 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2391
transform 1 0 2711 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2392
transform 1 0 2723 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2393
transform 1 0 2785 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2394
transform 1 0 2797 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2395
transform 1 0 2875 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2396
transform 1 0 2743 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2397
transform 1 0 2790 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2398
transform 1 0 2821 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2399
transform 1 0 2750 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2400
transform 1 0 2584 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2401
transform 1 0 2404 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2402
transform 1 0 1872 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2403
transform 1 0 1871 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2404
transform 1 0 1955 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2405
transform 1 0 1919 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2406
transform 1 0 2441 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2407
transform 1 0 2479 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2408
transform 1 0 2497 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2409
transform 1 0 1927 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2410
transform 1 0 1813 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2411
transform 1 0 1883 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2412
transform 1 0 1967 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2413
transform 1 0 2779 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2414
transform 1 0 2791 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2415
transform 1 0 2863 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2416
transform 1 0 2785 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2417
transform 1 0 2869 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2418
transform 1 0 2854 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2419
transform 1 0 1770 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2420
transform 1 0 1643 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2421
transform 1 0 2477 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2422
transform 1 0 2623 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2423
transform 1 0 2659 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2424
transform 1 0 2185 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2425
transform 1 0 2557 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2426
transform 1 0 1992 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2427
transform 1 0 2005 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2428
transform 1 0 2036 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2429
transform 1 0 2092 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2430
transform 1 0 2593 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2431
transform 1 0 2617 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2432
transform 1 0 2029 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2433
transform 1 0 2455 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2434
transform 1 0 2657 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2435
transform 1 0 2657 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2436
transform 1 0 2711 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2437
transform 1 0 2651 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2438
transform 1 0 2639 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2439
transform 1 0 2063 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2440
transform 1 0 2665 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2441
transform 1 0 2603 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2442
transform 1 0 2633 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2443
transform 1 0 2695 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2444
transform 1 0 2693 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2445
transform 1 0 2699 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2446
transform 1 0 2669 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2447
transform 1 0 2741 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2448
transform 1 0 2663 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2449
transform 1 0 2592 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2450
transform 1 0 2755 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2451
transform 1 0 2761 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2452
transform 1 0 2851 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2453
transform 1 0 2719 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2454
transform 1 0 2784 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2455
transform 1 0 2815 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2456
transform 1 0 2744 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2457
transform 1 0 2578 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2458
transform 1 0 2422 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2459
transform 1 0 2233 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2460
transform 1 0 2004 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2461
transform 1 0 1834 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2462
transform 1 0 1906 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2463
transform 1 0 2237 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2464
transform 1 0 1719 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2465
transform 1 0 1720 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2466
transform 1 0 2123 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2467
transform 1 0 2214 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2468
transform 1 0 1854 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2469
transform 1 0 1877 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2470
transform 1 0 1961 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2471
transform 1 0 2778 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2472
transform 1 0 2809 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2473
transform 1 0 2713 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2474
transform 1 0 2760 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2475
transform 1 0 2695 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2476
transform 1 0 2833 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2477
transform 1 0 2743 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2478
transform 1 0 2737 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2479
transform 1 0 2681 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2480
transform 1 0 2663 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2481
transform 1 0 2735 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2482
transform 1 0 2657 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2483
transform 1 0 2754 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2484
transform 1 0 2689 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2485
transform 1 0 2827 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2486
transform 1 0 2737 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2487
transform 1 0 2731 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2488
transform 1 0 2675 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2489
transform 1 0 2687 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2490
transform 1 0 2687 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2491
transform 1 0 2743 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2492
transform 1 0 2749 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2493
transform 1 0 2839 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2494
transform 1 0 2701 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2495
transform 1 0 2766 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2496
transform 1 0 2675 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2497
transform 1 0 2747 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2498
transform 1 0 2681 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2499
transform 1 0 1936 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2500
transform 1 0 1994 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2501
transform 1 0 1945 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2502
transform 1 0 1882 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2503
transform 1 0 2056 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2504
transform 1 0 1690 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2505
transform 1 0 1709 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2506
transform 1 0 2172 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2507
transform 1 0 1836 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2508
transform 1 0 1673 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2509
transform 1 0 2876 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2510
transform 1 0 2906 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2511
transform 1 0 2882 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2512
transform 1 0 2974 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2513
transform 1 0 2980 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2514
transform 1 0 3022 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2515
transform 1 0 2707 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2516
transform 1 0 2772 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2517
transform 1 0 2827 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2518
transform 1 0 2762 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2519
transform 1 0 2596 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2520
transform 1 0 1775 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2521
transform 1 0 1757 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2522
transform 1 0 1771 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2523
transform 1 0 1771 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2524
transform 1 0 1769 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2525
transform 1 0 1907 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2526
transform 1 0 1841 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2527
transform 1 0 1812 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2528
transform 1 0 1763 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2529
transform 1 0 1777 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2530
transform 1 0 1777 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2531
transform 1 0 2328 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2532
transform 1 0 1950 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2533
transform 1 0 2009 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2534
transform 1 0 2081 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2535
transform 1 0 2597 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2536
transform 1 0 2609 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2537
transform 1 0 2701 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2538
transform 1 0 2713 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2539
transform 1 0 2791 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2540
transform 1 0 2653 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2541
transform 1 0 2718 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2542
transform 1 0 2749 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2543
transform 1 0 2678 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2544
transform 1 0 2524 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2545
transform 1 0 2380 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2546
transform 1 0 2116 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2547
transform 1 0 1986 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2548
transform 1 0 2639 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2549
transform 1 0 2693 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2550
transform 1 0 2603 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2551
transform 1 0 2633 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2552
transform 1 0 2689 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2553
transform 1 0 2701 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2554
transform 1 0 2773 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2555
transform 1 0 2082 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2556
transform 1 0 2645 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2557
transform 1 0 2699 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2558
transform 1 0 2621 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2559
transform 1 0 2639 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2560
transform 1 0 2821 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2561
transform 1 0 2725 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2562
transform 1 0 2719 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2563
transform 1 0 2669 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2564
transform 1 0 2651 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2565
transform 1 0 2729 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2566
transform 1 0 2683 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2567
transform 1 0 2748 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2568
transform 1 0 2803 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2569
transform 1 0 2738 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2570
transform 1 0 2572 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2571
transform 1 0 2416 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2572
transform 1 0 2742 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2573
transform 1 0 2797 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2574
transform 1 0 2732 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2575
transform 1 0 2677 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2576
transform 1 0 2815 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2577
transform 1 0 2724 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2578
transform 1 0 2767 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2579
transform 1 0 2702 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2580
transform 1 0 2542 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2581
transform 1 0 2659 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2582
transform 1 0 2797 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2583
transform 1 0 2707 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2584
transform 1 0 2695 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2585
transform 1 0 2645 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2586
transform 1 0 2627 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2587
transform 1 0 2705 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2588
transform 1 0 2651 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2589
transform 1 0 2580 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2590
transform 1 0 2334 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2591
transform 1 0 2249 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2592
transform 1 0 2191 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2593
transform 1 0 2040 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2594
transform 1 0 2773 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2595
transform 1 0 2708 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2596
transform 1 0 2548 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2597
transform 1 0 2398 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2598
transform 1 0 1962 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2599
transform 1 0 2027 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2600
transform 1 0 2681 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2601
transform 1 0 2310 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2602
transform 1 0 2224 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2603
transform 1 0 2267 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2604
transform 1 0 2346 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2605
transform 1 0 2610 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2606
transform 1 0 2669 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2607
transform 1 0 2723 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2608
transform 1 0 2645 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2609
transform 1 0 2663 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2610
transform 1 0 2713 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2611
transform 1 0 2567 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2612
transform 1 0 2605 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2613
transform 1 0 2647 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2614
transform 1 0 2437 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2615
transform 1 0 2545 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2616
transform 1 0 2028 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2617
transform 1 0 2561 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2618
transform 1 0 2525 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2619
transform 1 0 2039 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2620
transform 1 0 1979 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2621
transform 1 0 1930 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2622
transform 1 0 2134 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2623
transform 1 0 2419 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2624
transform 1 0 2560 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2625
transform 1 0 2720 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2626
transform 1 0 2785 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2627
transform 1 0 1563 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-2628
transform 1 0 1789 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2629
transform 1 0 2001 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2630
transform 1 0 2161 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2631
transform 1 0 1735 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2632
transform 1 0 1896 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2633
transform 1 0 2158 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2634
transform 1 0 2213 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2635
transform 1 0 2280 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2636
transform 1 0 1980 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2637
transform 1 0 2332 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2638
transform 1 0 2074 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2639
transform 1 0 1954 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2640
transform 1 0 1560 0 1 732
box 0 0 3 6
use FEEDTHRU  F-2641
transform 1 0 2344 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2642
transform 1 0 2476 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2643
transform 1 0 2084 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2644
transform 1 0 2029 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2645
transform 1 0 1998 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2646
transform 1 0 2473 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2647
transform 1 0 2215 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2648
transform 1 0 2599 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2649
transform 1 0 2008 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2650
transform 1 0 1858 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2651
transform 1 0 1906 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2652
transform 1 0 1946 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2653
transform 1 0 1603 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2654
transform 1 0 1972 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2655
transform 1 0 1609 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2656
transform 1 0 1954 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2657
transform 1 0 1840 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2658
transform 1 0 1888 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2659
transform 1 0 1928 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2660
transform 1 0 1885 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2661
transform 1 0 1846 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2662
transform 1 0 1630 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2663
transform 1 0 1494 0 1 732
box 0 0 3 6
use FEEDTHRU  F-2664
transform 1 0 1636 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2665
transform 1 0 1689 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2666
transform 1 0 1750 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2667
transform 1 0 1642 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2668
transform 1 0 1701 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2669
transform 1 0 2483 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2670
transform 1 0 2581 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2671
transform 1 0 2581 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2672
transform 1 0 2047 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2673
transform 1 0 2305 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2674
transform 1 0 1962 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2675
transform 1 0 1987 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2676
transform 1 0 2465 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2677
transform 1 0 2015 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2678
transform 1 0 1961 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2679
transform 1 0 1473 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-2680
transform 1 0 1585 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2681
transform 1 0 1671 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2682
transform 1 0 1708 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2683
transform 1 0 1661 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2684
transform 1 0 1728 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2685
transform 1 0 1860 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2686
transform 1 0 1889 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2687
transform 1 0 1949 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2688
transform 1 0 1811 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2689
transform 1 0 1799 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2690
transform 1 0 1867 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2691
transform 1 0 2068 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2692
transform 1 0 2272 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2693
transform 1 0 2050 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2694
transform 1 0 2283 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2695
transform 1 0 2332 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2696
transform 1 0 2309 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2697
transform 1 0 1591 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2698
transform 1 0 1677 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2699
transform 1 0 1714 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2700
transform 1 0 1667 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2701
transform 1 0 1704 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2702
transform 1 0 1866 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2703
transform 1 0 1895 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2704
transform 1 0 1898 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2705
transform 1 0 1855 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2706
transform 1 0 1836 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2707
transform 1 0 1747 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2708
transform 1 0 1891 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2709
transform 1 0 1783 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2710
transform 1 0 1783 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2711
transform 1 0 1781 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2712
transform 1 0 1793 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2713
transform 1 0 2615 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2714
transform 1 0 2627 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2715
transform 1 0 2683 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2716
transform 1 0 2689 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2717
transform 1 0 2785 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2718
transform 1 0 2647 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2719
transform 1 0 2609 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2720
transform 1 0 2621 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2721
transform 1 0 2677 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2722
transform 1 0 2683 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2723
transform 1 0 2615 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2724
transform 1 0 2671 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2725
transform 1 0 2677 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2726
transform 1 0 2779 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2727
transform 1 0 2641 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2728
transform 1 0 2712 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2729
transform 1 0 2755 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2730
transform 1 0 2696 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2731
transform 1 0 2536 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2732
transform 1 0 2537 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2733
transform 1 0 2495 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2734
transform 1 0 2021 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2735
transform 1 0 1967 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2736
transform 1 0 1944 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2737
transform 1 0 2226 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2738
transform 1 0 2177 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2739
transform 1 0 1852 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2740
transform 1 0 1800 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2741
transform 1 0 2587 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2742
transform 1 0 2053 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2743
transform 1 0 2329 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2744
transform 1 0 1986 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2745
transform 1 0 1993 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2746
transform 1 0 2030 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2747
transform 1 0 2008 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2748
transform 1 0 2128 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2749
transform 1 0 2050 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2750
transform 1 0 1858 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2751
transform 1 0 2148 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2752
transform 1 0 2615 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2753
transform 1 0 2657 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2754
transform 1 0 2591 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2755
transform 1 0 2597 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2756
transform 1 0 2653 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2757
transform 1 0 2653 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2758
transform 1 0 2731 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2759
transform 1 0 2605 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2760
transform 1 0 2322 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2761
transform 1 0 2191 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2762
transform 1 0 2100 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2763
transform 1 0 2069 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2764
transform 1 0 2141 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2765
transform 1 0 2130 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2766
transform 1 0 2123 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2767
transform 1 0 2195 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2768
transform 1 0 2579 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2769
transform 1 0 2591 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2770
transform 1 0 2641 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2771
transform 1 0 2641 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2772
transform 1 0 2677 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2773
transform 1 0 2551 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2774
transform 1 0 2064 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2775
transform 1 0 2053 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2776
transform 1 0 2153 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2777
transform 1 0 2651 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2778
transform 1 0 1849 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2779
transform 1 0 1993 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2780
transform 1 0 2527 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2781
transform 1 0 2515 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2782
transform 1 0 2519 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2783
transform 1 0 2477 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2784
transform 1 0 1938 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2785
transform 1 0 1855 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2786
transform 1 0 1999 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2787
transform 1 0 2515 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2788
transform 1 0 2503 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2789
transform 1 0 2489 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2790
transform 1 0 1950 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2791
transform 1 0 1885 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2792
transform 1 0 2005 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2793
transform 1 0 2706 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2794
transform 1 0 2629 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2795
transform 1 0 2767 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2796
transform 1 0 2761 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2797
transform 1 0 2700 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2798
transform 1 0 2623 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2799
transform 1 0 2761 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2800
transform 1 0 2630 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2801
transform 1 0 2689 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2802
transform 1 0 2382 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2803
transform 1 0 2563 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2804
transform 1 0 2701 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2805
transform 1 0 2635 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2806
transform 1 0 2635 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2807
transform 1 0 2666 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2808
transform 1 0 2719 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2809
transform 1 0 2646 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2810
transform 1 0 2575 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2811
transform 1 0 2713 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2812
transform 1 0 2629 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2813
transform 1 0 2629 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2814
transform 1 0 2585 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2815
transform 1 0 2585 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2816
transform 1 0 2675 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2817
transform 1 0 2633 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2818
transform 1 0 2574 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2819
transform 1 0 2304 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2820
transform 1 0 2231 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2821
transform 1 0 2179 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2822
transform 1 0 2518 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2823
transform 1 0 2672 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2824
transform 1 0 2725 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2825
transform 1 0 2652 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2826
transform 1 0 2587 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2827
transform 1 0 2719 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2828
transform 1 0 2669 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2829
transform 1 0 2621 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2830
transform 1 0 2562 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2831
transform 1 0 2292 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2832
transform 1 0 2225 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2833
transform 1 0 2173 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2834
transform 1 0 2567 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2835
transform 1 0 2663 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2836
transform 1 0 2627 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2837
transform 1 0 2568 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2838
transform 1 0 2298 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2839
transform 1 0 2573 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2840
transform 1 0 2617 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2841
transform 1 0 2605 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2842
transform 1 0 2707 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2843
transform 1 0 2569 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2844
transform 1 0 2634 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2845
transform 1 0 2713 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2846
transform 1 0 2660 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2847
transform 1 0 2506 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2848
transform 1 0 2362 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2849
transform 1 0 2080 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2850
transform 1 0 1894 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2851
transform 1 0 1687 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2852
transform 1 0 1732 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2853
transform 1 0 1822 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2854
transform 1 0 1858 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2855
transform 1 0 1940 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2856
transform 1 0 1903 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2857
transform 1 0 1588 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2858
transform 1 0 1600 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2859
transform 1 0 1810 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2860
transform 1 0 1846 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2861
transform 1 0 1934 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2862
transform 1 0 1897 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2863
transform 1 0 1884 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2864
transform 1 0 1789 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2865
transform 1 0 1933 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2866
transform 1 0 1801 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2867
transform 1 0 1801 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2868
transform 1 0 1835 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2869
transform 1 0 1457 0 1 732
box 0 0 3 6
use FEEDTHRU  F-2870
transform 1 0 1594 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2871
transform 1 0 1678 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2872
transform 1 0 1816 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2873
transform 1 0 1852 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2874
transform 1 0 1942 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2875
transform 1 0 2026 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2876
transform 1 0 1948 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2877
transform 1 0 1996 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2878
transform 1 0 2042 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2879
transform 1 0 2017 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2880
transform 1 0 2004 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2881
transform 1 0 2377 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2882
transform 1 0 2065 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2883
transform 1 0 2521 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2884
transform 1 0 2509 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2885
transform 1 0 2495 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2886
transform 1 0 1960 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2887
transform 1 0 2002 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2888
transform 1 0 2048 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2889
transform 1 0 1969 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2890
transform 1 0 1819 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2891
transform 1 0 1932 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2892
transform 1 0 1957 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2893
transform 1 0 1988 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2894
transform 1 0 2353 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2895
transform 1 0 2329 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2896
transform 1 0 2303 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2897
transform 1 0 1841 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2898
transform 1 0 1997 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2899
transform 1 0 1949 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2900
transform 1 0 1920 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2901
transform 1 0 2160 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2902
transform 1 0 1685 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2903
transform 1 0 1726 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2904
transform 1 0 1975 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2905
transform 1 0 2191 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2906
transform 1 0 2221 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2907
transform 1 0 1871 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2908
transform 1 0 1835 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2909
transform 1 0 1991 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2910
transform 1 0 1943 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2911
transform 1 0 1914 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2912
transform 1 0 1782 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2913
transform 1 0 1679 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2914
transform 1 0 2268 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2915
transform 1 0 2154 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2916
transform 1 0 2171 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2917
transform 1 0 2213 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2918
transform 1 0 2549 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2919
transform 1 0 2262 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2920
transform 1 0 2556 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2921
transform 1 0 2609 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2922
transform 1 0 2645 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2923
transform 1 0 1864 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2924
transform 1 0 1834 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2925
transform 1 0 1870 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2926
transform 1 0 1952 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2927
transform 1 0 1909 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2928
transform 1 0 1896 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2929
transform 1 0 1801 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2930
transform 1 0 1957 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2931
transform 1 0 1807 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2932
transform 1 0 1831 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2933
transform 1 0 1829 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2934
transform 1 0 1823 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2935
transform 1 0 1985 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2936
transform 1 0 1937 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2937
transform 1 0 1876 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2938
transform 1 0 1964 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2939
transform 1 0 1933 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2940
transform 1 0 1908 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2941
transform 1 0 1893 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2942
transform 1 0 1738 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2943
transform 1 0 1691 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2944
transform 1 0 2106 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2945
transform 1 0 1938 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2946
transform 1 0 1744 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2947
transform 1 0 1703 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2948
transform 1 0 1800 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2949
transform 1 0 1915 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2950
transform 1 0 1958 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2951
transform 1 0 1921 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2952
transform 1 0 1927 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2953
transform 1 0 1902 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2954
transform 1 0 1795 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2955
transform 1 0 1951 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2956
transform 1 0 2688 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2957
transform 1 0 2743 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2958
transform 1 0 2690 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2959
transform 1 0 2530 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2960
transform 1 0 2503 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2961
transform 1 0 2676 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2962
transform 1 0 2599 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2963
transform 1 0 2743 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2964
transform 1 0 2197 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2965
transform 1 0 2101 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2966
transform 1 0 1711 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-2967
transform 1 0 1600 0 1 901
box 0 0 3 6
use FEEDTHRU  F-2968
transform 1 0 1900 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2969
transform 1 0 1982 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2970
transform 1 0 1951 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2971
transform 1 0 1926 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-2972
transform 1 0 2201 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2973
transform 1 0 2513 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2974
transform 1 0 2543 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2975
transform 1 0 2531 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2976
transform 1 0 2575 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2977
transform 1 0 2495 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2978
transform 1 0 2561 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2979
transform 1 0 2597 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-2980
transform 1 0 2532 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-2981
transform 1 0 2244 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-2982
transform 1 0 2201 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-2983
transform 1 0 2032 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-2984
transform 1 0 1866 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-2985
transform 1 0 1753 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-2986
transform 1 0 1560 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-2987
transform 1 0 2633 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-2988
transform 1 0 2537 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-2989
transform 1 0 2525 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-2990
transform 1 0 2569 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-2991
transform 1 0 2575 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-2992
transform 1 0 2671 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-2993
transform 1 0 2527 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-2994
transform 1 0 2131 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2995
transform 1 0 2138 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-2996
transform 1 0 2470 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-2997
transform 1 0 2326 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-2998
transform 1 0 2185 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-2999
transform 1 0 2100 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3000
transform 1 0 2521 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3001
transform 1 0 2563 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3002
transform 1 0 2563 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3003
transform 1 0 2557 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3004
transform 1 0 2513 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3005
transform 1 0 2513 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3006
transform 1 0 1741 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3007
transform 1 0 1842 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3008
transform 1 0 1924 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3009
transform 1 0 2195 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3010
transform 1 0 2232 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3011
transform 1 0 2268 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3012
transform 1 0 2501 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3013
transform 1 0 2573 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3014
transform 1 0 2519 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3015
transform 1 0 2501 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3016
transform 1 0 2551 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3017
transform 1 0 1860 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3018
transform 1 0 1990 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3019
transform 1 0 2593 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3020
transform 1 0 2737 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3021
transform 1 0 2623 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3022
transform 1 0 2611 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3023
transform 1 0 2682 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3024
transform 1 0 2697 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3025
transform 1 0 2475 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3026
transform 1 0 2384 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3027
transform 1 0 2251 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3028
transform 1 0 2067 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3029
transform 1 0 2604 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3030
transform 1 0 2687 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3031
transform 1 0 2573 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3032
transform 1 0 2555 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3033
transform 1 0 2599 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3034
transform 1 0 2611 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3035
transform 1 0 2725 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3036
transform 1 0 2581 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3037
transform 1 0 2670 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3038
transform 1 0 2737 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3039
transform 1 0 2684 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3040
transform 1 0 2069 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3041
transform 1 0 2190 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3042
transform 1 0 2022 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3043
transform 1 0 2033 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3044
transform 1 0 2099 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3045
transform 1 0 2387 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3046
transform 1 0 2423 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3047
transform 1 0 2449 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3048
transform 1 0 2467 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3049
transform 1 0 2023 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3050
transform 1 0 1879 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3051
transform 1 0 1980 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3052
transform 1 0 1799 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3053
transform 1 0 2178 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3054
transform 1 0 1992 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3055
transform 1 0 2063 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3056
transform 1 0 2117 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3057
transform 1 0 2363 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3058
transform 1 0 2369 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3059
transform 1 0 2419 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3060
transform 1 0 2437 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3061
transform 1 0 2017 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3062
transform 1 0 1873 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3063
transform 1 0 1974 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3064
transform 1 0 1999 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3065
transform 1 0 2024 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3066
transform 1 0 1948 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3067
transform 1 0 1900 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3068
transform 1 0 1918 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3069
transform 1 0 1654 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3070
transform 1 0 1618 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3071
transform 1 0 1882 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3072
transform 1 0 1876 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3073
transform 1 0 1924 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3074
transform 1 0 2000 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3075
transform 1 0 1981 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3076
transform 1 0 1956 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3077
transform 1 0 1837 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3078
transform 1 0 1491 0 1 732
box 0 0 3 6
use FEEDTHRU  F-3079
transform 1 0 1624 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3080
transform 1 0 2707 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3081
transform 1 0 2636 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3082
transform 1 0 2654 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3083
transform 1 0 2500 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3084
transform 1 0 2356 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3085
transform 1 0 1731 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3086
transform 1 0 1774 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3087
transform 1 0 1715 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3088
transform 1 0 2100 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3089
transform 1 0 1968 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3090
transform 1 0 2015 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3091
transform 1 0 2069 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3092
transform 1 0 1883 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3093
transform 1 0 1780 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3094
transform 1 0 1721 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3095
transform 1 0 1806 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3096
transform 1 0 1974 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3097
transform 1 0 2021 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3098
transform 1 0 2075 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3099
transform 1 0 1913 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3100
transform 1 0 1865 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3101
transform 1 0 2215 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3102
transform 1 0 2155 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3103
transform 1 0 1981 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3104
transform 1 0 1825 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3105
transform 1 0 1944 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3106
transform 1 0 1975 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3107
transform 1 0 2006 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3108
transform 1 0 1918 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3109
transform 1 0 1870 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3110
transform 1 0 1726 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3111
transform 1 0 2142 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3112
transform 1 0 2177 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3113
transform 1 0 2519 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3114
transform 1 0 2483 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3115
transform 1 0 2665 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3116
transform 1 0 2118 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3117
transform 1 0 2479 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3118
transform 1 0 2575 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3119
transform 1 0 2612 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3120
transform 1 0 2482 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3121
transform 1 0 2338 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3122
transform 1 0 2038 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3123
transform 1 0 2618 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3124
transform 1 0 2671 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3125
transform 1 0 2124 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3126
transform 1 0 2485 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3127
transform 1 0 2635 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3128
transform 1 0 2557 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3129
transform 1 0 2545 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3130
transform 1 0 2624 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3131
transform 1 0 2677 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3132
transform 1 0 2166 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3133
transform 1 0 2515 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3134
transform 1 0 2647 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3135
transform 1 0 2533 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3136
transform 1 0 2521 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3137
transform 1 0 2539 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3138
transform 1 0 2527 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3139
transform 1 0 2507 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3140
transform 1 0 2531 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3141
transform 1 0 1831 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3142
transform 1 0 1987 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3143
transform 1 0 2045 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3144
transform 1 0 1865 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3145
transform 1 0 1805 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3146
transform 1 0 1807 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3147
transform 1 0 1847 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3148
transform 1 0 1811 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3149
transform 1 0 2143 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3150
transform 1 0 2144 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3151
transform 1 0 2014 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3152
transform 1 0 1996 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3153
transform 1 0 1978 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3154
transform 1 0 2642 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3155
transform 1 0 2695 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3156
transform 1 0 2478 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3157
transform 1 0 2533 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3158
transform 1 0 2683 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3159
transform 1 0 2551 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3160
transform 1 0 2539 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3161
transform 1 0 2648 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3162
transform 1 0 2701 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3163
transform 1 0 2616 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3164
transform 1 0 2539 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3165
transform 1 0 2689 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3166
transform 1 0 2545 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3167
transform 1 0 2533 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3168
transform 1 0 1858 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3169
transform 1 0 2046 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3170
transform 1 0 2197 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3171
transform 1 0 1642 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3172
transform 1 0 1497 0 1 732
box 0 0 3 6
use FEEDTHRU  F-3173
transform 1 0 1636 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3174
transform 1 0 2047 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3175
transform 1 0 1894 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3176
transform 1 0 1942 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3177
transform 1 0 2054 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3178
transform 1 0 2023 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3179
transform 1 0 1956 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3180
transform 1 0 1991 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3181
transform 1 0 2051 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3182
transform 1 0 1853 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3183
transform 1 0 1710 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3184
transform 1 0 1997 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3185
transform 1 0 2057 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3186
transform 1 0 1859 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3187
transform 1 0 1817 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3188
transform 1 0 1813 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3189
transform 1 0 1813 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3190
transform 1 0 2003 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3191
transform 1 0 1597 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3192
transform 1 0 1707 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3193
transform 1 0 1762 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3194
transform 1 0 1697 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3195
transform 1 0 1603 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3196
transform 1 0 1713 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3197
transform 1 0 2011 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3198
transform 1 0 1843 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3199
transform 1 0 1968 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3200
transform 1 0 2002 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3201
transform 1 0 2110 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3202
transform 1 0 2080 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3203
transform 1 0 2600 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3204
transform 1 0 2611 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3205
transform 1 0 1846 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3206
transform 1 0 1984 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3207
transform 1 0 2026 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3208
transform 1 0 2074 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3209
transform 1 0 2576 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3210
transform 1 0 2269 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3211
transform 1 0 2136 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3212
transform 1 0 1852 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3213
transform 1 0 2467 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3214
transform 1 0 2453 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3215
transform 1 0 2471 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3216
transform 1 0 2485 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3217
transform 1 0 2533 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3218
transform 1 0 2413 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3219
transform 1 0 2112 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3220
transform 1 0 2161 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3221
transform 1 0 2204 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3222
transform 1 0 2035 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3223
transform 1 0 2066 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3224
transform 1 0 1954 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3225
transform 1 0 1906 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3226
transform 1 0 1870 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3227
transform 1 0 1708 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3228
transform 1 0 2041 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3229
transform 1 0 2078 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3230
transform 1 0 1960 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3231
transform 1 0 1924 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3232
transform 1 0 1864 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3233
transform 1 0 1690 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3234
transform 1 0 2047 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3235
transform 1 0 2434 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3236
transform 1 0 2320 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3237
transform 1 0 1996 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3238
transform 1 0 2464 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3239
transform 1 0 2071 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3240
transform 1 0 2077 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3241
transform 1 0 2046 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3242
transform 1 0 1969 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3243
transform 1 0 2125 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3244
transform 1 0 2407 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3245
transform 1 0 2413 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3246
transform 1 0 2333 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3247
transform 1 0 2345 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3248
transform 1 0 2177 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3249
transform 1 0 2105 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3250
transform 1 0 2028 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3251
transform 1 0 2112 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3252
transform 1 0 1967 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3253
transform 1 0 1858 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3254
transform 1 0 2126 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3255
transform 1 0 2119 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3256
transform 1 0 2058 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3257
transform 1 0 2251 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3258
transform 1 0 2161 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3259
transform 1 0 2389 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3260
transform 1 0 2389 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3261
transform 1 0 2321 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3262
transform 1 0 2279 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3263
transform 1 0 2165 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3264
transform 1 0 1900 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3265
transform 1 0 2075 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3266
transform 1 0 2130 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3267
transform 1 0 2094 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3268
transform 1 0 2135 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3269
transform 1 0 2497 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3270
transform 1 0 2509 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3271
transform 1 0 2665 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3272
transform 1 0 2509 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3273
transform 1 0 2491 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3274
transform 1 0 2503 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3275
transform 1 0 2659 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3276
transform 1 0 2497 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3277
transform 1 0 2238 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3278
transform 1 0 2659 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3279
transform 1 0 2606 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3280
transform 1 0 2458 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3281
transform 1 0 2314 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3282
transform 1 0 1990 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3283
transform 1 0 2485 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3284
transform 1 0 2471 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3285
transform 1 0 2489 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3286
transform 1 0 2639 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3287
transform 1 0 2603 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3288
transform 1 0 2550 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3289
transform 1 0 2059 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3290
transform 1 0 2072 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3291
transform 1 0 1966 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3292
transform 1 0 1918 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3293
transform 1 0 2065 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3294
transform 1 0 2010 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3295
transform 1 0 1891 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3296
transform 1 0 2059 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3297
transform 1 0 2339 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3298
transform 1 0 2357 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3299
transform 1 0 2189 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3300
transform 1 0 2141 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3301
transform 1 0 2106 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3302
transform 1 0 2148 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3303
transform 1 0 2087 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3304
transform 1 0 2114 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3305
transform 1 0 1990 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3306
transform 1 0 1936 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3307
transform 1 0 1816 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3308
transform 1 0 2107 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3309
transform 1 0 2052 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3310
transform 1 0 2071 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3311
transform 1 0 2131 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3312
transform 1 0 2359 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3313
transform 1 0 2353 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3314
transform 1 0 2237 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3315
transform 1 0 2255 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3316
transform 1 0 2120 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3317
transform 1 0 2113 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3318
transform 1 0 1860 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3319
transform 1 0 2034 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3320
transform 1 0 2075 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3321
transform 1 0 2123 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3322
transform 1 0 1925 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3323
transform 1 0 1787 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3324
transform 1 0 2040 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3325
transform 1 0 2081 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3326
transform 1 0 2129 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3327
transform 1 0 2075 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3328
transform 1 0 2195 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3329
transform 1 0 2323 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3330
transform 1 0 2347 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3331
transform 1 0 2101 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3332
transform 1 0 1963 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3333
transform 1 0 2034 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3334
transform 1 0 2095 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3335
transform 1 0 2090 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3336
transform 1 0 2058 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3337
transform 1 0 2087 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3338
transform 1 0 2135 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3339
transform 1 0 2117 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3340
transform 1 0 2201 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3341
transform 1 0 2317 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3342
transform 1 0 2329 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3343
transform 1 0 2095 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3344
transform 1 0 1933 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3345
transform 1 0 1909 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3346
transform 1 0 2040 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3347
transform 1 0 2101 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3348
transform 1 0 2096 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3349
transform 1 0 1903 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3350
transform 1 0 2077 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3351
transform 1 0 2197 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3352
transform 1 0 2287 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3353
transform 1 0 2182 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3354
transform 1 0 2224 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3355
transform 1 0 2252 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3356
transform 1 0 2203 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3357
transform 1 0 2272 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3358
transform 1 0 2416 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3359
transform 1 0 2552 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3360
transform 1 0 2239 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3361
transform 1 0 2335 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3362
transform 1 0 2260 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3363
transform 1 0 2410 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3364
transform 1 0 2348 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3365
transform 1 0 2209 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3366
transform 1 0 2130 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3367
transform 1 0 2365 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3368
transform 1 0 2527 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3369
transform 1 0 2443 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3370
transform 1 0 2431 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3371
transform 1 0 2435 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3372
transform 1 0 2453 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3373
transform 1 0 2549 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3374
transform 1 0 2381 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3375
transform 1 0 2172 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3376
transform 1 0 2184 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3377
transform 1 0 2159 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3378
transform 1 0 2128 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3379
transform 1 0 1960 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3380
transform 1 0 2254 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3381
transform 1 0 2380 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3382
transform 1 0 2258 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3383
transform 1 0 2240 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3384
transform 1 0 2128 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3385
transform 1 0 2188 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3386
transform 1 0 2140 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3387
transform 1 0 1912 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3388
transform 1 0 1927 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3389
transform 1 0 1557 0 1 732
box 0 0 3 6
use FEEDTHRU  F-3390
transform 1 0 2516 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3391
transform 1 0 2245 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3392
transform 1 0 2142 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3393
transform 1 0 2546 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3394
transform 1 0 2251 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3395
transform 1 0 2154 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3396
transform 1 0 2383 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3397
transform 1 0 2557 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3398
transform 1 0 2455 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3399
transform 1 0 2437 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3400
transform 1 0 1806 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3401
transform 1 0 1864 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3402
transform 1 0 1805 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3403
transform 1 0 2076 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3404
transform 1 0 1812 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3405
transform 1 0 1876 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3406
transform 1 0 1835 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3407
transform 1 0 2052 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3408
transform 1 0 1818 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3409
transform 1 0 1882 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3410
transform 1 0 1901 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3411
transform 1 0 2022 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3412
transform 1 0 2150 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3413
transform 1 0 2020 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3414
transform 1 0 1978 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3415
transform 1 0 1810 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3416
transform 1 0 1660 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3417
transform 1 0 2311 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3418
transform 1 0 2299 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3419
transform 1 0 2231 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3420
transform 1 0 2243 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3421
transform 1 0 2305 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3422
transform 1 0 2293 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3423
transform 1 0 2225 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3424
transform 1 0 1921 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3425
transform 1 0 2070 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3426
transform 1 0 2137 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3427
transform 1 0 2168 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3428
transform 1 0 2038 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3429
transform 1 0 2641 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3430
transform 1 0 2461 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3431
transform 1 0 2443 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3432
transform 1 0 2447 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3433
transform 1 0 1470 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-3434
transform 1 0 1633 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3435
transform 1 0 1467 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-3436
transform 1 0 1624 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3437
transform 1 0 1755 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3438
transform 1 0 1810 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3439
transform 1 0 1745 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3440
transform 1 0 1740 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3441
transform 1 0 1998 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3442
transform 1 0 2039 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3443
transform 1 0 2087 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3444
transform 1 0 1889 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3445
transform 1 0 1853 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3446
transform 1 0 1837 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3447
transform 1 0 1837 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3448
transform 1 0 1630 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3449
transform 1 0 1761 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3450
transform 1 0 1816 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3451
transform 1 0 1757 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3452
transform 1 0 1734 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3453
transform 1 0 2016 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3454
transform 1 0 2057 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3455
transform 1 0 2093 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3456
transform 1 0 1907 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3457
transform 1 0 2315 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3458
transform 1 0 2351 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3459
transform 1 0 2327 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3460
transform 1 0 2369 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3461
transform 1 0 1798 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3462
transform 1 0 1888 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3463
transform 1 0 2214 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3464
transform 1 0 2465 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3465
transform 1 0 2555 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3466
transform 1 0 2393 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3467
transform 1 0 2363 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3468
transform 1 0 2407 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3469
transform 1 0 2179 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3470
transform 1 0 2089 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3471
transform 1 0 2102 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3472
transform 1 0 2083 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3473
transform 1 0 2016 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3474
transform 1 0 1861 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3475
transform 1 0 2035 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3476
transform 1 0 1819 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3477
transform 1 0 1819 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3478
transform 1 0 1841 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3479
transform 1 0 1895 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3480
transform 1 0 2105 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3481
transform 1 0 2045 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3482
transform 1 0 2004 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3483
transform 1 0 1716 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3484
transform 1 0 1733 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3485
transform 1 0 1807 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3486
transform 1 0 1752 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3487
transform 1 0 1912 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3488
transform 1 0 1585 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3489
transform 1 0 1615 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3490
transform 1 0 1448 0 1 732
box 0 0 3 6
use FEEDTHRU  F-3491
transform 1 0 1978 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3492
transform 1 0 2108 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3493
transform 1 0 2089 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3494
transform 1 0 2022 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3495
transform 1 0 1867 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3496
transform 1 0 2041 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3497
transform 1 0 1825 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3498
transform 1 0 1825 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3499
transform 1 0 1847 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3500
transform 1 0 1901 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3501
transform 1 0 2111 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3502
transform 1 0 2051 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3503
transform 1 0 2010 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3504
transform 1 0 1722 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3505
transform 1 0 1739 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3506
transform 1 0 1804 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3507
transform 1 0 1749 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3508
transform 1 0 1621 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3509
transform 1 0 2171 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3510
transform 1 0 2166 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3511
transform 1 0 2514 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3512
transform 1 0 2591 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3513
transform 1 0 2627 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3514
transform 1 0 2447 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3515
transform 1 0 2417 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3516
transform 1 0 2557 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3517
transform 1 0 2564 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3518
transform 1 0 2422 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3519
transform 1 0 2278 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3520
transform 1 0 1930 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3521
transform 1 0 1840 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3522
transform 1 0 1578 0 1 732
box 0 0 3 6
use FEEDTHRU  F-3523
transform 1 0 2587 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3524
transform 1 0 2184 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3525
transform 1 0 2401 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3526
transform 1 0 2593 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3527
transform 1 0 2196 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3528
transform 1 0 2407 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3529
transform 1 0 2569 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3530
transform 1 0 2431 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3531
transform 1 0 2159 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3532
transform 1 0 2112 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3533
transform 1 0 2058 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3534
transform 1 0 2167 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3535
transform 1 0 2082 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3536
transform 1 0 1939 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3537
transform 1 0 2180 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3538
transform 1 0 2050 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3539
transform 1 0 2056 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3540
transform 1 0 1984 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3541
transform 1 0 1762 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3542
transform 1 0 2198 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3543
transform 1 0 2179 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3544
transform 1 0 2094 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3545
transform 1 0 1945 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3546
transform 1 0 2119 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3547
transform 1 0 2185 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3548
transform 1 0 2227 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3549
transform 1 0 2219 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3550
transform 1 0 2231 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3551
transform 1 0 2183 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3552
transform 1 0 2129 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3553
transform 1 0 2088 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3554
transform 1 0 1824 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3555
transform 1 0 1811 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3556
transform 1 0 1870 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3557
transform 1 0 2191 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3558
transform 1 0 2135 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3559
transform 1 0 1943 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3560
transform 1 0 2153 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3561
transform 1 0 2093 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3562
transform 1 0 2046 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3563
transform 1 0 1788 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3564
transform 1 0 1793 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3565
transform 1 0 2185 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3566
transform 1 0 1786 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3567
transform 1 0 1956 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3568
transform 1 0 2214 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3569
transform 1 0 2599 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3570
transform 1 0 2570 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3571
transform 1 0 2428 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3572
transform 1 0 2284 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3573
transform 1 0 1924 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3574
transform 1 0 2640 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3575
transform 1 0 2503 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3576
transform 1 0 2628 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3577
transform 1 0 2491 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3578
transform 1 0 2653 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3579
transform 1 0 2449 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3580
transform 1 0 2425 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3581
transform 1 0 2429 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3582
transform 1 0 2459 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3583
transform 1 0 2154 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3584
transform 1 0 2424 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3585
transform 1 0 2478 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3586
transform 1 0 2531 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3587
transform 1 0 2597 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3588
transform 1 0 2429 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3589
transform 1 0 2399 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3590
transform 1 0 2401 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3591
transform 1 0 2425 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3592
transform 1 0 2623 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3593
transform 1 0 2461 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3594
transform 1 0 2484 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3595
transform 1 0 2549 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3596
transform 1 0 2615 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3597
transform 1 0 2435 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3598
transform 1 0 2411 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3599
transform 1 0 2014 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3600
transform 1 0 2086 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3601
transform 1 0 2216 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3602
transform 1 0 2197 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3603
transform 1 0 2573 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3604
transform 1 0 2621 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3605
transform 1 0 2441 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3606
transform 1 0 2405 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3607
transform 1 0 2395 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3608
transform 1 0 2413 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3609
transform 1 0 1936 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3610
transform 1 0 2296 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3611
transform 1 0 2452 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3612
transform 1 0 2594 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3613
transform 1 0 2653 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3614
transform 1 0 2526 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3615
transform 1 0 2467 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3616
transform 1 0 2629 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3617
transform 1 0 2419 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3618
transform 1 0 2088 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3619
transform 1 0 2149 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3620
transform 1 0 2156 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3621
transform 1 0 2026 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3622
transform 1 0 1915 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3623
transform 1 0 2071 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3624
transform 1 0 1843 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3625
transform 1 0 1843 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3626
transform 1 0 1889 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3627
transform 1 0 1931 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3628
transform 1 0 2147 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3629
transform 1 0 2099 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3630
transform 1 0 2052 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3631
transform 1 0 1746 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3632
transform 1 0 1751 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3633
transform 1 0 1822 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3634
transform 1 0 1773 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3635
transform 1 0 2155 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3636
transform 1 0 2162 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3637
transform 1 0 2032 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3638
transform 1 0 1954 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3639
transform 1 0 2148 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3640
transform 1 0 2215 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3641
transform 1 0 2227 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3642
transform 1 0 2149 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3643
transform 1 0 2227 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3644
transform 1 0 2281 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3645
transform 1 0 2297 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3646
transform 1 0 2273 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3647
transform 1 0 2267 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3648
transform 1 0 2165 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3649
transform 1 0 2118 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3650
transform 1 0 1968 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3651
transform 1 0 1829 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3652
transform 1 0 1888 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3653
transform 1 0 2371 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3654
transform 1 0 2393 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3655
transform 1 0 2417 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3656
transform 1 0 2591 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3657
transform 1 0 2543 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3658
transform 1 0 2472 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3659
transform 1 0 2142 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3660
transform 1 0 2141 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3661
transform 1 0 2140 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3662
transform 1 0 2028 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3663
transform 1 0 2395 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3664
transform 1 0 2365 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3665
transform 1 0 2375 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3666
transform 1 0 2405 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3667
transform 1 0 1732 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3668
transform 1 0 1887 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3669
transform 1 0 1834 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3670
transform 1 0 1763 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3671
transform 1 0 1764 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3672
transform 1 0 2064 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3673
transform 1 0 1654 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3674
transform 1 0 1788 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3675
transform 1 0 1840 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3676
transform 1 0 1769 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3677
transform 1 0 1758 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3678
transform 1 0 2070 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3679
transform 1 0 2111 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3680
transform 1 0 2159 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3681
transform 1 0 1973 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3682
transform 1 0 2015 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3683
transform 1 0 1873 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3684
transform 1 0 1879 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3685
transform 1 0 2083 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3686
transform 1 0 1927 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3687
transform 1 0 2106 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3688
transform 1 0 2173 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3689
transform 1 0 2174 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3690
transform 1 0 2044 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3691
transform 1 0 1972 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3692
transform 1 0 1794 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3693
transform 1 0 1846 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3694
transform 1 0 1775 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3695
transform 1 0 1752 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3696
transform 1 0 2076 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3697
transform 1 0 2117 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3698
transform 1 0 2160 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3699
transform 1 0 2263 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3700
transform 1 0 2179 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3701
transform 1 0 2299 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3702
transform 1 0 2387 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3703
transform 1 0 2423 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3704
transform 1 0 2609 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3705
transform 1 0 2555 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3706
transform 1 0 2508 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3707
transform 1 0 2124 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3708
transform 1 0 2383 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3709
transform 1 0 1572 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-3710
transform 1 0 1822 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3711
transform 1 0 1986 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3712
transform 1 0 2068 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3713
transform 1 0 2099 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3714
transform 1 0 1575 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-3715
transform 1 0 1792 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3716
transform 1 0 1962 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3717
transform 1 0 1810 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3718
transform 1 0 1974 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3719
transform 1 0 2080 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3720
transform 1 0 2111 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3721
transform 1 0 2070 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3722
transform 1 0 2442 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3723
transform 1 0 2513 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3724
transform 1 0 2567 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3725
transform 1 0 1816 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3726
transform 1 0 1980 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3727
transform 1 0 2122 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3728
transform 1 0 2117 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3729
transform 1 0 2617 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3730
transform 1 0 2490 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3731
transform 1 0 2449 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3732
transform 1 0 2027 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3733
transform 1 0 1930 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3734
transform 1 0 1914 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3735
transform 1 0 1759 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3736
transform 1 0 1524 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-3737
transform 1 0 2316 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3738
transform 1 0 2179 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3739
transform 1 0 2083 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3740
transform 1 0 2159 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3741
transform 1 0 2113 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3742
transform 1 0 1951 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3743
transform 1 0 2335 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3744
transform 1 0 2521 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3745
transform 1 0 2371 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3746
transform 1 0 2220 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3747
transform 1 0 2563 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3748
transform 1 0 2540 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3749
transform 1 0 2386 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3750
transform 1 0 2233 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3751
transform 1 0 2339 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3752
transform 1 0 2501 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3753
transform 1 0 2261 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3754
transform 1 0 2333 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3755
transform 1 0 2441 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3756
transform 1 0 2321 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3757
transform 1 0 2178 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3758
transform 1 0 1950 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3759
transform 1 0 2003 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3760
transform 1 0 1966 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3761
transform 1 0 1920 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3762
transform 1 0 2291 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3763
transform 1 0 2327 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3764
transform 1 0 2417 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3765
transform 1 0 2297 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3766
transform 1 0 2208 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3767
transform 1 0 2768 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3768
transform 1 0 2538 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3769
transform 1 0 2411 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3770
transform 1 0 2381 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3771
transform 1 0 2377 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3772
transform 1 0 2401 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3773
transform 1 0 2603 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3774
transform 1 0 2585 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3775
transform 1 0 2544 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3776
transform 1 0 2136 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3777
transform 1 0 2153 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3778
transform 1 0 2185 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3779
transform 1 0 2070 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3780
transform 1 0 1867 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3781
transform 1 0 2617 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3782
transform 1 0 2443 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3783
transform 1 0 2556 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3784
transform 1 0 2441 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3785
transform 1 0 2274 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3786
transform 1 0 1986 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3787
transform 1 0 2051 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3788
transform 1 0 1996 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3789
transform 1 0 2453 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3790
transform 1 0 2321 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3791
transform 1 0 2285 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3792
transform 1 0 2275 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3793
transform 1 0 2287 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3794
transform 1 0 2297 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3795
transform 1 0 2243 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3796
transform 1 0 2263 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3797
transform 1 0 2137 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3798
transform 1 0 2308 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3799
transform 1 0 2446 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3800
transform 1 0 2588 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3801
transform 1 0 2647 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3802
transform 1 0 2580 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3803
transform 1 0 2431 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3804
transform 1 0 2605 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3805
transform 1 0 2377 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3806
transform 1 0 2347 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3807
transform 1 0 2351 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3808
transform 1 0 2375 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3809
transform 1 0 2585 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3810
transform 1 0 2567 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3811
transform 1 0 2526 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3812
transform 1 0 2118 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3813
transform 1 0 2135 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3814
transform 1 0 1933 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3815
transform 1 0 1942 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3816
transform 1 0 2302 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3817
transform 1 0 2440 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3818
transform 1 0 2582 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3819
transform 1 0 2623 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3820
transform 1 0 2586 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3821
transform 1 0 2419 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3822
transform 1 0 2599 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3823
transform 1 0 2365 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3824
transform 1 0 2335 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3825
transform 1 0 2345 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3826
transform 1 0 2369 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3827
transform 1 0 2579 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3828
transform 1 0 2561 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3829
transform 1 0 2520 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3830
transform 1 0 2275 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3831
transform 1 0 2510 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3832
transform 1 0 2236 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3833
transform 1 0 2299 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3834
transform 1 0 2256 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3835
transform 1 0 2341 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3836
transform 1 0 2491 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3837
transform 1 0 2293 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3838
transform 1 0 2269 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3839
transform 1 0 2273 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3840
transform 1 0 2315 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3841
transform 1 0 2365 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3842
transform 1 0 2262 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3843
transform 1 0 2381 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3844
transform 1 0 2136 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3845
transform 1 0 1776 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3846
transform 1 0 2341 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3847
transform 1 0 2371 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3848
transform 1 0 2611 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3849
transform 1 0 2437 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3850
transform 1 0 2622 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3851
transform 1 0 2233 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3852
transform 1 0 2281 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3853
transform 1 0 2293 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3854
transform 1 0 2239 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3855
transform 1 0 2233 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3856
transform 1 0 2311 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3857
transform 1 0 2244 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3858
transform 1 0 2293 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3859
transform 1 0 2324 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3860
transform 1 0 2189 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3861
transform 1 0 2177 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3862
transform 1 0 2167 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3863
transform 1 0 2173 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3864
transform 1 0 2233 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3865
transform 1 0 2178 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3866
transform 1 0 1975 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3867
transform 1 0 2137 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3868
transform 1 0 1849 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3869
transform 1 0 1849 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3870
transform 1 0 2107 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3871
transform 1 0 1855 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3872
transform 1 0 1861 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3873
transform 1 0 1883 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3874
transform 1 0 1937 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3875
transform 1 0 2171 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3876
transform 1 0 2147 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3877
transform 1 0 2124 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3878
transform 1 0 2962 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3879
transform 1 0 2598 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3880
transform 1 0 2425 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3881
transform 1 0 2593 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3882
transform 1 0 2341 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3883
transform 1 0 1817 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3884
transform 1 0 1912 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3885
transform 1 0 1854 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3886
transform 1 0 1714 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-3887
transform 1 0 2275 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3888
transform 1 0 2485 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3889
transform 1 0 2359 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3890
transform 1 0 2316 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3891
transform 1 0 2539 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3892
transform 1 0 2462 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3893
transform 1 0 2356 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3894
transform 1 0 2212 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3895
transform 1 0 1894 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3896
transform 1 0 2251 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3897
transform 1 0 2239 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3898
transform 1 0 2267 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3899
transform 1 0 2303 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3900
transform 1 0 2507 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3901
transform 1 0 2489 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3902
transform 1 0 2376 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3903
transform 1 0 2034 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3904
transform 1 0 2057 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3905
transform 1 0 1889 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3906
transform 1 0 1942 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3907
transform 1 0 1902 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3908
transform 1 0 1871 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3909
transform 1 0 1948 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3910
transform 1 0 2525 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3911
transform 1 0 2507 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3912
transform 1 0 2448 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3913
transform 1 0 2064 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3914
transform 1 0 2279 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3915
transform 1 0 2161 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3916
transform 1 0 2137 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3917
transform 1 0 2171 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3918
transform 1 0 2147 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3919
transform 1 0 2219 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3920
transform 1 0 2195 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3921
transform 1 0 2160 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3922
transform 1 0 2155 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3923
transform 1 0 1999 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3924
transform 1 0 2190 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3925
transform 1 0 1993 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3926
transform 1 0 2279 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-3927
transform 1 0 2202 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3928
transform 1 0 1878 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3929
transform 1 0 2327 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-3930
transform 1 0 2225 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-3931
transform 1 0 2183 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3932
transform 1 0 2173 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3933
transform 1 0 2165 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3934
transform 1 0 2269 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3935
transform 1 0 2251 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3936
transform 1 0 2221 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3937
transform 1 0 2353 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3938
transform 1 0 2342 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3939
transform 1 0 2230 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3940
transform 1 0 2020 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3941
transform 1 0 1979 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3942
transform 1 0 2010 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-3943
transform 1 0 2298 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-3944
transform 1 0 2016 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-3945
transform 1 0 2146 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3946
transform 1 0 2081 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-3947
transform 1 0 2152 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-3948
transform 1 0 2098 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3949
transform 1 0 2002 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3950
transform 1 0 1774 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3951
transform 1 0 2104 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3952
transform 1 0 2228 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3953
transform 1 0 2257 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3954
transform 1 0 2208 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3955
transform 1 0 2287 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3956
transform 1 0 2292 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3957
transform 1 0 2377 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3958
transform 1 0 2384 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3959
transform 1 0 2326 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3960
transform 1 0 2206 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3961
transform 1 0 1876 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3962
transform 1 0 1804 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3963
transform 1 0 2304 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3964
transform 1 0 2533 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3965
transform 1 0 1524 0 1 732
box 0 0 3 6
use FEEDTHRU  F-3966
transform 1 0 1762 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3967
transform 1 0 1828 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3968
transform 1 0 2062 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3969
transform 1 0 2186 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3970
transform 1 0 2221 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3971
transform 1 0 1966 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3972
transform 1 0 2068 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3973
transform 1 0 2192 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3974
transform 1 0 2227 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3975
transform 1 0 2172 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3976
transform 1 0 2191 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3977
transform 1 0 2107 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3978
transform 1 0 2250 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3979
transform 1 0 2341 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3980
transform 1 0 2264 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-3981
transform 1 0 2212 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-3982
transform 1 0 2116 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-3983
transform 1 0 1804 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-3984
transform 1 0 1714 0 1 901
box 0 0 3 6
use FEEDTHRU  F-3985
transform 1 0 2315 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3986
transform 1 0 2311 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3987
transform 1 0 2323 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3988
transform 1 0 2587 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3989
transform 1 0 2395 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3990
transform 1 0 2610 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3991
transform 1 0 2641 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3992
transform 1 0 2309 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-3993
transform 1 0 2305 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-3994
transform 1 0 2317 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-3995
transform 1 0 2581 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-3996
transform 1 0 2389 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-3997
transform 1 0 2604 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-3998
transform 1 0 2635 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-3999
transform 1 0 1711 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-4000
transform 1 0 1890 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4001
transform 1 0 1954 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4002
transform 1 0 1847 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4003
transform 1 0 1812 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4004
transform 1 0 2190 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4005
transform 1 0 2207 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4006
transform 1 0 2291 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4007
transform 1 0 2183 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4008
transform 1 0 1765 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-4009
transform 1 0 2044 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4010
transform 1 0 2281 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4011
transform 1 0 2246 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4012
transform 1 0 2122 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4013
transform 1 0 2020 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4014
transform 1 0 2543 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4015
transform 1 0 2309 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4016
transform 1 0 2261 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4017
transform 1 0 2245 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4018
transform 1 0 2269 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4019
transform 1 0 2515 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4020
transform 1 0 2323 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4021
transform 1 0 2472 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4022
transform 1 0 2569 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4023
transform 1 0 2522 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4024
transform 1 0 2404 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4025
transform 1 0 2388 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4026
transform 1 0 2317 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4027
transform 1 0 2497 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4028
transform 1 0 2245 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4029
transform 1 0 2310 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4030
transform 1 0 2275 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4031
transform 1 0 2431 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4032
transform 1 0 2209 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4033
transform 1 0 2197 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4034
transform 1 0 2213 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4035
transform 1 0 2261 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4036
transform 1 0 2489 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4037
transform 1 0 2399 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4038
transform 1 0 2395 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4039
transform 1 0 2360 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4040
transform 1 0 2266 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4041
transform 1 0 2200 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4042
transform 1 0 1822 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4043
transform 1 0 1750 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4044
transform 1 0 1554 0 1 732
box 0 0 3 6
use FEEDTHRU  F-4045
transform 1 0 2537 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4046
transform 1 0 2502 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4047
transform 1 0 2094 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4048
transform 1 0 2105 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4049
transform 1 0 2309 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4050
transform 1 0 2226 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4051
transform 1 0 1938 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4052
transform 1 0 1943 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4053
transform 1 0 2002 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4054
transform 1 0 1908 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4055
transform 1 0 1747 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-4056
transform 1 0 2213 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4057
transform 1 0 2551 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4058
transform 1 0 2492 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4059
transform 1 0 2362 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4060
transform 1 0 2236 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4061
transform 1 0 1858 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4062
transform 1 0 2504 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4063
transform 1 0 2374 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4064
transform 1 0 2248 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4065
transform 1 0 1852 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4066
transform 1 0 1780 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4067
transform 1 0 2183 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4068
transform 1 0 2201 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4069
transform 1 0 1955 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4070
transform 1 0 2189 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4071
transform 1 0 2166 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4072
transform 1 0 1794 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4073
transform 1 0 1823 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4074
transform 1 0 1936 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4075
transform 1 0 1848 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4076
transform 1 0 1693 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-4077
transform 1 0 1464 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-4078
transform 1 0 2207 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4079
transform 1 0 1949 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4080
transform 1 0 1877 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4081
transform 1 0 1855 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4082
transform 1 0 1861 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4083
transform 1 0 2143 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4084
transform 1 0 1957 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4085
transform 1 0 2202 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4086
transform 1 0 2263 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4087
transform 1 0 2234 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4088
transform 1 0 2110 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4089
transform 1 0 2008 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4090
transform 1 0 2226 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4091
transform 1 0 1981 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4092
transform 1 0 2167 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4093
transform 1 0 2065 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4094
transform 1 0 1879 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4095
transform 1 0 2087 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4096
transform 1 0 2039 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4097
transform 1 0 2261 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4098
transform 1 0 2255 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4099
transform 1 0 2196 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4100
transform 1 0 1818 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4101
transform 1 0 1841 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4102
transform 1 0 1960 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4103
transform 1 0 1872 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4104
transform 1 0 2287 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4105
transform 1 0 2232 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4106
transform 1 0 1987 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4107
transform 1 0 2173 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4108
transform 1 0 1993 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4109
transform 1 0 1927 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4110
transform 1 0 2081 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4111
transform 1 0 2027 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4112
transform 1 0 2255 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4113
transform 1 0 2249 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4114
transform 1 0 1846 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4115
transform 1 0 2242 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4116
transform 1 0 2368 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4117
transform 1 0 2498 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4118
transform 1 0 2545 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4119
transform 1 0 2334 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4120
transform 1 0 2281 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4121
transform 1 0 2479 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4122
transform 1 0 2215 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4123
transform 1 0 2209 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4124
transform 1 0 2207 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4125
transform 1 0 2237 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4126
transform 1 0 2465 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4127
transform 1 0 2453 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4128
transform 1 0 2388 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4129
transform 1 0 2028 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4130
transform 1 0 2045 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4131
transform 1 0 2203 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4132
transform 1 0 1786 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4133
transform 1 0 1834 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4134
transform 1 0 2562 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4135
transform 1 0 2605 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4136
transform 1 0 2558 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4137
transform 1 0 2568 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4138
transform 1 0 2347 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4139
transform 1 0 2539 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4140
transform 1 0 2263 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4141
transform 1 0 2257 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4142
transform 1 0 2255 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4143
transform 1 0 2291 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4144
transform 1 0 2537 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4145
transform 1 0 2525 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4146
transform 1 0 2496 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4147
transform 1 0 2088 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4148
transform 1 0 2093 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4149
transform 1 0 2164 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4150
transform 1 0 2082 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4151
transform 1 0 2574 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4152
transform 1 0 2353 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4153
transform 1 0 2545 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4154
transform 1 0 2257 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4155
transform 1 0 2251 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4156
transform 1 0 2249 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4157
transform 1 0 2285 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4158
transform 1 0 2531 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4159
transform 1 0 2519 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4160
transform 1 0 2490 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4161
transform 1 0 2082 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4162
transform 1 0 2231 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4163
transform 1 0 2237 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4164
transform 1 0 1991 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4165
transform 1 0 1949 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4166
transform 1 0 1891 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4167
transform 1 0 2153 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4168
transform 1 0 2161 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4169
transform 1 0 2167 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4170
transform 1 0 2245 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4171
transform 1 0 2288 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4172
transform 1 0 2335 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4173
transform 1 0 2286 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4174
transform 1 0 2077 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4175
transform 1 0 2209 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4176
transform 1 0 2023 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4177
transform 1 0 1975 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4178
transform 1 0 2063 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4179
transform 1 0 2203 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4180
transform 1 0 1981 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4181
transform 1 0 1963 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4182
transform 1 0 1979 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4183
transform 1 0 2009 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4184
transform 1 0 2249 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4185
transform 1 0 2243 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4186
transform 1 0 2041 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4187
transform 1 0 2268 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4188
transform 1 0 2305 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4189
transform 1 0 2270 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4190
transform 1 0 2134 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4191
transform 1 0 2068 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4192
transform 1 0 1708 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4193
transform 1 0 2029 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4194
transform 1 0 2197 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4195
transform 1 0 1963 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4196
transform 1 0 1957 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4197
transform 1 0 1955 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4198
transform 1 0 2011 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4199
transform 1 0 2274 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4200
transform 1 0 2311 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4201
transform 1 0 2276 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4202
transform 1 0 2140 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4203
transform 1 0 2098 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4204
transform 1 0 1702 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4205
transform 1 0 2005 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4206
transform 1 0 2280 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4207
transform 1 0 2329 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4208
transform 1 0 2282 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4209
transform 1 0 2176 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4210
transform 1 0 2014 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4211
transform 1 0 1907 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4212
transform 1 0 1890 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4213
transform 1 0 2392 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4214
transform 1 0 2528 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4215
transform 1 0 2575 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4216
transform 1 0 2532 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4217
transform 1 0 2293 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4218
transform 1 0 2503 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4219
transform 1 0 1840 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4220
transform 1 0 2266 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4221
transform 1 0 2398 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4222
transform 1 0 2534 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4223
transform 1 0 2581 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4224
transform 1 0 2550 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4225
transform 1 0 2299 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4226
transform 1 0 2509 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4227
transform 1 0 2203 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4228
transform 1 0 2203 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4229
transform 1 0 2189 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4230
transform 1 0 2249 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4231
transform 1 0 2495 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4232
transform 1 0 1873 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4233
transform 1 0 1885 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4234
transform 1 0 2551 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4235
transform 1 0 2335 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4236
transform 1 0 2592 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4237
transform 1 0 2095 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4238
transform 1 0 2149 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4239
transform 1 0 2425 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4240
transform 1 0 2209 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4241
transform 1 0 2364 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4242
transform 1 0 2497 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4243
transform 1 0 2456 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4244
transform 1 0 2320 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4245
transform 1 0 2131 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4246
transform 1 0 2407 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4247
transform 1 0 2197 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4248
transform 1 0 2071 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4249
transform 1 0 2299 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4250
transform 1 0 2131 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4251
transform 1 0 2346 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4252
transform 1 0 2407 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4253
transform 1 0 2402 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4254
transform 1 0 2296 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4255
transform 1 0 2194 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4256
transform 1 0 1768 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4257
transform 1 0 2184 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4258
transform 1 0 2213 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4259
transform 1 0 2298 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4260
transform 1 0 2023 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4261
transform 1 0 2159 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4262
transform 1 0 2129 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4263
transform 1 0 2131 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4264
transform 1 0 2107 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4265
transform 1 0 2353 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4266
transform 1 0 2185 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4267
transform 1 0 2358 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4268
transform 1 0 2491 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4269
transform 1 0 2432 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4270
transform 1 0 2314 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4271
transform 1 0 2363 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4272
transform 1 0 2315 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4273
transform 1 0 2280 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4274
transform 1 0 1962 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4275
transform 1 0 1973 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4276
transform 1 0 2105 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4277
transform 1 0 2113 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4278
transform 1 0 2083 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4279
transform 1 0 2305 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4280
transform 1 0 2137 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4281
transform 1 0 2352 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4282
transform 1 0 2473 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4283
transform 1 0 1732 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4284
transform 1 0 1750 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4285
transform 1 0 2152 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4286
transform 1 0 2242 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4287
transform 1 0 2372 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4288
transform 1 0 2383 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4289
transform 1 0 2340 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4290
transform 1 0 2083 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4291
transform 1 0 2263 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4292
transform 1 0 2059 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4293
transform 1 0 2035 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4294
transform 1 0 2069 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4295
transform 1 0 2093 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4296
transform 1 0 2303 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4297
transform 1 0 2291 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4298
transform 1 0 2232 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4299
transform 1 0 1932 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4300
transform 1 0 1931 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4301
transform 1 0 1515 0 1 732
box 0 0 3 6
use FEEDTHRU  F-4302
transform 1 0 1726 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4303
transform 1 0 1738 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4304
transform 1 0 1798 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4305
transform 1 0 2230 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4306
transform 1 0 2350 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4307
transform 1 0 2486 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4308
transform 1 0 2509 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4309
transform 1 0 2412 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4310
transform 1 0 2203 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4311
transform 1 0 2419 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4312
transform 1 0 2137 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4313
transform 1 0 2149 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4314
transform 1 0 2147 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4315
transform 1 0 2195 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4316
transform 1 0 2435 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4317
transform 1 0 2387 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4318
transform 1 0 2346 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4319
transform 1 0 1998 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4320
transform 1 0 2015 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4321
transform 1 0 2086 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4322
transform 1 0 1792 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4323
transform 1 0 2224 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4324
transform 1 0 2344 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4325
transform 1 0 2468 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4326
transform 1 0 2503 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4327
transform 1 0 1648 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4328
transform 1 0 1672 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4329
transform 1 0 2062 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4330
transform 1 0 2146 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4331
transform 1 0 1684 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4332
transform 1 0 2086 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4333
transform 1 0 2182 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4334
transform 1 0 2306 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4335
transform 1 0 2514 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4336
transform 1 0 2257 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4337
transform 1 0 2443 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4338
transform 1 0 1902 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4339
transform 1 0 1925 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4340
transform 1 0 2238 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4341
transform 1 0 1920 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4342
transform 1 0 2093 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4343
transform 1 0 2101 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4344
transform 1 0 2077 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4345
transform 1 0 2329 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4346
transform 1 0 2155 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4347
transform 1 0 2376 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4348
transform 1 0 2425 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4349
transform 1 0 2390 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4350
transform 1 0 2254 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4351
transform 1 0 2170 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4352
transform 1 0 1744 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4353
transform 1 0 2450 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4354
transform 1 0 2308 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4355
transform 1 0 1985 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4356
transform 1 0 1907 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4357
transform 1 0 1897 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4358
transform 1 0 2292 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4359
transform 1 0 1774 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4360
transform 1 0 1756 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4361
transform 1 0 2188 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4362
transform 1 0 2302 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4363
transform 1 0 2438 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4364
transform 1 0 2479 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4365
transform 1 0 2394 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4366
transform 1 0 2191 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4367
transform 1 0 2401 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4368
transform 1 0 2101 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4369
transform 1 0 2107 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4370
transform 1 0 2099 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4371
transform 1 0 2165 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4372
transform 1 0 2405 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4373
transform 1 0 1933 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4374
transform 1 0 1903 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4375
transform 1 0 1937 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4376
transform 1 0 1979 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4377
transform 1 0 2227 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4378
transform 1 0 1909 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4379
transform 1 0 1921 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4380
transform 1 0 1919 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4381
transform 1 0 1951 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4382
transform 1 0 1951 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4383
transform 1 0 2239 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4384
transform 1 0 2035 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4385
transform 1 0 2318 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4386
transform 1 0 1810 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4387
transform 1 0 1786 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4388
transform 1 0 2218 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4389
transform 1 0 2332 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4390
transform 1 0 2474 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4391
transform 1 0 2515 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4392
transform 1 0 2520 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4393
transform 1 0 2215 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4394
transform 1 0 1654 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4395
transform 1 0 1666 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4396
transform 1 0 1648 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4397
transform 1 0 2038 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4398
transform 1 0 2158 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4399
transform 1 0 2300 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4400
transform 1 0 2323 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4401
transform 1 0 2328 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4402
transform 1 0 2017 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4403
transform 1 0 2221 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4404
transform 1 0 1897 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4405
transform 1 0 1909 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4406
transform 1 0 1901 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4407
transform 1 0 1961 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4408
transform 1 0 2225 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4409
transform 1 0 2219 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4410
transform 1 0 1678 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4411
transform 1 0 1612 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4412
transform 1 0 2032 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4413
transform 1 0 2152 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4414
transform 1 0 2294 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4415
transform 1 0 2317 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4416
transform 1 0 2009 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4417
transform 1 0 2011 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4418
transform 1 0 2017 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4419
transform 1 0 2164 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4420
transform 1 0 2050 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4421
transform 1 0 1618 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4422
transform 1 0 1684 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4423
transform 1 0 2338 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4424
transform 1 0 2480 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4425
transform 1 0 2527 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4426
transform 1 0 2544 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4427
transform 1 0 2245 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4428
transform 1 0 2473 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4429
transform 1 0 2143 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4430
transform 1 0 2155 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4431
transform 1 0 2141 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4432
transform 1 0 2219 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4433
transform 1 0 2483 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4434
transform 1 0 2483 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4435
transform 1 0 2454 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4436
transform 1 0 2097 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4437
transform 1 0 2281 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4438
transform 1 0 2044 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4439
transform 1 0 1606 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4440
transform 1 0 1672 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4441
transform 1 0 2225 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4442
transform 1 0 2231 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4443
transform 1 0 1967 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4444
transform 1 0 1895 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4445
transform 1 0 1915 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4446
transform 1 0 1891 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4447
transform 1 0 2443 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4448
transform 1 0 2448 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4449
transform 1 0 2179 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4450
transform 1 0 2371 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4451
transform 1 0 2041 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4452
transform 1 0 2071 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4453
transform 1 0 2033 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4454
transform 1 0 2105 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4455
transform 1 0 2123 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4456
transform 1 0 2201 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4457
transform 1 0 2471 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4458
transform 1 0 2471 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4459
transform 1 0 2460 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4460
transform 1 0 2040 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4461
transform 1 0 2108 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4462
transform 1 0 2125 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4463
transform 1 0 2461 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4464
transform 1 0 2239 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4465
transform 1 0 2538 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4466
transform 1 0 2521 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4467
transform 1 0 2243 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4468
transform 1 0 2237 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4469
transform 1 0 2220 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4470
transform 1 0 1830 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4471
transform 1 0 2065 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4472
transform 1 0 2257 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4473
transform 1 0 1927 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4474
transform 1 0 1939 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4475
transform 1 0 1913 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4476
transform 1 0 2119 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4477
transform 1 0 2467 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4478
transform 1 0 2233 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4479
transform 1 0 2113 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4480
transform 1 0 2143 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4481
transform 1 0 2117 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4482
transform 1 0 2207 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4483
transform 1 0 2477 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4484
transform 1 0 2477 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4485
transform 1 0 2466 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4486
transform 1 0 2358 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4487
transform 1 0 2369 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4488
transform 1 0 2393 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4489
transform 1 0 2129 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4490
transform 1 0 2045 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4491
transform 1 0 2053 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4492
transform 1 0 2035 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4493
transform 1 0 2389 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4494
transform 1 0 2364 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4495
transform 1 0 2375 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4496
transform 1 0 2399 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4497
transform 1 0 2141 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4498
transform 1 0 2051 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4499
transform 1 0 2041 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4500
transform 1 0 2029 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4501
transform 1 0 2377 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4502
transform 1 0 2167 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4503
transform 1 0 2454 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4504
transform 1 0 2461 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4505
transform 1 0 2420 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4506
transform 1 0 2284 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4507
transform 1 0 2164 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4508
transform 1 0 1720 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4509
transform 1 0 1756 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4510
transform 1 0 1563 0 1 732
box 0 0 3 6
use FEEDTHRU  F-4511
transform 1 0 2039 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4512
transform 1 0 2016 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4513
transform 1 0 2430 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4514
transform 1 0 2447 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4515
transform 1 0 2447 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4516
transform 1 0 2177 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4517
transform 1 0 2033 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4518
transform 1 0 2134 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4519
transform 1 0 2010 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4520
transform 1 0 1828 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-4521
transform 1 0 1554 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-4522
transform 1 0 2146 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4523
transform 1 0 2260 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4524
transform 1 0 2396 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4525
transform 1 0 2437 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4526
transform 1 0 2442 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4527
transform 1 0 2149 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4528
transform 1 0 2359 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4529
transform 1 0 2005 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4530
transform 1 0 2023 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4531
transform 1 0 2021 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4532
transform 1 0 2111 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4533
transform 1 0 2375 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4534
transform 1 0 2339 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4535
transform 1 0 2328 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4536
transform 1 0 1944 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4537
transform 1 0 1961 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4538
transform 1 0 2056 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4539
transform 1 0 1944 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4540
transform 1 0 1854 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4541
transform 1 0 1865 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4542
transform 1 0 1984 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4543
transform 1 0 2256 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4544
transform 1 0 2273 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4545
transform 1 0 2285 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4546
transform 1 0 2003 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4547
transform 1 0 1931 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4548
transform 1 0 1933 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4549
transform 1 0 1915 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4550
transform 1 0 2269 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4551
transform 1 0 2047 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4552
transform 1 0 1840 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-4553
transform 1 0 1485 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-4554
transform 1 0 1723 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-4555
transform 1 0 1878 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4556
transform 1 0 1972 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4557
transform 1 0 1853 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4558
transform 1 0 1836 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4559
transform 1 0 2244 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4560
transform 1 0 1482 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-4561
transform 1 0 1729 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-4562
transform 1 0 1884 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4563
transform 1 0 1978 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4564
transform 1 0 1859 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4565
transform 1 0 1842 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4566
transform 1 0 2250 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4567
transform 1 0 2267 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4568
transform 1 0 2273 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4569
transform 1 0 1997 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4570
transform 1 0 1925 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4571
transform 1 0 2111 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4572
transform 1 0 2125 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4573
transform 1 0 2095 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4574
transform 1 0 2455 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4575
transform 1 0 2119 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4576
transform 1 0 2089 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4577
transform 1 0 2449 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4578
transform 1 0 2221 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4579
transform 1 0 1991 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4580
transform 1 0 1981 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4581
transform 1 0 2077 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4582
transform 1 0 2047 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4583
transform 1 0 2413 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4584
transform 1 0 2411 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4585
transform 1 0 2394 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4586
transform 1 0 1992 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4587
transform 1 0 2009 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4588
transform 1 0 2110 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4589
transform 1 0 1998 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4590
transform 1 0 2435 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4591
transform 1 0 2418 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4592
transform 1 0 1991 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4593
transform 1 0 2104 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4594
transform 1 0 1980 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4595
transform 1 0 2400 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4596
transform 1 0 2417 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4597
transform 1 0 2429 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4598
transform 1 0 2153 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4599
transform 1 0 2057 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4600
transform 1 0 1488 0 1 732
box 0 0 3 6
use FEEDTHRU  F-4601
transform 1 0 1696 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4602
transform 1 0 1642 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4603
transform 1 0 1485 0 1 732
box 0 0 3 6
use FEEDTHRU  F-4604
transform 1 0 1702 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4605
transform 1 0 1624 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4606
transform 1 0 2074 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4607
transform 1 0 2200 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4608
transform 1 0 2330 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4609
transform 1 0 2359 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4610
transform 1 0 2370 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4611
transform 1 0 2053 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4612
transform 1 0 2275 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4613
transform 1 0 1921 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4614
transform 1 0 1945 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4615
transform 1 0 1943 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4616
transform 1 0 2015 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4617
transform 1 0 2297 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4618
transform 1 0 2303 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4619
transform 1 0 2286 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4620
transform 1 0 1866 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4621
transform 1 0 1877 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4622
transform 1 0 2419 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4623
transform 1 0 2430 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4624
transform 1 0 2119 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4625
transform 1 0 2341 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4626
transform 1 0 1975 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4627
transform 1 0 2005 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4628
transform 1 0 2003 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4629
transform 1 0 2099 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4630
transform 1 0 1581 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-4631
transform 1 0 1798 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-4632
transform 1 0 1968 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4633
transform 1 0 2092 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4634
transform 1 0 1804 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-4635
transform 1 0 2021 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4636
transform 1 0 2004 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4637
transform 1 0 2436 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4638
transform 1 0 2459 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4639
transform 1 0 2459 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4640
transform 1 0 2171 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4641
transform 1 0 2075 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4642
transform 1 0 2089 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4643
transform 1 0 2053 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4644
transform 1 0 1969 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4645
transform 1 0 1961 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4646
transform 1 0 2033 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4647
transform 1 0 2321 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4648
transform 1 0 2262 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4649
transform 1 0 2285 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4650
transform 1 0 2279 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4651
transform 1 0 2378 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4652
transform 1 0 2413 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4653
transform 1 0 2418 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4654
transform 1 0 2113 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4655
transform 1 0 2335 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4656
transform 1 0 1957 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4657
transform 1 0 1999 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4658
transform 1 0 1985 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4659
transform 1 0 2069 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4660
transform 1 0 2345 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4661
transform 1 0 2357 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4662
transform 1 0 2122 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4663
transform 1 0 1660 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4664
transform 1 0 2008 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4665
transform 1 0 1774 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-4666
transform 1 0 1926 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4667
transform 1 0 2050 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4668
transform 1 0 1913 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4669
transform 1 0 1896 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4670
transform 1 0 2322 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4671
transform 1 0 2345 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4672
transform 1 0 2333 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4673
transform 1 0 2057 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4674
transform 1 0 1973 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4675
transform 1 0 1993 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4676
transform 1 0 1945 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4677
transform 1 0 2323 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4678
transform 1 0 2101 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4679
transform 1 0 2400 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4680
transform 1 0 2080 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4681
transform 1 0 2194 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4682
transform 1 0 1768 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4683
transform 1 0 1696 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4684
transform 1 0 2158 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4685
transform 1 0 2272 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4686
transform 1 0 2414 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4687
transform 1 0 2455 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4688
transform 1 0 2460 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4689
transform 1 0 2143 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4690
transform 1 0 2365 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4691
transform 1 0 1987 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4692
transform 1 0 2444 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4693
transform 1 0 2485 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4694
transform 1 0 2502 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4695
transform 1 0 2173 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4696
transform 1 0 2395 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4697
transform 1 0 2011 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4698
transform 1 0 2059 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4699
transform 1 0 2039 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4700
transform 1 0 2135 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4701
transform 1 0 2423 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4702
transform 1 0 2429 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4703
transform 1 0 2412 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4704
transform 1 0 1974 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4705
transform 1 0 1997 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4706
transform 1 0 1597 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4707
transform 1 0 2056 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4708
transform 1 0 2170 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4709
transform 1 0 2312 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4710
transform 1 0 2347 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4711
transform 1 0 2304 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4712
transform 1 0 2333 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4713
transform 1 0 1950 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4714
transform 1 0 2074 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4715
transform 1 0 1937 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4716
transform 1 0 1908 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4717
transform 1 0 2352 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4718
transform 1 0 2021 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4719
transform 1 0 2309 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4720
transform 1 0 2327 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4721
transform 1 0 2310 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4722
transform 1 0 1872 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4723
transform 1 0 1895 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4724
transform 1 0 2038 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4725
transform 1 0 2508 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4726
transform 1 0 1992 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4727
transform 1 0 2116 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4728
transform 1 0 1985 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4729
transform 1 0 1956 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4730
transform 1 0 2406 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4731
transform 1 0 2423 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4732
transform 1 0 2411 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4733
transform 1 0 2123 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4734
transform 1 0 2027 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4735
transform 1 0 2047 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4736
transform 1 0 1999 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4737
transform 1 0 2383 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4738
transform 1 0 2161 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4739
transform 1 0 2496 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4740
transform 1 0 2467 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4741
transform 1 0 2426 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4742
transform 1 0 2278 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4743
transform 1 0 1636 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4744
transform 1 0 2092 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4745
transform 1 0 2206 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4746
transform 1 0 2354 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4747
transform 1 0 2389 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4748
transform 1 0 2424 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4749
transform 1 0 2095 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4750
transform 1 0 2311 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4751
transform 1 0 2065 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4752
transform 1 0 2357 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4753
transform 1 0 2063 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4754
transform 1 0 2026 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4755
transform 1 0 1883 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4756
transform 1 0 1848 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4757
transform 1 0 2408 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4758
transform 1 0 2449 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4759
transform 1 0 2484 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4760
transform 1 0 1497 0 1 11264
box 0 0 3 6
use FEEDTHRU  F-4761
transform 1 0 1768 0 1 11105
box 0 0 3 6
use FEEDTHRU  F-4762
transform 1 0 1938 0 1 10850
box 0 0 3 6
use FEEDTHRU  F-4763
transform 1 0 2062 0 1 10509
box 0 0 3 6
use FEEDTHRU  F-4764
transform 1 0 1919 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4765
transform 1 0 1884 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4766
transform 1 0 2334 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4767
transform 1 0 2351 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4768
transform 1 0 2339 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4769
transform 1 0 2045 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4770
transform 1 0 1949 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4771
transform 1 0 1914 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4772
transform 1 0 2370 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4773
transform 1 0 2393 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4774
transform 1 0 2381 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4775
transform 1 0 2081 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4776
transform 1 0 1997 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4777
transform 1 0 2017 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4778
transform 1 0 1969 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4779
transform 1 0 2347 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4780
transform 1 0 2125 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4781
transform 1 0 2466 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4782
transform 1 0 2431 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4783
transform 1 0 1714 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4784
transform 1 0 2176 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4785
transform 1 0 2290 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4786
transform 1 0 2248 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4787
transform 1 0 2134 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4788
transform 1 0 1666 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4789
transform 1 0 2340 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4790
transform 1 0 2363 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4791
transform 1 0 2351 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4792
transform 1 0 2051 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4793
transform 1 0 1967 0 1 6808
box 0 0 3 6
use FEEDTHRU  F-4794
transform 1 0 1987 0 1 6171
box 0 0 3 6
use FEEDTHRU  F-4795
transform 1 0 1939 0 1 5572
box 0 0 3 6
use FEEDTHRU  F-4796
transform 1 0 2317 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4797
transform 1 0 2089 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4798
transform 1 0 2436 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4799
transform 1 0 2401 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4800
transform 1 0 2366 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4801
transform 1 0 2218 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-4802
transform 1 0 2104 0 1 1571
box 0 0 3 6
use FEEDTHRU  F-4803
transform 1 0 2087 0 1 7369
box 0 0 3 6
use FEEDTHRU  F-4804
transform 1 0 2387 0 1 8006
box 0 0 3 6
use FEEDTHRU  F-4805
transform 1 0 2405 0 1 8585
box 0 0 3 6
use FEEDTHRU  F-4806
transform 1 0 2382 0 1 9128
box 0 0 3 6
use FEEDTHRU  F-4807
transform 1 0 1926 0 1 9631
box 0 0 3 6
use FEEDTHRU  F-4808
transform 1 0 1955 0 1 10092
box 0 0 3 6
use FEEDTHRU  F-4809
transform 1 0 1630 0 1 1182
box 0 0 3 6
use FEEDTHRU  F-4810
transform 1 0 1720 0 1 901
box 0 0 3 6
use FEEDTHRU  F-4811
transform 1 0 2336 0 1 2557
box 0 0 3 6
use FEEDTHRU  F-4812
transform 1 0 2371 0 1 3126
box 0 0 3 6
use FEEDTHRU  F-4813
transform 1 0 2406 0 1 3699
box 0 0 3 6
use FEEDTHRU  F-4814
transform 1 0 2059 0 1 4294
box 0 0 3 6
use FEEDTHRU  F-4815
transform 1 0 2287 0 1 4917
box 0 0 3 6
use FEEDTHRU  F-4816
transform 1 0 1903 0 1 5572
box 0 0 3 6
<< metal1 >>
rect 1423 683 1562 684
rect 1426 685 1595 686
rect 1430 687 1438 688
rect 1433 689 1450 690
rect 1440 691 1459 692
rect 1443 693 1487 694
rect 1446 695 1490 696
rect 1452 697 1598 698
rect 1455 699 1493 700
rect 1461 701 1499 702
rect 1464 703 1568 704
rect 1468 705 1517 706
rect 1471 707 1556 708
rect 1495 709 1630 710
rect 1507 711 1520 712
rect 1510 713 1514 714
rect 1525 713 1601 714
rect 1543 715 1607 716
rect 1546 717 1550 718
rect 1552 717 1619 718
rect 1558 719 1637 720
rect 1564 721 1633 722
rect 1579 723 1640 724
rect 1582 725 1623 726
rect 1603 727 1610 728
rect 1612 727 1626 728
rect 1615 729 1643 730
rect 1423 739 1683 740
rect 1423 741 1686 742
rect 1426 743 1722 744
rect 1426 745 1725 746
rect 1430 747 1710 748
rect 1430 749 1680 750
rect 1433 751 1650 752
rect 1433 753 1668 754
rect 1437 755 1590 756
rect 1436 757 2030 758
rect 1440 759 1689 760
rect 1439 761 1806 762
rect 1443 763 1716 764
rect 1443 765 1707 766
rect 1446 767 1923 768
rect 1446 769 1635 770
rect 1455 771 1962 772
rect 1464 773 1896 774
rect 1465 775 1662 776
rect 1468 777 1734 778
rect 1471 779 1782 780
rect 1474 781 1965 782
rect 1481 783 1542 784
rect 1484 785 1536 786
rect 1486 787 1704 788
rect 1489 789 1698 790
rect 1505 791 1598 792
rect 1507 793 1818 794
rect 1510 795 1746 796
rect 1511 797 1514 798
rect 1516 797 1728 798
rect 1477 799 1518 800
rect 1519 799 1794 800
rect 1523 801 1583 802
rect 1525 803 1764 804
rect 1543 805 2000 806
rect 1546 807 1833 808
rect 1547 809 1890 810
rect 1552 811 1878 812
rect 1555 813 1752 814
rect 1558 815 1929 816
rect 1561 817 1956 818
rect 1564 819 1758 820
rect 1567 821 1836 822
rect 1549 823 1569 824
rect 1550 825 1740 826
rect 1571 827 1640 828
rect 1579 829 1842 830
rect 1594 831 1821 832
rect 1458 833 1596 834
rect 1600 833 1959 834
rect 1601 835 1604 836
rect 1606 835 1908 836
rect 1609 837 1911 838
rect 1612 839 1938 840
rect 1615 841 1917 842
rect 1449 843 1617 844
rect 1450 845 1611 846
rect 1618 845 1987 846
rect 1452 847 1620 848
rect 1453 849 1605 850
rect 1622 849 2013 850
rect 1625 851 1800 852
rect 1492 853 1626 854
rect 1493 855 1953 856
rect 1629 857 1692 858
rect 1632 859 1770 860
rect 1495 861 1632 862
rect 1496 863 1830 864
rect 1636 865 1737 866
rect 1498 867 1638 868
rect 1642 867 2010 868
rect 1461 869 1644 870
rect 1462 871 1932 872
rect 1655 873 2033 874
rect 1673 875 1997 876
rect 1775 877 1968 878
rect 1787 879 1972 880
rect 1811 881 2016 882
rect 1847 883 1993 884
rect 1853 885 1990 886
rect 1859 887 2023 888
rect 1913 889 1920 890
rect 1925 889 2037 890
rect 1934 891 2040 892
rect 1940 893 2019 894
rect 1943 895 2007 896
rect 1974 897 2026 898
rect 1977 899 2004 900
rect 1417 908 1557 909
rect 1430 910 1644 911
rect 1443 912 1902 913
rect 1448 914 2289 915
rect 1450 916 2220 917
rect 1455 918 1575 919
rect 1459 920 1632 921
rect 1474 922 1527 923
rect 1477 924 1512 925
rect 1481 926 2064 927
rect 1484 928 2214 929
rect 1483 930 1569 931
rect 1486 932 1944 933
rect 1490 934 1854 935
rect 1493 936 2160 937
rect 1474 938 1494 939
rect 1502 938 2241 939
rect 1505 940 1515 941
rect 1505 942 2238 943
rect 1517 944 1533 945
rect 1520 946 1524 947
rect 1535 946 2112 947
rect 1541 948 2130 949
rect 1547 950 1911 951
rect 1550 952 2184 953
rect 1420 954 1551 955
rect 1586 954 1617 955
rect 1592 956 2277 957
rect 1601 958 1713 959
rect 1589 960 1602 961
rect 1496 962 1590 963
rect 1607 962 1674 963
rect 1613 964 1680 965
rect 1595 966 1680 967
rect 1595 968 2283 969
rect 1619 970 1884 971
rect 1619 972 1686 973
rect 1439 974 1686 975
rect 1438 976 1569 977
rect 1625 976 2346 977
rect 1625 978 1704 979
rect 1423 980 1704 981
rect 1424 982 1980 983
rect 1631 984 1722 985
rect 1637 986 2049 987
rect 1471 988 1638 989
rect 1643 988 1698 989
rect 1649 990 1674 991
rect 1649 992 1668 993
rect 1667 994 2375 995
rect 1676 996 1683 997
rect 1691 996 1866 997
rect 1697 998 1770 999
rect 1709 1000 1872 1001
rect 1436 1002 1710 1003
rect 1721 1002 1758 1003
rect 1724 1004 2046 1005
rect 1739 1006 2178 1007
rect 1727 1008 1740 1009
rect 1727 1010 2425 1011
rect 1745 1012 2094 1013
rect 1431 1014 1746 1015
rect 1751 1014 1824 1015
rect 1733 1016 1752 1017
rect 1688 1018 1734 1019
rect 1757 1018 1776 1019
rect 1465 1020 1776 1021
rect 1769 1022 2016 1023
rect 1426 1024 2016 1025
rect 1427 1026 1599 1027
rect 1781 1026 1854 1027
rect 1793 1028 2070 1029
rect 1793 1030 2365 1031
rect 1817 1032 2088 1033
rect 1462 1034 1818 1035
rect 1462 1036 2325 1037
rect 1820 1038 2217 1039
rect 1829 1040 2154 1041
rect 1763 1042 1830 1043
rect 1763 1044 2372 1045
rect 1832 1046 2166 1047
rect 1835 1048 2142 1049
rect 1787 1050 1836 1051
rect 1787 1052 1812 1053
rect 1661 1054 1812 1055
rect 1859 1054 2052 1055
rect 1859 1056 2023 1057
rect 1706 1058 2022 1059
rect 1877 1060 2100 1061
rect 1805 1062 1878 1063
rect 1715 1064 1806 1065
rect 1715 1066 2422 1067
rect 1889 1068 2172 1069
rect 1799 1070 1890 1071
rect 1799 1072 2368 1073
rect 1895 1074 2082 1075
rect 1895 1076 1968 1077
rect 1907 1078 2322 1079
rect 1571 1080 1908 1081
rect 1913 1080 2443 1081
rect 1913 1082 1929 1083
rect 1916 1084 2106 1085
rect 1919 1086 2256 1087
rect 1655 1088 1920 1089
rect 1433 1090 1656 1091
rect 1434 1092 2328 1093
rect 1922 1094 2253 1095
rect 1736 1096 1923 1097
rect 1441 1098 1737 1099
rect 1925 1098 2292 1099
rect 1925 1100 2030 1101
rect 1931 1102 2439 1103
rect 1841 1104 1932 1105
rect 1841 1106 2019 1107
rect 1934 1108 1944 1109
rect 1937 1110 2331 1111
rect 1937 1112 2033 1113
rect 1446 1114 2034 1115
rect 1445 1116 1662 1117
rect 1940 1116 2124 1117
rect 1952 1118 2340 1119
rect 1955 1120 2076 1121
rect 1610 1122 1956 1123
rect 1958 1122 2259 1123
rect 1961 1124 2196 1125
rect 1961 1126 2390 1127
rect 1964 1128 2058 1129
rect 1974 1130 2295 1131
rect 1604 1132 1974 1133
rect 1977 1132 2334 1133
rect 1986 1134 2250 1135
rect 1847 1136 1986 1137
rect 1847 1138 1972 1139
rect 1992 1138 2028 1139
rect 1991 1140 2000 1141
rect 1996 1142 2235 1143
rect 1997 1144 2349 1145
rect 2003 1146 2202 1147
rect 1989 1148 2004 1149
rect 2006 1148 2208 1149
rect 2009 1150 2359 1151
rect 1453 1152 2010 1153
rect 1452 1154 1581 1155
rect 2012 1154 2362 1155
rect 1634 1156 2013 1157
rect 2025 1156 2118 1157
rect 2039 1158 2139 1159
rect 2036 1160 2040 1161
rect 2036 1162 2432 1163
rect 2135 1164 2436 1165
rect 2189 1166 2446 1167
rect 2231 1168 2429 1169
rect 2297 1170 2353 1171
rect 2336 1172 2393 1173
rect 2342 1174 2356 1175
rect 2383 1174 2411 1175
rect 2386 1176 2408 1177
rect 2401 1178 2418 1179
rect 2404 1180 2415 1181
rect 1417 1189 1590 1190
rect 1417 1191 1968 1192
rect 1420 1193 2067 1194
rect 1427 1195 2283 1196
rect 1427 1197 2061 1198
rect 1434 1199 1740 1200
rect 1438 1201 2055 1202
rect 1438 1203 1656 1204
rect 1448 1205 2584 1206
rect 1448 1207 1836 1208
rect 1455 1209 2037 1210
rect 1455 1211 1572 1212
rect 1462 1213 2079 1214
rect 1466 1215 1632 1216
rect 1474 1217 2253 1218
rect 1473 1219 2157 1220
rect 1476 1221 2670 1222
rect 1480 1223 1521 1224
rect 1483 1225 1902 1226
rect 1483 1227 1590 1228
rect 1490 1229 1974 1230
rect 1471 1231 1974 1232
rect 1493 1233 1836 1234
rect 1502 1235 1887 1236
rect 1505 1237 1593 1238
rect 1514 1239 1584 1240
rect 1523 1241 1677 1242
rect 1529 1243 2550 1244
rect 1547 1245 1923 1246
rect 1550 1247 1971 1248
rect 1559 1249 2353 1250
rect 1577 1251 2325 1252
rect 1631 1253 2238 1254
rect 1643 1255 2422 1256
rect 1712 1257 2103 1258
rect 1781 1259 2016 1260
rect 1486 1261 2016 1262
rect 1487 1263 2058 1264
rect 1598 1265 2058 1266
rect 1793 1267 2226 1268
rect 1793 1269 2190 1270
rect 1757 1271 2190 1272
rect 1757 1273 2022 1274
rect 1829 1275 2368 1276
rect 1829 1277 2088 1278
rect 1685 1279 2088 1280
rect 1685 1281 2214 1282
rect 1841 1283 2643 1284
rect 1841 1285 1956 1286
rect 1847 1287 2244 1288
rect 1459 1289 1848 1290
rect 1459 1291 2064 1292
rect 1673 1293 2064 1294
rect 1574 1295 1674 1296
rect 1859 1295 2238 1296
rect 1859 1297 2010 1298
rect 1424 1299 2010 1300
rect 1424 1301 1500 1302
rect 1889 1301 2375 1302
rect 1595 1303 2376 1304
rect 1595 1305 2277 1306
rect 1889 1307 2100 1308
rect 1703 1309 2100 1310
rect 1703 1311 2112 1312
rect 1895 1313 2214 1314
rect 1895 1315 2049 1316
rect 1901 1317 1920 1318
rect 1420 1319 1920 1320
rect 1925 1319 2286 1320
rect 1865 1321 1926 1322
rect 1865 1323 2094 1324
rect 1637 1325 2094 1326
rect 1452 1327 1638 1328
rect 1452 1329 1908 1330
rect 1871 1331 1908 1332
rect 1727 1333 1872 1334
rect 1727 1335 2154 1336
rect 1751 1337 2154 1338
rect 1751 1339 2034 1340
rect 1613 1341 2034 1342
rect 1613 1343 2241 1344
rect 1931 1345 2280 1346
rect 1931 1347 2106 1348
rect 1943 1349 2304 1350
rect 1943 1351 2028 1352
rect 1949 1353 2544 1354
rect 1985 1355 2028 1356
rect 1763 1357 1986 1358
rect 1763 1359 2178 1360
rect 1715 1361 2178 1362
rect 1715 1363 2220 1364
rect 1787 1365 2220 1366
rect 1431 1367 1788 1368
rect 1431 1369 1506 1370
rect 1991 1369 2316 1370
rect 1991 1371 2636 1372
rect 2003 1373 2112 1374
rect 1775 1375 2004 1376
rect 1775 1377 2184 1378
rect 2012 1379 2025 1380
rect 2045 1379 2109 1380
rect 1607 1381 2046 1382
rect 2105 1381 2372 1382
rect 2117 1383 2382 1384
rect 1805 1385 2118 1386
rect 1805 1387 2070 1388
rect 1709 1389 2070 1390
rect 1709 1391 2130 1392
rect 2051 1393 2130 1394
rect 1619 1395 2052 1396
rect 1526 1397 1620 1398
rect 2123 1397 2352 1398
rect 1661 1399 2124 1400
rect 1556 1401 1662 1402
rect 2135 1401 2421 1402
rect 1667 1403 2136 1404
rect 1568 1405 1668 1406
rect 2138 1405 2310 1406
rect 2141 1407 2370 1408
rect 1913 1409 2142 1410
rect 1586 1411 1914 1412
rect 2183 1411 2393 1412
rect 2195 1413 2454 1414
rect 1769 1415 2196 1416
rect 1462 1417 1770 1418
rect 2198 1417 2217 1418
rect 2204 1419 2256 1420
rect 1961 1421 2256 1422
rect 1961 1423 2541 1424
rect 2207 1425 2448 1426
rect 1877 1427 2208 1428
rect 1877 1429 1884 1430
rect 1490 1431 1884 1432
rect 2231 1431 2478 1432
rect 1799 1433 2232 1434
rect 2249 1433 2502 1434
rect 1853 1435 2250 1436
rect 2258 1435 2508 1436
rect 2261 1437 2337 1438
rect 2267 1439 2640 1440
rect 2273 1441 2390 1442
rect 2288 1443 2496 1444
rect 2291 1445 2499 1446
rect 2291 1447 2633 1448
rect 2294 1449 2538 1450
rect 2297 1451 2514 1452
rect 1937 1453 2298 1454
rect 1817 1455 1938 1456
rect 1679 1457 1818 1458
rect 1580 1459 1680 1460
rect 2321 1459 2379 1460
rect 1997 1461 2322 1462
rect 1979 1463 1998 1464
rect 1811 1465 1980 1466
rect 1601 1467 1812 1468
rect 1441 1469 1602 1470
rect 1441 1471 1956 1472
rect 2327 1471 2565 1472
rect 2327 1473 2704 1474
rect 2330 1475 2466 1476
rect 2333 1477 2571 1478
rect 2075 1479 2334 1480
rect 1625 1481 2076 1482
rect 1532 1483 1626 1484
rect 1532 1485 2148 1486
rect 2339 1485 2547 1486
rect 2039 1487 2340 1488
rect 1649 1489 2040 1490
rect 1649 1491 1737 1492
rect 2342 1491 2520 1492
rect 2345 1493 2688 1494
rect 2345 1495 2580 1496
rect 2348 1497 2574 1498
rect 2355 1499 2526 1500
rect 2358 1501 2596 1502
rect 1469 1503 2358 1504
rect 2361 1503 2532 1504
rect 2364 1505 2425 1506
rect 2081 1507 2364 1508
rect 1445 1509 2082 1510
rect 1445 1511 2022 1512
rect 2234 1511 2424 1512
rect 2383 1513 2436 1514
rect 2386 1515 2608 1516
rect 2393 1517 2701 1518
rect 2399 1519 2446 1520
rect 2401 1521 2652 1522
rect 2404 1523 2646 1524
rect 2405 1525 2711 1526
rect 2407 1527 2623 1528
rect 2410 1529 2620 1530
rect 2414 1531 2667 1532
rect 2417 1533 2664 1534
rect 2417 1535 2715 1536
rect 2428 1537 2484 1538
rect 2431 1539 2487 1540
rect 2438 1541 2708 1542
rect 2442 1543 2505 1544
rect 2201 1545 2442 1546
rect 1823 1547 2202 1548
rect 1733 1549 1824 1550
rect 1733 1551 2160 1552
rect 1697 1553 2160 1554
rect 1434 1555 1698 1556
rect 2459 1555 2673 1556
rect 2489 1557 2587 1558
rect 2558 1559 2724 1560
rect 2561 1561 2721 1562
rect 2576 1563 2718 1564
rect 2601 1565 2629 1566
rect 2604 1567 2626 1568
rect 2675 1567 2694 1568
rect 2690 1569 2697 1570
rect 1424 1578 1518 1579
rect 1417 1580 1425 1581
rect 1427 1580 2175 1581
rect 1431 1582 2046 1583
rect 1445 1584 1932 1585
rect 1448 1586 1470 1587
rect 1448 1588 1620 1589
rect 1452 1590 1788 1591
rect 1452 1592 1866 1593
rect 1455 1594 1782 1595
rect 1466 1596 2319 1597
rect 1476 1598 2247 1599
rect 1469 1600 1477 1601
rect 1483 1600 1584 1601
rect 1485 1602 2124 1603
rect 1487 1604 1884 1605
rect 1502 1606 2370 1607
rect 1505 1608 1542 1609
rect 1532 1610 2901 1611
rect 1565 1612 2079 1613
rect 1577 1614 1608 1615
rect 1547 1616 1578 1617
rect 1473 1618 1548 1619
rect 1473 1620 2526 1621
rect 1625 1622 1656 1623
rect 1480 1624 1626 1625
rect 1643 1624 1887 1625
rect 1661 1626 1692 1627
rect 1631 1628 1662 1629
rect 1589 1630 1632 1631
rect 1679 1630 2779 1631
rect 1667 1632 1680 1633
rect 1709 1632 1740 1633
rect 1685 1634 1710 1635
rect 1745 1634 1782 1635
rect 1715 1636 1746 1637
rect 1751 1636 1800 1637
rect 1721 1638 1752 1639
rect 1703 1640 1722 1641
rect 1673 1642 1704 1643
rect 1649 1644 1674 1645
rect 1613 1646 1650 1647
rect 1571 1648 1614 1649
rect 1571 1650 2157 1651
rect 1763 1652 1788 1653
rect 1727 1654 1764 1655
rect 1697 1656 1728 1657
rect 1637 1658 1698 1659
rect 1595 1660 1638 1661
rect 1559 1662 1596 1663
rect 1523 1664 1560 1665
rect 1523 1666 2061 1667
rect 1805 1668 1884 1669
rect 1434 1670 1806 1671
rect 1817 1670 1854 1671
rect 1775 1672 1818 1673
rect 1601 1674 1776 1675
rect 1835 1674 1866 1675
rect 1835 1676 2868 1677
rect 1889 1678 2827 1679
rect 1841 1680 1890 1681
rect 1841 1682 2636 1683
rect 1931 1684 2292 1685
rect 1943 1686 2544 1687
rect 1895 1688 1944 1689
rect 1970 1688 2073 1689
rect 1973 1690 2046 1691
rect 1793 1692 1974 1693
rect 1455 1694 1794 1695
rect 1991 1694 2772 1695
rect 1937 1696 1992 1697
rect 1490 1698 1938 1699
rect 2021 1698 2124 1699
rect 1979 1700 2022 1701
rect 1417 1702 1980 1703
rect 2054 1702 2169 1703
rect 2066 1704 2163 1705
rect 2108 1706 2223 1707
rect 2177 1708 2292 1709
rect 1441 1710 2178 1711
rect 1441 1712 1848 1713
rect 1811 1714 1848 1715
rect 1757 1716 1812 1717
rect 2198 1716 2325 1717
rect 2102 1718 2199 1719
rect 2204 1718 2271 1719
rect 1529 1720 2205 1721
rect 1499 1722 1530 1723
rect 1499 1724 2742 1725
rect 2243 1726 2370 1727
rect 2153 1728 2244 1729
rect 2033 1730 2154 1731
rect 1955 1732 2034 1733
rect 1907 1734 1956 1735
rect 1859 1736 1908 1737
rect 1823 1738 1860 1739
rect 1459 1740 1824 1741
rect 1459 1742 2127 1743
rect 2261 1742 2412 1743
rect 2147 1744 2262 1745
rect 2063 1746 2148 1747
rect 1420 1748 2064 1749
rect 1420 1750 1914 1751
rect 1829 1752 1914 1753
rect 1769 1754 1830 1755
rect 1733 1756 1770 1757
rect 1427 1758 1734 1759
rect 2285 1758 2430 1759
rect 2165 1760 2286 1761
rect 2051 1762 2166 1763
rect 1488 1764 2052 1765
rect 2321 1764 2436 1765
rect 1492 1766 2322 1767
rect 2327 1766 2472 1767
rect 2207 1768 2328 1769
rect 2093 1770 2208 1771
rect 2093 1772 2841 1773
rect 2333 1774 2580 1775
rect 2219 1776 2334 1777
rect 2105 1778 2220 1779
rect 1466 1780 2106 1781
rect 2378 1780 2493 1781
rect 2381 1782 2526 1783
rect 2255 1784 2382 1785
rect 2171 1786 2256 1787
rect 2057 1788 2172 1789
rect 1985 1790 2058 1791
rect 1462 1792 1986 1793
rect 1462 1794 2025 1795
rect 2387 1794 2776 1795
rect 2423 1796 2580 1797
rect 2279 1798 2424 1799
rect 2279 1800 2769 1801
rect 2441 1802 2708 1803
rect 2303 1804 2442 1805
rect 2189 1806 2304 1807
rect 2141 1808 2190 1809
rect 2099 1810 2142 1811
rect 2003 1812 2100 1813
rect 1961 1814 2004 1815
rect 1925 1816 1962 1817
rect 1877 1818 1926 1819
rect 1431 1820 1878 1821
rect 2447 1820 2556 1821
rect 2309 1822 2448 1823
rect 2309 1824 2919 1825
rect 2459 1826 2616 1827
rect 2315 1828 2460 1829
rect 2486 1828 2631 1829
rect 2498 1830 2584 1831
rect 2501 1832 2655 1833
rect 2357 1834 2502 1835
rect 2213 1836 2358 1837
rect 2117 1838 2214 1839
rect 2117 1840 2394 1841
rect 2393 1842 2640 1843
rect 2489 1844 2640 1845
rect 2375 1846 2490 1847
rect 2249 1848 2376 1849
rect 2135 1850 2250 1851
rect 2069 1852 2136 1853
rect 1967 1854 2070 1855
rect 1919 1856 1968 1857
rect 1871 1858 1920 1859
rect 1434 1860 1872 1861
rect 2507 1860 2658 1861
rect 2363 1862 2508 1863
rect 2237 1864 2364 1865
rect 2237 1866 2643 1867
rect 2540 1868 2673 1869
rect 2543 1870 2908 1871
rect 2546 1872 2745 1873
rect 2549 1874 2748 1875
rect 2399 1876 2550 1877
rect 2267 1878 2400 1879
rect 2201 1880 2268 1881
rect 2075 1882 2202 1883
rect 2027 1884 2076 1885
rect 2027 1886 2838 1887
rect 2564 1888 2757 1889
rect 2570 1890 2831 1891
rect 2573 1892 2633 1893
rect 2417 1894 2574 1895
rect 2273 1896 2418 1897
rect 2159 1898 2274 1899
rect 2039 1900 2160 1901
rect 1495 1902 2040 1903
rect 2465 1902 2634 1903
rect 2465 1904 2871 1905
rect 2576 1906 2912 1907
rect 2591 1908 2670 1909
rect 2513 1910 2670 1911
rect 2595 1912 2788 1913
rect 2597 1914 2824 1915
rect 2601 1916 2821 1917
rect 2604 1918 2782 1919
rect 2453 1920 2604 1921
rect 2297 1922 2454 1923
rect 2195 1924 2298 1925
rect 2081 1926 2196 1927
rect 2081 1928 2112 1929
rect 2009 1930 2112 1931
rect 2009 1932 2130 1933
rect 2129 1934 2905 1935
rect 2607 1936 2800 1937
rect 2609 1938 2718 1939
rect 2619 1940 2812 1941
rect 2622 1942 2815 1943
rect 2477 1944 2622 1945
rect 2345 1946 2478 1947
rect 2225 1948 2346 1949
rect 2183 1950 2226 1951
rect 2087 1952 2184 1953
rect 2015 1954 2088 1955
rect 1997 1956 2016 1957
rect 1949 1958 1998 1959
rect 1901 1960 1950 1961
rect 1445 1962 1902 1963
rect 2625 1962 2818 1963
rect 2628 1964 2926 1965
rect 2483 1966 2628 1967
rect 2339 1968 2484 1969
rect 2339 1970 2704 1971
rect 2645 1972 2844 1973
rect 2651 1974 2850 1975
rect 2651 1976 2929 1977
rect 2663 1978 2862 1979
rect 2495 1980 2664 1981
rect 2351 1982 2496 1983
rect 2231 1984 2352 1985
rect 2231 1986 2709 1987
rect 2666 1988 2865 1989
rect 2586 1990 2667 1991
rect 2405 1992 2586 1993
rect 2405 1994 2922 1995
rect 2675 1996 2874 1997
rect 2519 1998 2676 1999
rect 2519 2000 2898 2001
rect 2687 2002 2697 2003
rect 2531 2004 2697 2005
rect 2504 2006 2532 2007
rect 2690 2006 2895 2007
rect 2693 2008 2892 2009
rect 2537 2010 2694 2011
rect 1438 2012 2538 2013
rect 1438 2014 2316 2015
rect 2700 2014 2703 2015
rect 2710 2014 2880 2015
rect 1583 2016 2712 2017
rect 2714 2016 2766 2017
rect 2561 2018 2715 2019
rect 2420 2020 2562 2021
rect 2720 2020 2727 2021
rect 2558 2022 2721 2023
rect 2723 2022 2883 2023
rect 2738 2024 2915 2025
rect 2762 2026 2834 2027
rect 1417 2035 2104 2036
rect 1420 2037 1990 2038
rect 1424 2039 3019 2040
rect 1427 2041 1900 2042
rect 1431 2043 1491 2044
rect 1432 2045 2338 2046
rect 1434 2047 1866 2048
rect 1436 2049 1960 2050
rect 1438 2051 2166 2052
rect 1443 2053 1854 2054
rect 1445 2055 1690 2056
rect 1448 2057 2199 2058
rect 1450 2059 1734 2060
rect 1452 2061 2175 2062
rect 1453 2063 1780 2064
rect 1455 2065 2290 2066
rect 1457 2067 1822 2068
rect 1462 2069 2709 2070
rect 1464 2071 2200 2072
rect 1466 2073 2100 2074
rect 1467 2075 2058 2076
rect 1469 2077 2098 2078
rect 1471 2079 2122 2080
rect 1473 2081 2022 2082
rect 1474 2083 1674 2084
rect 1476 2085 2152 2086
rect 1483 2087 1804 2088
rect 1485 2089 1588 2090
rect 1488 2091 2380 2092
rect 1492 2093 1932 2094
rect 1497 2095 1608 2096
rect 1499 2097 2014 2098
rect 1500 2099 1612 2100
rect 1502 2101 1978 2102
rect 1515 2103 2127 2104
rect 1486 2105 2128 2106
rect 1521 2107 1548 2108
rect 1523 2109 2779 2110
rect 1529 2111 1534 2112
rect 1541 2111 1552 2112
rect 1545 2113 1566 2114
rect 1557 2115 1572 2116
rect 1559 2117 1570 2118
rect 1563 2119 2163 2120
rect 1575 2121 1578 2122
rect 1583 2121 1600 2122
rect 1593 2123 1596 2124
rect 1613 2123 1630 2124
rect 1623 2125 2319 2126
rect 1429 2127 2320 2128
rect 1625 2129 1642 2130
rect 1631 2131 1648 2132
rect 1637 2133 1654 2134
rect 1643 2135 1660 2136
rect 1649 2137 1672 2138
rect 1655 2139 1684 2140
rect 1661 2141 1666 2142
rect 1677 2141 1776 2142
rect 1691 2143 1738 2144
rect 1692 2145 2020 2146
rect 1695 2147 1710 2148
rect 1697 2149 1720 2150
rect 1701 2151 1722 2152
rect 1703 2153 1726 2154
rect 1707 2155 1740 2156
rect 1727 2157 1774 2158
rect 1743 2159 1746 2160
rect 1749 2159 2223 2160
rect 1751 2161 1786 2162
rect 1761 2163 2670 2164
rect 1763 2165 1810 2166
rect 1769 2167 1816 2168
rect 1781 2169 1828 2170
rect 1787 2171 1852 2172
rect 1791 2173 2667 2174
rect 1793 2175 1834 2176
rect 1797 2177 2634 2178
rect 1799 2179 1840 2180
rect 1805 2181 1870 2182
rect 1811 2183 1846 2184
rect 1817 2185 1876 2186
rect 1823 2187 1858 2188
rect 1829 2189 1864 2190
rect 1835 2191 1882 2192
rect 1841 2193 1888 2194
rect 1847 2195 1936 2196
rect 1859 2197 1942 2198
rect 1871 2199 1954 2200
rect 1877 2201 1966 2202
rect 1883 2203 1912 2204
rect 1889 2205 1930 2206
rect 1893 2207 1974 2208
rect 1901 2209 1984 2210
rect 1905 2211 1986 2212
rect 1907 2213 1948 2214
rect 1913 2215 1924 2216
rect 1919 2217 2008 2218
rect 1925 2219 2002 2220
rect 1937 2221 1996 2222
rect 1943 2223 2056 2224
rect 1949 2225 2026 2226
rect 1955 2227 2068 2228
rect 1961 2229 2080 2230
rect 1971 2231 2118 2232
rect 1979 2233 2110 2234
rect 1991 2235 2116 2236
rect 1997 2237 2044 2238
rect 2003 2239 2050 2240
rect 2009 2241 2032 2242
rect 2015 2243 2146 2244
rect 2027 2245 2158 2246
rect 2033 2247 2164 2248
rect 2037 2249 2094 2250
rect 2045 2251 2176 2252
rect 2051 2253 2182 2254
rect 2061 2255 2640 2256
rect 2063 2257 2188 2258
rect 2069 2259 2194 2260
rect 2075 2261 2578 2262
rect 2081 2263 2602 2264
rect 2085 2265 2478 2266
rect 2087 2267 2218 2268
rect 2091 2269 2769 2270
rect 2105 2271 2230 2272
rect 2111 2273 2236 2274
rect 2129 2275 2242 2276
rect 2133 2277 3013 2278
rect 2139 2279 2472 2280
rect 2141 2281 2278 2282
rect 2147 2283 2917 2284
rect 2153 2285 2296 2286
rect 2159 2287 2302 2288
rect 2171 2289 2314 2290
rect 2177 2291 2284 2292
rect 2183 2293 2308 2294
rect 2189 2295 2968 2296
rect 2195 2297 2772 2298
rect 2072 2299 2197 2300
rect 1967 2301 2074 2302
rect 2201 2301 2332 2302
rect 2207 2303 2356 2304
rect 2211 2305 3119 2306
rect 2213 2307 2266 2308
rect 2219 2309 2368 2310
rect 2225 2311 2254 2312
rect 2231 2313 2344 2314
rect 2237 2315 2512 2316
rect 2243 2317 2374 2318
rect 2249 2319 2712 2320
rect 1459 2321 2251 2322
rect 1460 2323 2169 2324
rect 2039 2325 2170 2326
rect 2255 2325 2392 2326
rect 2259 2327 2382 2328
rect 2261 2329 2398 2330
rect 2267 2331 2362 2332
rect 2273 2333 2416 2334
rect 2279 2335 2428 2336
rect 2285 2337 2422 2338
rect 2291 2339 2905 2340
rect 2297 2341 2404 2342
rect 2303 2343 2440 2344
rect 2309 2345 2452 2346
rect 2310 2347 2919 2348
rect 2315 2349 2434 2350
rect 1517 2351 2317 2352
rect 2321 2351 2458 2352
rect 1679 2353 2323 2354
rect 2327 2353 2386 2354
rect 2333 2355 2476 2356
rect 2204 2357 2335 2358
rect 1495 2359 2206 2360
rect 2339 2359 2482 2360
rect 1446 2361 2341 2362
rect 2345 2361 2470 2362
rect 2349 2363 2412 2364
rect 2351 2365 2488 2366
rect 2357 2367 2464 2368
rect 2369 2369 2500 2370
rect 1441 2371 2371 2372
rect 2375 2371 2506 2372
rect 2246 2373 2377 2374
rect 2123 2375 2248 2376
rect 2387 2375 2542 2376
rect 2393 2377 2530 2378
rect 2399 2379 2536 2380
rect 2400 2381 2493 2382
rect 2363 2383 2494 2384
rect 2270 2385 2365 2386
rect 2135 2387 2272 2388
rect 2405 2387 2524 2388
rect 2409 2389 2776 2390
rect 2417 2391 2554 2392
rect 2423 2393 2566 2394
rect 2429 2395 2572 2396
rect 2435 2397 2871 2398
rect 2436 2399 3115 2400
rect 2441 2401 2584 2402
rect 2445 2403 2841 2404
rect 1493 2405 2842 2406
rect 2447 2407 2590 2408
rect 2453 2409 2596 2410
rect 2459 2411 2608 2412
rect 2324 2413 2461 2414
rect 2325 2415 2824 2416
rect 2465 2417 2838 2418
rect 2483 2419 2614 2420
rect 2489 2421 2827 2422
rect 2495 2423 3016 2424
rect 2507 2425 2662 2426
rect 2508 2427 2664 2428
rect 2517 2429 3058 2430
rect 2519 2431 2674 2432
rect 2525 2433 2680 2434
rect 2531 2435 2692 2436
rect 2547 2437 3055 2438
rect 2549 2439 2710 2440
rect 2555 2441 3025 2442
rect 2559 2443 3129 2444
rect 2585 2445 2752 2446
rect 2591 2447 2770 2448
rect 2603 2449 2776 2450
rect 2619 2451 3065 2452
rect 2625 2453 3062 2454
rect 2627 2455 2794 2456
rect 2630 2457 2797 2458
rect 2631 2459 2901 2460
rect 2637 2461 3122 2462
rect 2643 2463 3108 2464
rect 2649 2465 3105 2466
rect 2651 2467 2824 2468
rect 2654 2469 2926 2470
rect 2501 2471 2656 2472
rect 2667 2471 2898 2472
rect 2675 2473 2836 2474
rect 2685 2475 3112 2476
rect 2696 2477 2887 2478
rect 2537 2479 2698 2480
rect 2720 2479 2899 2480
rect 2561 2481 2722 2482
rect 2726 2481 2905 2482
rect 2727 2483 3028 2484
rect 2733 2485 2868 2486
rect 2741 2487 2869 2488
rect 2756 2489 2947 2490
rect 2757 2491 2908 2492
rect 2762 2493 2953 2494
rect 2597 2495 2764 2496
rect 2781 2495 2971 2496
rect 2609 2497 2782 2498
rect 2787 2497 2983 2498
rect 2615 2499 2788 2500
rect 2799 2499 2989 2500
rect 1439 2501 2800 2502
rect 2805 2501 3126 2502
rect 2811 2503 3001 2504
rect 2811 2505 2965 2506
rect 2814 2507 3004 2508
rect 2817 2509 3007 2510
rect 2820 2511 3010 2512
rect 2826 2513 2929 2514
rect 2738 2515 2929 2516
rect 2573 2517 2740 2518
rect 2830 2517 2920 2518
rect 2657 2519 2830 2520
rect 2833 2519 3022 2520
rect 2843 2521 3031 2522
rect 2847 2523 3101 2524
rect 2849 2525 3037 2526
rect 2853 2527 3098 2528
rect 2861 2529 3049 2530
rect 2864 2531 3052 2532
rect 2693 2533 2866 2534
rect 2873 2533 3080 2534
rect 2702 2535 2875 2536
rect 2543 2537 2704 2538
rect 2879 2537 3077 2538
rect 2744 2539 2881 2540
rect 2579 2541 2746 2542
rect 2891 2541 3092 2542
rect 2714 2543 2893 2544
rect 2621 2545 2716 2546
rect 2894 2545 3095 2546
rect 2911 2547 2944 2548
rect 2882 2549 2911 2550
rect 2747 2551 2884 2552
rect 2914 2551 2941 2552
rect 2921 2553 3074 2554
rect 2765 2555 2923 2556
rect 1420 2564 2260 2565
rect 1434 2566 1605 2567
rect 1436 2568 2152 2569
rect 1439 2570 2320 2571
rect 1441 2572 2178 2573
rect 1443 2574 2308 2575
rect 1450 2576 1774 2577
rect 1438 2578 1451 2579
rect 1457 2578 1948 2579
rect 1456 2580 1642 2581
rect 1464 2582 2182 2583
rect 1463 2584 2323 2585
rect 1474 2586 2116 2587
rect 1473 2588 1864 2589
rect 1486 2590 2794 2591
rect 1488 2592 1924 2593
rect 1427 2594 1923 2595
rect 1490 2596 1840 2597
rect 1491 2598 2050 2599
rect 1493 2600 2859 2601
rect 1497 2602 1594 2603
rect 1498 2604 2049 2605
rect 1500 2606 2401 2607
rect 1521 2608 3115 2609
rect 1526 2610 1546 2611
rect 1533 2612 1539 2613
rect 1569 2612 1581 2613
rect 1568 2614 1576 2615
rect 1563 2616 1575 2617
rect 1551 2618 1563 2619
rect 1550 2620 1558 2621
rect 1417 2622 1557 2623
rect 1587 2622 1593 2623
rect 1601 2622 2985 2623
rect 1611 2624 2442 2625
rect 1616 2626 3165 2627
rect 1629 2628 1635 2629
rect 1677 2628 1767 2629
rect 1676 2630 1684 2631
rect 1665 2632 1683 2633
rect 1653 2634 1665 2635
rect 1623 2636 1653 2637
rect 1689 2636 3031 2637
rect 1688 2638 1720 2639
rect 1695 2640 1713 2641
rect 1694 2642 1726 2643
rect 1701 2644 1725 2645
rect 1707 2646 1731 2647
rect 1706 2648 1738 2649
rect 1718 2650 1750 2651
rect 1736 2652 1744 2653
rect 1453 2654 1743 2655
rect 1748 2654 1780 2655
rect 1754 2656 1786 2657
rect 1761 2658 2991 2659
rect 1671 2660 1761 2661
rect 1659 2662 1671 2663
rect 1647 2664 1659 2665
rect 1772 2664 1834 2665
rect 1784 2666 1846 2667
rect 1797 2668 2913 2669
rect 1796 2670 1858 2671
rect 1832 2672 1852 2673
rect 1838 2674 1876 2675
rect 1844 2676 1972 2677
rect 1850 2678 1882 2679
rect 1856 2680 1900 2681
rect 1862 2682 1978 2683
rect 1880 2684 1894 2685
rect 1887 2686 3156 2687
rect 1886 2688 1930 2689
rect 1424 2690 1929 2691
rect 1892 2692 1906 2693
rect 1898 2694 1936 2695
rect 1904 2696 1942 2697
rect 1911 2698 2965 2699
rect 1910 2700 1954 2701
rect 1916 2702 1960 2703
rect 1934 2704 1966 2705
rect 1940 2706 3028 2707
rect 1946 2708 1996 2709
rect 1952 2710 1984 2711
rect 1958 2712 1990 2713
rect 1964 2714 3025 2715
rect 1970 2716 3016 2717
rect 1976 2718 2008 2719
rect 1982 2720 2002 2721
rect 1988 2722 3108 2723
rect 1994 2724 2032 2725
rect 2000 2726 2026 2727
rect 2006 2728 2038 2729
rect 2019 2730 2793 2731
rect 2018 2732 2044 2733
rect 2024 2734 2056 2735
rect 2030 2736 2086 2737
rect 2036 2738 2068 2739
rect 2042 2740 2080 2741
rect 1483 2742 2079 2743
rect 1446 2744 1483 2745
rect 2054 2744 3227 2745
rect 2061 2746 2931 2747
rect 2060 2748 2074 2749
rect 1432 2750 2073 2751
rect 1431 2752 1600 2753
rect 1598 2754 2944 2755
rect 2084 2756 2104 2757
rect 2097 2758 2103 2759
rect 2091 2760 2097 2761
rect 2090 2762 2110 2763
rect 1471 2764 2109 2765
rect 1470 2766 2067 2767
rect 2114 2766 2122 2767
rect 2120 2768 2128 2769
rect 1495 2770 2127 2771
rect 2150 2770 2158 2771
rect 2156 2772 2164 2773
rect 2162 2774 2206 2775
rect 2180 2776 2200 2777
rect 2187 2778 2223 2779
rect 2186 2780 3153 2781
rect 2196 2782 2232 2783
rect 2198 2784 2218 2785
rect 2204 2786 2254 2787
rect 2216 2788 3186 2789
rect 2229 2790 2259 2791
rect 2193 2792 2229 2793
rect 2192 2794 3108 2795
rect 2241 2796 2968 2797
rect 2240 2798 2554 2799
rect 2250 2800 2286 2801
rect 2252 2802 2548 2803
rect 2271 2804 2307 2805
rect 2270 2806 2578 2807
rect 2295 2808 2319 2809
rect 2294 2810 2326 2811
rect 2301 2812 2325 2813
rect 2316 2814 2352 2815
rect 2364 2814 2877 2815
rect 2334 2816 2364 2817
rect 2310 2818 2334 2819
rect 2370 2818 2406 2819
rect 2376 2820 2388 2821
rect 2340 2822 2376 2823
rect 2436 2822 2496 2823
rect 2451 2824 2920 2825
rect 2409 2826 2451 2827
rect 2403 2828 2409 2829
rect 2367 2830 2403 2831
rect 2460 2830 2502 2831
rect 2493 2832 2553 2833
rect 2433 2834 2493 2835
rect 1429 2836 2433 2837
rect 2499 2836 2547 2837
rect 2457 2838 2499 2839
rect 2415 2840 2457 2841
rect 2379 2842 2415 2843
rect 2378 2844 2386 2845
rect 2373 2846 2385 2847
rect 2337 2848 2373 2849
rect 2289 2850 2337 2851
rect 2529 2850 2577 2851
rect 2481 2852 2529 2853
rect 2439 2854 2481 2855
rect 2397 2856 2439 2857
rect 2361 2858 2397 2859
rect 2331 2860 2361 2861
rect 2283 2862 2331 2863
rect 2247 2864 2283 2865
rect 2246 2866 2518 2867
rect 2475 2868 2517 2869
rect 2474 2870 2917 2871
rect 2613 2872 3062 2873
rect 2601 2874 2613 2875
rect 2571 2876 2601 2877
rect 2523 2878 2571 2879
rect 1586 2880 2523 2881
rect 2655 2880 3230 2881
rect 2595 2882 2655 2883
rect 2594 2884 3190 2885
rect 2745 2886 2817 2887
rect 2691 2888 2745 2889
rect 2631 2890 2691 2891
rect 2787 2890 3241 2891
rect 2721 2892 2787 2893
rect 2667 2894 2721 2895
rect 2666 2896 3065 2897
rect 2796 2898 2889 2899
rect 2805 2900 2937 2901
rect 2739 2902 2805 2903
rect 2685 2904 2739 2905
rect 2211 2906 2685 2907
rect 2210 2908 2350 2909
rect 2313 2910 2349 2911
rect 2277 2912 2313 2913
rect 2276 2914 2512 2915
rect 2487 2916 2511 2917
rect 2445 2918 2487 2919
rect 1692 2920 2445 2921
rect 2811 2920 2943 2921
rect 1505 2922 2811 2923
rect 2826 2922 2907 2923
rect 2829 2924 2919 2925
rect 2763 2926 2829 2927
rect 2762 2928 3248 2929
rect 2835 2930 3027 2931
rect 2757 2932 2835 2933
rect 2697 2934 2757 2935
rect 2643 2936 2697 2937
rect 2642 2938 3234 2939
rect 2841 2940 3098 2941
rect 2775 2942 2841 2943
rect 2709 2944 2775 2945
rect 2637 2946 2709 2947
rect 2636 2948 2895 2949
rect 2847 2950 2955 2951
rect 2781 2952 2847 2953
rect 2727 2954 2781 2955
rect 2673 2956 2727 2957
rect 2619 2958 2673 2959
rect 2618 2960 3220 2961
rect 2853 2962 2949 2963
rect 2769 2964 2853 2965
rect 2703 2966 2769 2967
rect 2649 2968 2703 2969
rect 2589 2970 2649 2971
rect 2588 2972 3193 2973
rect 2865 2974 2961 2975
rect 2799 2976 2865 2977
rect 2733 2978 2799 2979
rect 2133 2980 2733 2981
rect 2132 2982 2140 2983
rect 2138 2984 2170 2985
rect 1467 2986 2169 2987
rect 1466 2988 1641 2989
rect 2868 2988 2967 2989
rect 2870 2990 3223 2991
rect 2883 2992 3060 2993
rect 2886 2994 3033 2995
rect 2898 2996 3015 2997
rect 2910 2998 3058 2999
rect 2823 3000 2910 3001
rect 2751 3002 2823 3003
rect 2679 3004 2751 3005
rect 2625 3006 2679 3007
rect 2583 3008 2625 3009
rect 2535 3010 2583 3011
rect 2534 3012 2898 3013
rect 2880 3014 3057 3015
rect 1803 3016 2880 3017
rect 1802 3018 1816 3019
rect 1502 3020 1815 3021
rect 2924 3020 3126 3021
rect 2928 3022 3072 3023
rect 2940 3024 3069 3025
rect 2946 3026 3087 3027
rect 2963 3028 3119 3029
rect 2972 3030 3101 3031
rect 2996 3032 3244 3033
rect 3000 3034 3141 3035
rect 3003 3036 3144 3037
rect 2508 3038 3003 3039
rect 3006 3038 3147 3039
rect 1791 3040 3006 3041
rect 1790 3042 1810 3043
rect 1808 3044 1822 3045
rect 1820 3046 1828 3047
rect 1826 3048 1870 3049
rect 1868 3050 2014 3051
rect 2012 3052 3013 3053
rect 3009 3054 3150 3055
rect 2892 3056 3009 3057
rect 2715 3058 2892 3059
rect 2661 3060 2715 3061
rect 2607 3062 2661 3063
rect 2559 3064 2607 3065
rect 2558 3066 2566 3067
rect 2541 3068 2565 3069
rect 2463 3070 2541 3071
rect 2421 3072 2463 3073
rect 1589 3074 2421 3075
rect 3018 3074 3159 3075
rect 3021 3076 3162 3077
rect 2904 3078 3021 3079
rect 3036 3078 3180 3079
rect 3044 3080 3168 3081
rect 3048 3082 3055 3083
rect 3051 3084 3177 3085
rect 2874 3086 3051 3087
rect 3073 3086 3214 3087
rect 2366 3088 3075 3089
rect 3076 3088 3217 3089
rect 2300 3090 3078 3091
rect 3079 3090 3112 3091
rect 2922 3092 3081 3093
rect 2970 3094 3111 3095
rect 3091 3096 3202 3097
rect 2952 3098 3093 3099
rect 3094 3098 3205 3099
rect 3104 3100 3183 3101
rect 2505 3102 3105 3103
rect 2469 3104 2505 3105
rect 2427 3106 2469 3107
rect 2391 3108 2427 3109
rect 2355 3110 2391 3111
rect 2343 3112 2355 3113
rect 2265 3114 2343 3115
rect 2235 3116 2265 3117
rect 1460 3118 2235 3119
rect 1459 3120 2289 3121
rect 3121 3120 3237 3121
rect 2982 3122 3123 3123
rect 3128 3122 3251 3123
rect 2988 3124 3129 3125
rect 1417 3133 1923 3134
rect 1420 3135 2049 3136
rect 1427 3137 1917 3138
rect 1431 3139 2388 3140
rect 1431 3141 2157 3142
rect 1441 3143 2303 3144
rect 1459 3145 1947 3146
rect 1463 3147 1689 3148
rect 1427 3149 1688 3150
rect 1450 3151 1463 3152
rect 1438 3153 1451 3154
rect 1438 3155 2613 3156
rect 1466 3157 1905 3158
rect 1468 3159 3038 3160
rect 1473 3161 2061 3162
rect 1485 3163 2283 3164
rect 1488 3165 2223 3166
rect 1491 3167 2115 3168
rect 1495 3169 2043 3170
rect 1482 3171 1495 3172
rect 1498 3171 2037 3172
rect 1502 3173 2073 3174
rect 1505 3175 2013 3176
rect 1507 3177 1569 3178
rect 1514 3179 1520 3180
rect 1526 3179 1532 3180
rect 1525 3181 1617 3182
rect 1528 3183 2502 3184
rect 1538 3185 1544 3186
rect 1562 3185 1568 3186
rect 1556 3187 1562 3188
rect 1478 3189 1556 3190
rect 1586 3189 2025 3190
rect 1580 3191 1586 3192
rect 1574 3193 1580 3194
rect 1475 3195 1574 3196
rect 1592 3195 1616 3196
rect 1601 3197 1605 3198
rect 1434 3199 1604 3200
rect 1434 3201 1613 3202
rect 1609 3203 3045 3204
rect 1658 3205 3075 3206
rect 1652 3207 1658 3208
rect 1694 3207 1700 3208
rect 1712 3207 3244 3208
rect 1706 3209 1712 3210
rect 1724 3209 2423 3210
rect 1723 3211 3248 3212
rect 1748 3213 1778 3214
rect 1736 3215 1748 3216
rect 1844 3215 1922 3216
rect 1802 3217 1844 3218
rect 1772 3219 1802 3220
rect 1742 3221 1772 3222
rect 1730 3223 1742 3224
rect 1424 3225 1730 3226
rect 1424 3227 1694 3228
rect 1862 3227 3153 3228
rect 1820 3229 1862 3230
rect 1819 3231 1827 3232
rect 1825 3233 1833 3234
rect 1796 3235 1832 3236
rect 1795 3237 1851 3238
rect 1790 3239 1850 3240
rect 1789 3241 1809 3242
rect 1807 3243 1839 3244
rect 1837 3245 1857 3246
rect 1873 3245 1881 3246
rect 1879 3247 1893 3248
rect 1868 3249 1892 3250
rect 1814 3251 1868 3252
rect 1784 3253 1814 3254
rect 1903 3253 1929 3254
rect 1915 3255 2793 3256
rect 1927 3257 1953 3258
rect 1621 3259 1952 3260
rect 1945 3261 1977 3262
rect 1975 3263 2001 3264
rect 1999 3265 2031 3266
rect 1482 3267 2030 3268
rect 2011 3269 2067 3270
rect 2023 3271 2091 3272
rect 2035 3273 2097 3274
rect 2041 3275 2103 3276
rect 2047 3277 2079 3278
rect 2054 3279 2066 3280
rect 2053 3281 2109 3282
rect 2059 3283 2121 3284
rect 2071 3285 2139 3286
rect 2080 3287 2880 3288
rect 2089 3289 2151 3290
rect 2095 3291 2181 3292
rect 2101 3293 2187 3294
rect 2107 3295 2175 3296
rect 2113 3297 2163 3298
rect 1598 3299 2162 3300
rect 1510 3301 1598 3302
rect 2119 3301 2667 3302
rect 2132 3303 3156 3304
rect 2131 3305 2211 3306
rect 2137 3307 2271 3308
rect 2149 3309 2217 3310
rect 2155 3311 2253 3312
rect 2173 3313 2229 3314
rect 1456 3315 2228 3316
rect 1456 3317 2178 3318
rect 2176 3319 2232 3320
rect 2179 3321 2235 3322
rect 2185 3323 2589 3324
rect 2194 3325 2286 3326
rect 2204 3327 3137 3328
rect 2203 3329 2265 3330
rect 2206 3331 2352 3332
rect 2209 3333 2259 3334
rect 2215 3335 2601 3336
rect 2221 3337 2565 3338
rect 2233 3339 2289 3340
rect 2240 3341 3190 3342
rect 2239 3343 2661 3344
rect 2198 3345 2660 3346
rect 2197 3347 2595 3348
rect 2251 3349 2343 3350
rect 2257 3351 2301 3352
rect 1441 3353 2300 3354
rect 2263 3355 2367 3356
rect 2269 3357 2307 3358
rect 2276 3359 3078 3360
rect 1886 3361 3077 3362
rect 1885 3363 1899 3364
rect 1897 3365 1911 3366
rect 1909 3367 1935 3368
rect 1933 3369 1959 3370
rect 1957 3371 1983 3372
rect 1589 3373 1982 3374
rect 2275 3373 2313 3374
rect 2281 3375 2331 3376
rect 2284 3377 2334 3378
rect 2287 3379 2337 3380
rect 2305 3381 2535 3382
rect 2311 3383 2898 3384
rect 2324 3385 2330 3386
rect 2192 3387 2324 3388
rect 1417 3389 2192 3390
rect 2335 3389 2547 3390
rect 2341 3391 2385 3392
rect 2354 3393 2663 3394
rect 2353 3395 2475 3396
rect 2365 3397 2499 3398
rect 2375 3399 2411 3400
rect 2363 3401 2375 3402
rect 2383 3401 2691 3402
rect 2396 3403 2895 3404
rect 2395 3405 2481 3406
rect 2434 3407 2496 3408
rect 2441 3409 2447 3410
rect 2405 3411 2441 3412
rect 1550 3413 2405 3414
rect 2468 3413 2498 3414
rect 2432 3415 2468 3416
rect 2420 3417 2432 3418
rect 2414 3419 2420 3420
rect 2413 3421 2511 3422
rect 2470 3423 2877 3424
rect 2473 3425 2571 3426
rect 2479 3427 2697 3428
rect 2126 3429 2696 3430
rect 2125 3431 2673 3432
rect 2504 3433 3186 3434
rect 2486 3435 2504 3436
rect 2450 3437 2486 3438
rect 2444 3439 2450 3440
rect 2438 3441 2444 3442
rect 2402 3443 2438 3444
rect 1500 3445 2402 3446
rect 2509 3445 3183 3446
rect 2528 3447 2546 3448
rect 2527 3449 2655 3450
rect 2533 3451 2577 3452
rect 2552 3453 3105 3454
rect 2551 3455 2583 3456
rect 2558 3457 3193 3458
rect 2557 3459 3108 3460
rect 2563 3461 2607 3462
rect 2569 3463 3199 3464
rect 2575 3465 3196 3466
rect 2581 3467 2649 3468
rect 2587 3469 2625 3470
rect 2599 3471 2964 3472
rect 2605 3473 2637 3474
rect 2611 3475 2643 3476
rect 2623 3477 3237 3478
rect 2629 3479 3241 3480
rect 2635 3481 2715 3482
rect 2647 3483 2721 3484
rect 2653 3485 2727 3486
rect 2665 3487 3119 3488
rect 2671 3489 2739 3490
rect 1970 3491 2738 3492
rect 1420 3493 1970 3494
rect 2684 3493 3116 3494
rect 1503 3495 2684 3496
rect 2689 3495 2745 3496
rect 2708 3497 3227 3498
rect 2707 3499 3251 3500
rect 2713 3501 2757 3502
rect 2719 3503 2751 3504
rect 2725 3505 2769 3506
rect 2743 3507 2799 3508
rect 2749 3509 2805 3510
rect 2755 3511 3189 3512
rect 2767 3513 3230 3514
rect 2774 3515 3171 3516
rect 2773 3517 2829 3518
rect 1940 3519 2828 3520
rect 1624 3521 1940 3522
rect 2791 3521 2823 3522
rect 2797 3523 2835 3524
rect 2803 3525 3220 3526
rect 2641 3527 3220 3528
rect 2821 3529 2847 3530
rect 2833 3531 2913 3532
rect 2845 3533 2865 3534
rect 2852 3535 2864 3536
rect 2870 3535 2885 3536
rect 2869 3537 3153 3538
rect 2875 3539 2925 3540
rect 2881 3541 2892 3542
rect 2888 3543 3074 3544
rect 2887 3545 2931 3546
rect 2893 3547 2937 3548
rect 2911 3549 2943 3550
rect 2918 3551 3156 3552
rect 2917 3553 2973 3554
rect 2923 3555 3006 3556
rect 2935 3557 2967 3558
rect 1470 3559 2966 3560
rect 1471 3561 2349 3562
rect 2347 3563 2409 3564
rect 2372 3565 2408 3566
rect 2360 3567 2372 3568
rect 2359 3569 2493 3570
rect 2491 3571 2619 3572
rect 2617 3573 2703 3574
rect 2701 3575 2763 3576
rect 2761 3577 3192 3578
rect 2944 3579 2961 3580
rect 2948 3581 3053 3582
rect 2947 3583 2985 3584
rect 2971 3585 3009 3586
rect 2977 3587 3015 3588
rect 2983 3589 3021 3590
rect 3002 3591 3041 3592
rect 3001 3593 3027 3594
rect 3013 3595 3165 3596
rect 3019 3597 3057 3598
rect 3022 3599 3060 3600
rect 3034 3601 3072 3602
rect 3043 3603 3081 3604
rect 3050 3605 3168 3606
rect 2144 3607 3050 3608
rect 2143 3609 2247 3610
rect 2245 3611 2295 3612
rect 2293 3613 2379 3614
rect 2377 3615 2427 3616
rect 2390 3617 2426 3618
rect 2389 3619 3134 3620
rect 3055 3621 3087 3622
rect 3061 3623 3093 3624
rect 3079 3625 3111 3626
rect 3091 3627 3123 3628
rect 3097 3629 3144 3630
rect 2996 3631 3143 3632
rect 2995 3633 3033 3634
rect 3031 3635 3069 3636
rect 3109 3635 3147 3636
rect 2786 3637 3146 3638
rect 2785 3639 2817 3640
rect 1964 3641 2816 3642
rect 1963 3643 1989 3644
rect 1987 3645 1995 3646
rect 1993 3647 2007 3648
rect 2005 3649 2019 3650
rect 2017 3651 2085 3652
rect 2083 3653 2169 3654
rect 2167 3655 2679 3656
rect 2677 3657 3210 3658
rect 3112 3659 3150 3660
rect 3121 3661 3159 3662
rect 3124 3663 3162 3664
rect 3128 3665 3223 3666
rect 3127 3667 3174 3668
rect 3130 3669 3141 3670
rect 3139 3671 3180 3672
rect 3164 3673 3202 3674
rect 2318 3675 3203 3676
rect 2317 3677 2541 3678
rect 2522 3679 2540 3680
rect 2516 3681 2522 3682
rect 2515 3683 3149 3684
rect 3167 3683 3205 3684
rect 2593 3685 3206 3686
rect 3176 3687 3234 3688
rect 3182 3689 3214 3690
rect 2941 3691 3213 3692
rect 3185 3693 3217 3694
rect 2954 3695 3217 3696
rect 2953 3697 2991 3698
rect 1417 3706 1928 3707
rect 1434 3708 2090 3709
rect 1434 3710 1586 3711
rect 1438 3712 1520 3713
rect 1438 3714 1574 3715
rect 1468 3716 2210 3717
rect 1475 3718 2195 3719
rect 1478 3720 1532 3721
rect 1485 3722 1814 3723
rect 1468 3724 1815 3725
rect 1485 3726 2738 3727
rect 1503 3728 1910 3729
rect 1503 3730 1844 3731
rect 1507 3732 1575 3733
rect 1507 3734 1616 3735
rect 1510 3736 3228 3737
rect 1514 3738 3222 3739
rect 1517 3740 2174 3741
rect 1528 3742 3113 3743
rect 1592 3744 1598 3745
rect 1598 3746 1766 3747
rect 1612 3748 2150 3749
rect 1624 3750 2666 3751
rect 1628 3752 1664 3753
rect 1424 3754 1665 3755
rect 1417 3756 1425 3757
rect 1633 3756 2004 3757
rect 1652 3758 2435 3759
rect 1675 3760 3199 3761
rect 1706 3762 1880 3763
rect 1717 3764 1785 3765
rect 1669 3766 1719 3767
rect 1670 3768 1688 3769
rect 1688 3770 1694 3771
rect 1529 3772 1695 3773
rect 1736 3772 1772 3773
rect 1482 3774 1773 3775
rect 1482 3776 2144 3777
rect 1844 3778 1970 3779
rect 1856 3780 1940 3781
rect 1871 3782 2177 3783
rect 1880 3784 1982 3785
rect 1910 3786 2042 3787
rect 1928 3788 2108 3789
rect 1940 3790 2084 3791
rect 1961 3792 2207 3793
rect 1970 3794 2048 3795
rect 1982 3796 2228 3797
rect 1609 3798 2229 3799
rect 1510 3800 1611 3801
rect 2027 3800 2303 3801
rect 2042 3802 2270 3803
rect 2051 3804 2285 3805
rect 2063 3806 2411 3807
rect 2078 3808 2288 3809
rect 2084 3810 2342 3811
rect 2090 3812 2438 3813
rect 2099 3814 2441 3815
rect 2105 3816 2405 3817
rect 2108 3818 2252 3819
rect 2059 3820 2253 3821
rect 2060 3822 2408 3823
rect 2137 3824 3217 3825
rect 2138 3826 2354 3827
rect 2144 3828 2462 3829
rect 2150 3830 2444 3831
rect 2174 3832 2504 3833
rect 2197 3834 2409 3835
rect 1500 3836 2199 3837
rect 2210 3836 2366 3837
rect 2131 3838 2367 3839
rect 2132 3840 2348 3841
rect 2215 3842 3253 3843
rect 2216 3844 2522 3845
rect 2101 3846 2523 3847
rect 2102 3848 2402 3849
rect 2185 3850 2403 3851
rect 2186 3852 2360 3853
rect 2257 3854 2343 3855
rect 2258 3856 2516 3857
rect 2167 3858 2517 3859
rect 2168 3860 2456 3861
rect 2263 3862 3292 3863
rect 2161 3864 2265 3865
rect 2162 3866 2498 3867
rect 2239 3868 2499 3869
rect 2240 3870 2540 3871
rect 2270 3872 2663 3873
rect 2288 3874 2294 3875
rect 2294 3876 2534 3877
rect 2317 3878 2361 3879
rect 2318 3880 2390 3881
rect 2348 3882 2570 3883
rect 2354 3884 2576 3885
rect 2390 3886 2606 3887
rect 2323 3888 2607 3889
rect 2324 3890 2474 3891
rect 1999 3892 2475 3893
rect 2000 3894 2192 3895
rect 2192 3896 2396 3897
rect 2396 3898 2612 3899
rect 2422 3900 2613 3901
rect 2438 3902 2624 3903
rect 2444 3904 2558 3905
rect 1993 3906 2559 3907
rect 2446 3908 2928 3909
rect 2456 3910 3289 3911
rect 2462 3912 3203 3913
rect 2479 3914 2535 3915
rect 2119 3916 2481 3917
rect 2120 3918 2432 3919
rect 2432 3920 2582 3921
rect 2485 3922 3232 3923
rect 2125 3924 2487 3925
rect 2126 3926 2468 3927
rect 2468 3928 2528 3929
rect 2504 3930 2642 3931
rect 2509 3932 3206 3933
rect 2510 3934 3268 3935
rect 2528 3936 3074 3937
rect 2540 3938 2618 3939
rect 1849 3940 2619 3941
rect 1621 3942 1851 3943
rect 2563 3942 3196 3943
rect 2383 3944 2565 3945
rect 2155 3946 2385 3947
rect 2156 3948 2378 3949
rect 2005 3950 2379 3951
rect 2006 3952 2282 3953
rect 2282 3954 2336 3955
rect 2336 3956 2594 3957
rect 2570 3958 2636 3959
rect 1753 3960 2637 3961
rect 1478 3962 1755 3963
rect 2576 3962 2648 3963
rect 2582 3964 2672 3965
rect 2594 3966 3306 3967
rect 2624 3968 2702 3969
rect 2642 3970 2714 3971
rect 2659 3972 2898 3973
rect 2660 3974 3171 3975
rect 2666 3976 3119 3977
rect 2672 3978 2732 3979
rect 2683 3980 3303 3981
rect 2684 3982 2750 3983
rect 2689 3984 3213 3985
rect 2690 3986 2756 3987
rect 2695 3988 3116 3989
rect 2696 3990 2762 3991
rect 2702 3992 2768 3993
rect 2714 3994 3189 3995
rect 2725 3996 3174 3997
rect 1861 3998 2727 3999
rect 1862 4000 2018 4001
rect 2018 4002 2330 4003
rect 1987 4004 2331 4005
rect 1988 4006 2234 4007
rect 2234 4008 3235 4009
rect 2732 4010 2804 4011
rect 2743 4012 3285 4013
rect 2744 4014 2792 4015
rect 2750 4016 2798 4017
rect 2756 4018 2810 4019
rect 2762 4020 2816 4021
rect 1807 4022 2817 4023
rect 1808 4024 1868 4025
rect 1868 4026 2024 4027
rect 2024 4028 2300 4029
rect 2300 4030 2552 4031
rect 2065 4032 2553 4033
rect 1475 4034 2067 4035
rect 2768 4034 2822 4035
rect 1795 4036 2823 4037
rect 1796 4038 1904 4039
rect 1500 4040 1905 4041
rect 2779 4040 3192 4041
rect 1825 4042 2781 4043
rect 1826 4044 1946 4045
rect 1946 4046 2096 4047
rect 2096 4048 2426 4049
rect 2426 4050 2600 4051
rect 2600 4052 2678 4053
rect 2678 4054 3282 4055
rect 2792 4056 2846 4057
rect 1709 4058 2847 4059
rect 2798 4060 3250 4061
rect 2804 4062 2858 4063
rect 2080 4064 2859 4065
rect 2081 4066 2375 4067
rect 2810 4066 2864 4067
rect 1747 4068 2865 4069
rect 1748 4070 1838 4071
rect 1838 4072 1958 4073
rect 1958 4074 2204 4075
rect 2204 4076 2414 4077
rect 2113 4078 2415 4079
rect 2114 4080 2420 4081
rect 2420 4082 2588 4083
rect 2588 4084 2654 4085
rect 2654 4086 2720 4087
rect 2720 4088 2786 4089
rect 1921 4090 2787 4091
rect 1922 4092 2072 4093
rect 2053 4094 2073 4095
rect 2054 4096 2372 4097
rect 2221 4098 2373 4099
rect 2222 4100 3299 4101
rect 2839 4102 3275 4103
rect 1741 4104 2841 4105
rect 1742 4106 1778 4107
rect 1723 4108 1779 4109
rect 1724 4110 1802 4111
rect 1802 4112 1898 4113
rect 1891 4114 1899 4115
rect 1892 4116 2012 4117
rect 2012 4118 2276 4119
rect 2276 4120 2312 4121
rect 2245 4122 2313 4123
rect 2246 4124 2546 4125
rect 2029 4126 2547 4127
rect 2852 4126 2882 4127
rect 2855 4128 3134 4129
rect 2869 4130 2883 4131
rect 2875 4132 3156 4133
rect 2876 4134 2906 4135
rect 2879 4136 2909 4137
rect 2884 4138 3278 4139
rect 2900 4140 3271 4141
rect 2906 4142 3216 4143
rect 2917 4144 2991 4145
rect 2918 4146 3053 4147
rect 2923 4148 3077 4149
rect 1601 4150 2925 4151
rect 2941 4150 2970 4151
rect 1525 4152 2943 4153
rect 1526 4154 1658 4155
rect 1427 4156 1659 4157
rect 1427 4158 2844 4159
rect 2971 4158 3027 4159
rect 2893 4160 2973 4161
rect 1759 4162 2895 4163
rect 1760 4164 1832 4165
rect 1681 4166 1833 4167
rect 1682 4168 1712 4169
rect 1699 4170 1713 4171
rect 1700 4172 1730 4173
rect 1730 4174 1820 4175
rect 1820 4176 1934 4177
rect 1934 4178 3159 4179
rect 3001 4180 3069 4181
rect 2947 4182 3003 4183
rect 2944 4184 2949 4185
rect 2470 4186 2946 4187
rect 3008 4186 3220 4187
rect 3019 4188 3105 4189
rect 3020 4190 3296 4191
rect 3022 4192 3108 4193
rect 3031 4194 3102 4195
rect 2977 4196 3033 4197
rect 2911 4198 2979 4199
rect 2912 4200 3137 4201
rect 3034 4202 3087 4203
rect 3040 4204 3114 4205
rect 3043 4206 3135 4207
rect 3044 4208 3143 4209
rect 2648 4210 3144 4211
rect 3049 4212 3146 4213
rect 2965 4214 3051 4215
rect 2966 4216 3210 4217
rect 3055 4218 3147 4219
rect 3061 4220 3204 4221
rect 2995 4222 3063 4223
rect 2887 4224 2997 4225
rect 1915 4226 2889 4227
rect 1431 4228 1917 4229
rect 1431 4230 1587 4231
rect 3091 4230 3177 4231
rect 3109 4232 3198 4233
rect 3037 4234 3111 4235
rect 2983 4236 3039 4237
rect 2935 4238 2985 4239
rect 2936 4240 3149 4241
rect 3121 4242 3201 4243
rect 3122 4244 3225 4245
rect 3124 4246 3162 4247
rect 3127 4248 3207 4249
rect 1420 4250 3129 4251
rect 1420 4252 1995 4253
rect 3130 4252 3210 4253
rect 3139 4254 3219 4255
rect 2305 4256 3141 4257
rect 1963 4258 2307 4259
rect 1964 4260 2036 4261
rect 1471 4262 2037 4263
rect 1471 4264 2031 4265
rect 3152 4264 3195 4265
rect 3164 4266 3244 4267
rect 3079 4268 3165 4269
rect 3013 4270 3081 4271
rect 2953 4272 3015 4273
rect 2833 4274 2955 4275
rect 1789 4276 2835 4277
rect 1790 4278 1886 4279
rect 1886 4280 1952 4281
rect 1441 4282 1953 4283
rect 1441 4284 2049 4285
rect 3167 4284 3247 4285
rect 3182 4286 3262 4287
rect 3097 4288 3183 4289
rect 3098 4290 3213 4291
rect 3185 4292 3265 4293
rect 1431 4301 1581 4302
rect 1441 4303 1551 4304
rect 1441 4305 2025 4306
rect 1468 4307 2043 4308
rect 1468 4309 2007 4310
rect 1503 4311 1911 4312
rect 1510 4313 1623 4314
rect 1510 4315 1923 4316
rect 1517 4317 3312 4318
rect 1517 4319 1941 4320
rect 1526 4321 1653 4322
rect 1485 4323 1527 4324
rect 1485 4325 2001 4326
rect 1541 4327 2829 4328
rect 1586 4329 1617 4330
rect 1601 4331 3244 4332
rect 1610 4333 1635 4334
rect 1434 4335 1611 4336
rect 1628 4335 1653 4336
rect 1507 4337 1629 4338
rect 1507 4339 1839 4340
rect 1500 4341 1839 4342
rect 1500 4343 1779 4344
rect 1640 4345 1677 4346
rect 1604 4347 1641 4348
rect 1661 4347 3033 4348
rect 1709 4349 2859 4350
rect 1514 4351 2859 4352
rect 1478 4353 1515 4354
rect 1778 4353 2865 4354
rect 1856 4355 2001 4356
rect 1434 4357 1857 4358
rect 1868 4357 2043 4358
rect 1754 4359 1869 4360
rect 1424 4361 1755 4362
rect 1424 4363 1743 4364
rect 1712 4365 1743 4366
rect 1712 4367 1833 4368
rect 1832 4369 2847 4370
rect 1871 4371 2046 4372
rect 1880 4373 2025 4374
rect 1772 4375 1881 4376
rect 1682 4377 1773 4378
rect 1886 4377 2007 4378
rect 1886 4379 2835 4380
rect 1898 4381 1923 4382
rect 1898 4383 2823 4384
rect 1940 4385 3301 4386
rect 1961 4387 2148 4388
rect 2003 4389 2160 4390
rect 2027 4391 2232 4392
rect 2051 4393 2274 4394
rect 2063 4395 2292 4396
rect 2081 4397 2280 4398
rect 2099 4399 2322 4400
rect 2105 4401 2328 4402
rect 2216 4403 3235 4404
rect 2216 4405 2475 4406
rect 2246 4407 2475 4408
rect 2288 4409 3144 4410
rect 2060 4411 2289 4412
rect 1892 4413 2061 4414
rect 1748 4415 1893 4416
rect 1748 4417 1785 4418
rect 1784 4419 2613 4420
rect 2357 4421 2898 4422
rect 2402 4423 3371 4424
rect 2192 4425 2403 4426
rect 2108 4427 2193 4428
rect 2429 4427 2844 4428
rect 2438 4429 2613 4430
rect 2438 4431 2547 4432
rect 2354 4433 2547 4434
rect 2186 4435 2355 4436
rect 2186 4437 2559 4438
rect 2384 4439 2559 4440
rect 2162 4441 2385 4442
rect 2162 4443 2253 4444
rect 2252 4445 2271 4446
rect 2048 4447 2271 4448
rect 2048 4449 2307 4450
rect 2138 4451 2307 4452
rect 1976 4453 2139 4454
rect 1478 4455 1977 4456
rect 2450 4455 3396 4456
rect 2222 4457 2451 4458
rect 2018 4459 2223 4460
rect 1874 4461 2019 4462
rect 1760 4463 1875 4464
rect 1503 4465 1761 4466
rect 2504 4465 3368 4466
rect 2294 4467 2505 4468
rect 1427 4469 2295 4470
rect 1427 4471 2109 4472
rect 2594 4471 2739 4472
rect 2426 4473 2595 4474
rect 2210 4475 2427 4476
rect 2078 4477 2211 4478
rect 1904 4479 2079 4480
rect 1808 4481 1905 4482
rect 1420 4483 1809 4484
rect 1420 4485 2247 4486
rect 2684 4485 3282 4486
rect 2534 4487 2685 4488
rect 2414 4489 2535 4490
rect 2414 4491 3327 4492
rect 2690 4493 2829 4494
rect 2540 4495 2691 4496
rect 2348 4497 2541 4498
rect 2126 4499 2349 4500
rect 1970 4501 2127 4502
rect 1820 4503 1971 4504
rect 1820 4505 2925 4506
rect 2696 4507 2835 4508
rect 2696 4509 2727 4510
rect 2582 4511 2727 4512
rect 2390 4513 2583 4514
rect 1417 4515 2391 4516
rect 1417 4517 1483 4518
rect 1482 4519 1995 4520
rect 1850 4521 1995 4522
rect 1475 4523 1851 4524
rect 2708 4523 3024 4524
rect 2570 4525 2709 4526
rect 2408 4527 2571 4528
rect 2198 4529 2409 4530
rect 2030 4531 2199 4532
rect 2030 4533 2457 4534
rect 2456 4535 3399 4536
rect 2714 4537 3334 4538
rect 2576 4539 2715 4540
rect 2480 4541 2577 4542
rect 2282 4543 2481 4544
rect 1438 4545 2283 4546
rect 2786 4545 2925 4546
rect 2648 4547 2787 4548
rect 2516 4549 2649 4550
rect 2324 4551 2517 4552
rect 2102 4553 2325 4554
rect 1964 4555 2103 4556
rect 1538 4557 1965 4558
rect 2792 4557 2931 4558
rect 2654 4559 2793 4560
rect 2492 4561 2655 4562
rect 2342 4563 2493 4564
rect 2120 4565 2343 4566
rect 1946 4567 2121 4568
rect 1946 4569 3253 4570
rect 2822 4571 3285 4572
rect 2840 4573 3375 4574
rect 2702 4575 2841 4576
rect 2564 4577 2703 4578
rect 2522 4579 2565 4580
rect 2372 4581 2523 4582
rect 2180 4583 2373 4584
rect 2180 4585 2265 4586
rect 2084 4587 2265 4588
rect 1928 4589 2085 4590
rect 1814 4591 1929 4592
rect 1814 4593 2637 4594
rect 2486 4595 2637 4596
rect 2360 4597 2487 4598
rect 2150 4599 2361 4600
rect 2150 4601 2229 4602
rect 1438 4603 2229 4604
rect 2855 4603 2871 4604
rect 2864 4605 3324 4606
rect 2876 4607 3271 4608
rect 2744 4609 2877 4610
rect 2600 4611 2745 4612
rect 2420 4613 2601 4614
rect 2204 4615 2421 4616
rect 1471 4617 2205 4618
rect 1471 4619 2013 4620
rect 1844 4621 2013 4622
rect 1724 4623 1845 4624
rect 1664 4625 1725 4626
rect 1529 4627 1665 4628
rect 1529 4629 1605 4630
rect 2906 4629 3159 4630
rect 2906 4631 3292 4632
rect 2918 4633 3216 4634
rect 2816 4635 2919 4636
rect 2678 4637 2817 4638
rect 2552 4639 2679 4640
rect 2336 4641 2553 4642
rect 2114 4643 2337 4644
rect 1952 4645 2115 4646
rect 1796 4647 1953 4648
rect 1796 4649 2895 4650
rect 2762 4651 2895 4652
rect 2624 4653 2763 4654
rect 2462 4655 2625 4656
rect 2240 4657 2463 4658
rect 2036 4659 2241 4660
rect 1862 4661 2037 4662
rect 1730 4663 1863 4664
rect 1670 4665 1731 4666
rect 2921 4665 2928 4666
rect 2945 4665 3000 4666
rect 2966 4667 3093 4668
rect 2966 4669 3238 4670
rect 2969 4671 3096 4672
rect 3002 4673 3117 4674
rect 2852 4675 3003 4676
rect 2720 4677 2853 4678
rect 2588 4679 2721 4680
rect 2396 4681 2589 4682
rect 2174 4683 2397 4684
rect 1988 4685 2175 4686
rect 1431 4687 1989 4688
rect 3005 4687 3289 4688
rect 3014 4689 3033 4690
rect 3014 4691 3213 4692
rect 3038 4693 3296 4694
rect 2972 4695 3039 4696
rect 1706 4697 2973 4698
rect 1706 4699 1719 4700
rect 1658 4701 1719 4702
rect 1658 4703 3306 4704
rect 2996 4705 3305 4706
rect 2942 4707 2997 4708
rect 2942 4709 3275 4710
rect 3056 4711 3378 4712
rect 3062 4713 3159 4714
rect 2936 4715 3063 4716
rect 2798 4717 2937 4718
rect 2660 4719 2799 4720
rect 2498 4721 2661 4722
rect 2318 4723 2499 4724
rect 2090 4725 2319 4726
rect 2090 4727 3299 4728
rect 3068 4729 3153 4730
rect 2948 4731 3069 4732
rect 2804 4733 2949 4734
rect 2672 4735 2805 4736
rect 2528 4737 2673 4738
rect 2366 4739 2529 4740
rect 2144 4741 2367 4742
rect 1958 4743 2145 4744
rect 1802 4745 1959 4746
rect 1802 4747 2901 4748
rect 2768 4749 2901 4750
rect 2630 4751 2769 4752
rect 2468 4753 2631 4754
rect 2234 4755 2469 4756
rect 2234 4757 2313 4758
rect 2096 4759 2313 4760
rect 1934 4761 2097 4762
rect 1790 4763 1935 4764
rect 1700 4765 1791 4766
rect 1598 4767 1701 4768
rect 1568 4769 1599 4770
rect 3074 4769 3278 4770
rect 3080 4771 3250 4772
rect 2990 4773 3081 4774
rect 2990 4775 3385 4776
rect 3098 4777 3189 4778
rect 2978 4779 3099 4780
rect 2888 4781 2979 4782
rect 2756 4783 2889 4784
rect 2666 4785 2757 4786
rect 2510 4787 2667 4788
rect 2300 4789 2511 4790
rect 2132 4791 2301 4792
rect 2072 4793 2133 4794
rect 1916 4795 2073 4796
rect 1916 4797 2619 4798
rect 2444 4799 2619 4800
rect 2258 4801 2445 4802
rect 2066 4803 2259 4804
rect 2066 4805 2379 4806
rect 2168 4807 2379 4808
rect 1982 4809 2169 4810
rect 1826 4811 1983 4812
rect 1736 4813 1827 4814
rect 1688 4815 1737 4816
rect 1688 4817 1695 4818
rect 3101 4817 3192 4818
rect 3104 4819 3216 4820
rect 2984 4821 3105 4822
rect 3128 4821 3225 4822
rect 3050 4823 3129 4824
rect 2912 4825 3051 4826
rect 2774 4827 2913 4828
rect 2774 4829 3303 4830
rect 3134 4831 3228 4832
rect 3026 4833 3135 4834
rect 2882 4835 3027 4836
rect 2750 4837 2883 4838
rect 2750 4839 2781 4840
rect 2642 4841 2781 4842
rect 2642 4843 3361 4844
rect 3140 4845 3162 4846
rect 3164 4845 3244 4846
rect 3107 4847 3165 4848
rect 3176 4847 3321 4848
rect 3086 4849 3177 4850
rect 3194 4849 3274 4850
rect 3110 4851 3195 4852
rect 3008 4853 3111 4854
rect 2954 4855 3009 4856
rect 2810 4857 2955 4858
rect 2732 4859 2811 4860
rect 2606 4861 2733 4862
rect 2432 4863 2607 4864
rect 2276 4865 2433 4866
rect 2054 4867 2277 4868
rect 2054 4869 2331 4870
rect 2156 4871 2331 4872
rect 2156 4873 3232 4874
rect 3170 4875 3231 4876
rect 3197 4877 3277 4878
rect 3113 4879 3198 4880
rect 3200 4879 3295 4880
rect 3200 4881 3222 4882
rect 3203 4883 3225 4884
rect 3044 4885 3204 4886
rect 1475 4887 3045 4888
rect 3206 4887 3286 4888
rect 3122 4889 3207 4890
rect 3020 4891 3123 4892
rect 2879 4893 3021 4894
rect 3209 4893 3289 4894
rect 3212 4895 3308 4896
rect 3218 4897 3234 4898
rect 3146 4899 3219 4900
rect 3240 4899 3315 4900
rect 3246 4901 3318 4902
rect 3261 4903 3355 4904
rect 3182 4905 3262 4906
rect 3264 4905 3358 4906
rect 3267 4907 3298 4908
rect 3291 4909 3364 4910
rect 3330 4911 3382 4912
rect 3336 4913 3389 4914
rect 3342 4915 3392 4916
rect 1434 4924 1953 4925
rect 1438 4926 2139 4927
rect 1447 4928 2061 4929
rect 1471 4930 2007 4931
rect 1478 4932 1971 4933
rect 1477 4934 1989 4935
rect 1482 4936 2157 4937
rect 1488 4938 2328 4939
rect 1491 4940 2283 4941
rect 1503 4942 1749 4943
rect 1514 4944 2313 4945
rect 1510 4946 2313 4947
rect 1517 4948 2880 4949
rect 1519 4950 2193 4951
rect 1526 4952 1905 4953
rect 1526 4954 2505 4955
rect 1529 4956 3015 4957
rect 1538 4958 1887 4959
rect 1541 4960 1839 4961
rect 1468 4962 1839 4963
rect 1462 4964 1469 4965
rect 1456 4966 1463 4967
rect 1450 4968 1457 4969
rect 1556 4968 2826 4969
rect 1574 4970 1587 4971
rect 1580 4972 2148 4973
rect 1634 4974 1647 4975
rect 1622 4976 1635 4977
rect 1610 4978 1623 4979
rect 1598 4980 1611 4981
rect 1562 4982 1599 4983
rect 1550 4984 1563 4985
rect 1652 4984 1671 4985
rect 1640 4986 1653 4987
rect 1628 4988 1641 4989
rect 1616 4990 1629 4991
rect 1694 4990 1719 4991
rect 1742 4990 1767 4991
rect 1742 4992 1791 4993
rect 1748 4994 1755 4995
rect 1688 4996 1755 4997
rect 1481 4998 1689 4999
rect 1790 4998 1845 4999
rect 1829 5000 2046 5001
rect 1844 5002 2073 5003
rect 1904 5004 2289 5005
rect 1661 5006 2289 5007
rect 1907 5008 2292 5009
rect 1910 5010 2229 5011
rect 1937 5012 2232 5013
rect 1952 5014 2241 5015
rect 1970 5016 2349 5017
rect 1976 5018 2193 5019
rect 1976 5020 2343 5021
rect 1982 5022 2157 5023
rect 1982 5024 2205 5025
rect 1988 5026 2367 5027
rect 2006 5028 2361 5029
rect 2060 5030 2265 5031
rect 2069 5032 2274 5033
rect 2072 5034 2301 5035
rect 2102 5036 2349 5037
rect 2102 5038 2403 5039
rect 2132 5040 2361 5041
rect 2132 5042 2409 5043
rect 2126 5044 2409 5045
rect 2126 5046 2463 5047
rect 2138 5048 2421 5049
rect 2150 5050 2229 5051
rect 2150 5052 2427 5053
rect 2159 5054 2574 5055
rect 2180 5056 2301 5057
rect 2090 5058 2181 5059
rect 2090 5060 2451 5061
rect 2204 5062 2511 5063
rect 2234 5064 2241 5065
rect 2234 5066 3327 5067
rect 2264 5068 2541 5069
rect 2282 5070 2295 5071
rect 2294 5072 2493 5073
rect 1868 5074 2493 5075
rect 2342 5076 2595 5077
rect 1760 5078 2595 5079
rect 1760 5080 1863 5081
rect 1862 5082 2145 5083
rect 2144 5084 2475 5085
rect 1874 5086 2475 5087
rect 1658 5088 1875 5089
rect 1604 5090 1659 5091
rect 1592 5092 1605 5093
rect 1433 5094 1593 5095
rect 2357 5094 3036 5095
rect 2279 5096 2358 5097
rect 2366 5096 2601 5097
rect 2216 5098 2601 5099
rect 2216 5100 2481 5101
rect 1856 5102 2481 5103
rect 1856 5104 2109 5105
rect 2108 5106 2355 5107
rect 1475 5108 2355 5109
rect 1474 5110 2115 5111
rect 2114 5112 3452 5113
rect 2402 5114 3469 5115
rect 2420 5116 2631 5117
rect 2426 5118 2625 5119
rect 2444 5120 3305 5121
rect 2444 5122 2529 5123
rect 1994 5124 2529 5125
rect 1994 5126 2175 5127
rect 1889 5128 2175 5129
rect 2450 5128 2655 5129
rect 2462 5130 2643 5131
rect 2468 5132 3455 5133
rect 2024 5134 2469 5135
rect 2024 5136 2211 5137
rect 2210 5138 2433 5139
rect 2432 5140 2571 5141
rect 1880 5142 2571 5143
rect 1880 5144 2085 5145
rect 2084 5146 2307 5147
rect 1507 5148 2307 5149
rect 2504 5148 2661 5149
rect 2186 5150 2661 5151
rect 2120 5152 2187 5153
rect 2120 5154 3324 5155
rect 2510 5156 2667 5157
rect 1541 5158 2667 5159
rect 2540 5160 3334 5161
rect 2552 5162 3382 5163
rect 2552 5164 2685 5165
rect 2576 5166 3459 5167
rect 2576 5168 2673 5169
rect 1940 5170 2673 5171
rect 1940 5172 2319 5173
rect 2318 5174 2583 5175
rect 2048 5176 2583 5177
rect 2048 5178 2415 5179
rect 2414 5180 3368 5181
rect 2618 5182 3371 5183
rect 2030 5184 2619 5185
rect 2030 5186 2379 5187
rect 2378 5188 2607 5189
rect 2606 5190 2709 5191
rect 2624 5192 2739 5193
rect 2630 5194 2715 5195
rect 2642 5196 2679 5197
rect 2654 5198 2733 5199
rect 1850 5200 2733 5201
rect 1424 5202 1851 5203
rect 1423 5204 1557 5205
rect 2678 5204 2781 5205
rect 1512 5206 2781 5207
rect 2684 5208 3308 5209
rect 2708 5210 2799 5211
rect 2714 5212 2793 5213
rect 2738 5214 2829 5215
rect 2744 5216 3408 5217
rect 2744 5218 2835 5219
rect 2762 5220 3430 5221
rect 2762 5222 2853 5223
rect 2768 5224 3364 5225
rect 2756 5226 2769 5227
rect 2792 5226 2865 5227
rect 2798 5228 2877 5229
rect 1500 5230 2877 5231
rect 1494 5232 1501 5233
rect 2816 5232 3462 5233
rect 1946 5234 2817 5235
rect 1946 5236 2325 5237
rect 2324 5238 2589 5239
rect 2054 5240 2589 5241
rect 2054 5242 3466 5243
rect 2828 5244 2901 5245
rect 2834 5246 2907 5247
rect 2846 5248 2889 5249
rect 2750 5250 2889 5251
rect 2750 5252 2841 5253
rect 1916 5254 2841 5255
rect 1916 5256 2271 5257
rect 2270 5258 2517 5259
rect 2000 5260 2517 5261
rect 2000 5262 2385 5263
rect 1427 5264 2385 5265
rect 1426 5266 1878 5267
rect 2852 5266 2895 5267
rect 2858 5268 3401 5269
rect 2858 5270 2931 5271
rect 1898 5272 2931 5273
rect 1898 5274 2223 5275
rect 2222 5276 2253 5277
rect 2252 5278 3328 5279
rect 2864 5280 2937 5281
rect 2870 5282 3445 5283
rect 2870 5284 2913 5285
rect 2894 5286 2949 5287
rect 1706 5288 2949 5289
rect 1706 5290 1731 5291
rect 1730 5292 2322 5293
rect 2900 5292 2955 5293
rect 1832 5294 2955 5295
rect 1431 5296 1833 5297
rect 1430 5298 1539 5299
rect 2912 5298 2967 5299
rect 2921 5300 3108 5301
rect 2924 5302 3241 5303
rect 2918 5304 2925 5305
rect 2918 5306 3238 5307
rect 2942 5308 3385 5309
rect 1964 5310 2943 5311
rect 1964 5312 2199 5313
rect 2078 5314 2199 5315
rect 2078 5316 2331 5317
rect 2096 5318 2331 5319
rect 2096 5320 2457 5321
rect 2456 5322 2559 5323
rect 2558 5324 2637 5325
rect 2636 5326 2703 5327
rect 2702 5328 2775 5329
rect 2774 5330 2805 5331
rect 2804 5332 2883 5333
rect 2696 5334 2883 5335
rect 2696 5336 3324 5337
rect 2960 5338 3003 5339
rect 1712 5340 3003 5341
rect 1712 5342 1737 5343
rect 1664 5344 1737 5345
rect 2963 5344 3006 5345
rect 2966 5346 2973 5347
rect 1808 5348 2973 5349
rect 1808 5350 1959 5351
rect 1958 5352 2337 5353
rect 2336 5354 2523 5355
rect 2066 5356 2523 5357
rect 2066 5358 2169 5359
rect 2168 5360 2247 5361
rect 2246 5362 2499 5363
rect 1928 5364 2499 5365
rect 1928 5366 2259 5367
rect 2258 5368 2547 5369
rect 2546 5370 2691 5371
rect 2690 5372 2787 5373
rect 2786 5374 3448 5375
rect 2981 5376 3024 5377
rect 2429 5378 3024 5379
rect 2984 5380 3027 5381
rect 1778 5382 3027 5383
rect 1444 5384 1779 5385
rect 2999 5384 3222 5385
rect 3014 5386 3057 5387
rect 3032 5388 3147 5389
rect 1796 5390 3033 5391
rect 1796 5392 1827 5393
rect 1826 5394 2043 5395
rect 2042 5396 2373 5397
rect 2372 5398 2613 5399
rect 2612 5400 2727 5401
rect 2726 5402 2823 5403
rect 1515 5404 2823 5405
rect 3050 5404 3375 5405
rect 1820 5406 3051 5407
rect 1820 5408 2037 5409
rect 2036 5410 2391 5411
rect 2162 5412 2391 5413
rect 1485 5414 2163 5415
rect 1484 5416 1677 5417
rect 1676 5418 3423 5419
rect 3056 5420 3069 5421
rect 3068 5422 3298 5423
rect 3098 5424 3141 5425
rect 3116 5426 3420 5427
rect 3104 5428 3117 5429
rect 1700 5430 3105 5431
rect 1700 5432 1725 5433
rect 1724 5434 1773 5435
rect 1417 5436 1773 5437
rect 3170 5436 3279 5437
rect 3170 5438 3312 5439
rect 3182 5440 3315 5441
rect 3188 5442 3249 5443
rect 3128 5444 3189 5445
rect 3038 5446 3129 5447
rect 1437 5448 3039 5449
rect 3203 5448 3264 5449
rect 3206 5450 3267 5451
rect 3158 5452 3207 5453
rect 3134 5454 3159 5455
rect 3044 5456 3135 5457
rect 1802 5458 3045 5459
rect 1802 5460 1935 5461
rect 1441 5462 1935 5463
rect 1440 5464 2013 5465
rect 2012 5466 2397 5467
rect 2396 5468 3427 5469
rect 3212 5470 3309 5471
rect 3164 5472 3213 5473
rect 3122 5474 3165 5475
rect 3080 5476 3123 5477
rect 3074 5478 3081 5479
rect 3062 5480 3075 5481
rect 1522 5482 3063 5483
rect 3215 5482 3312 5483
rect 3218 5484 3315 5485
rect 2996 5486 3219 5487
rect 1814 5488 2997 5489
rect 1529 5490 1815 5491
rect 3224 5490 3297 5491
rect 3176 5492 3225 5493
rect 3236 5492 3378 5493
rect 3243 5494 3334 5495
rect 3251 5496 3396 5497
rect 2990 5498 3397 5499
rect 2990 5500 3394 5501
rect 3273 5502 3370 5503
rect 3272 5504 3301 5505
rect 3276 5506 3373 5507
rect 3194 5508 3276 5509
rect 3194 5510 3198 5511
rect 3285 5510 3382 5511
rect 3230 5512 3285 5513
rect 3191 5514 3231 5515
rect 3288 5514 3385 5515
rect 3317 5516 3414 5517
rect 3320 5518 3340 5519
rect 2720 5520 3321 5521
rect 1922 5522 2721 5523
rect 1922 5524 2277 5525
rect 2276 5526 2487 5527
rect 2486 5528 2535 5529
rect 2534 5530 2649 5531
rect 2438 5532 2649 5533
rect 2018 5534 2439 5535
rect 1886 5536 2019 5537
rect 3330 5536 3399 5537
rect 2936 5538 3331 5539
rect 3336 5538 3442 5539
rect 3342 5540 3439 5541
rect 3354 5542 3392 5543
rect 3294 5544 3391 5545
rect 3357 5546 3389 5547
rect 3261 5548 3358 5549
rect 3200 5550 3261 5551
rect 3152 5552 3201 5553
rect 3110 5554 3153 5555
rect 3008 5556 3111 5557
rect 2978 5558 3009 5559
rect 2978 5560 3021 5561
rect 1784 5562 3021 5563
rect 1784 5564 1893 5565
rect 1420 5566 1893 5567
rect 3291 5566 3388 5567
rect 3233 5568 3291 5569
rect 3360 5568 3417 5569
rect 3403 5570 3411 5571
rect 1420 5579 1833 5580
rect 1423 5581 1920 5582
rect 1433 5583 1908 5584
rect 1434 5585 1695 5586
rect 1437 5587 1968 5588
rect 1438 5589 2781 5590
rect 1440 5591 2595 5592
rect 1441 5593 1593 5594
rect 1444 5595 1653 5596
rect 1445 5597 1581 5598
rect 1481 5599 2574 5600
rect 1482 5601 2181 5602
rect 1477 5603 2181 5604
rect 1484 5605 2568 5606
rect 1488 5607 2247 5608
rect 1515 5609 2997 5610
rect 1519 5611 1557 5612
rect 1522 5613 3021 5614
rect 1532 5615 1659 5616
rect 1535 5617 1653 5618
rect 1541 5619 2673 5620
rect 1544 5621 1551 5622
rect 1544 5623 2769 5624
rect 1547 5625 2235 5626
rect 1556 5627 1563 5628
rect 1568 5627 1878 5628
rect 1580 5629 1587 5630
rect 1592 5629 1605 5630
rect 1604 5631 1890 5632
rect 1426 5633 1890 5634
rect 1427 5635 1875 5636
rect 1616 5637 1623 5638
rect 1622 5639 1629 5640
rect 1598 5641 1629 5642
rect 1598 5643 1611 5644
rect 1430 5645 1611 5646
rect 1664 5645 1677 5646
rect 1676 5647 1689 5648
rect 1682 5649 1701 5650
rect 1688 5651 1707 5652
rect 1694 5653 1713 5654
rect 1700 5655 1731 5656
rect 1712 5657 1725 5658
rect 1526 5659 1725 5660
rect 1525 5661 2073 5662
rect 1718 5663 1767 5664
rect 1730 5665 1743 5666
rect 1742 5667 1749 5668
rect 1670 5669 1749 5670
rect 1754 5669 3397 5670
rect 1754 5671 2877 5672
rect 1766 5673 1797 5674
rect 1736 5675 1797 5676
rect 1431 5677 1737 5678
rect 1808 5677 1833 5678
rect 1485 5679 1809 5680
rect 1868 5679 2070 5680
rect 1874 5681 1881 5682
rect 1880 5683 2067 5684
rect 1886 5685 2958 5686
rect 1424 5687 1887 5688
rect 1925 5687 1938 5688
rect 1988 5687 3462 5688
rect 1940 5689 1989 5690
rect 1928 5691 1941 5692
rect 1928 5693 1995 5694
rect 1946 5695 1995 5696
rect 1922 5697 1947 5698
rect 1910 5699 1923 5700
rect 1898 5701 1911 5702
rect 1417 5703 1899 5704
rect 2033 5703 2241 5704
rect 2042 5705 2073 5706
rect 2030 5707 2043 5708
rect 2120 5707 3455 5708
rect 2090 5709 2121 5710
rect 2054 5711 2091 5712
rect 2036 5713 2055 5714
rect 2036 5715 2061 5716
rect 2012 5717 2061 5718
rect 2012 5719 2019 5720
rect 1970 5721 2019 5722
rect 1489 5723 1971 5724
rect 2234 5723 2283 5724
rect 2228 5725 2283 5726
rect 2186 5727 2229 5728
rect 2240 5727 2253 5728
rect 2246 5729 2271 5730
rect 2252 5731 2259 5732
rect 2258 5733 2265 5734
rect 2264 5735 3362 5736
rect 2270 5737 2295 5738
rect 2276 5739 3328 5740
rect 2276 5741 2289 5742
rect 2198 5743 2289 5744
rect 2198 5745 2211 5746
rect 2210 5747 2217 5748
rect 2156 5749 2217 5750
rect 2144 5751 2157 5752
rect 2114 5753 2145 5754
rect 2084 5755 2115 5756
rect 1474 5757 2085 5758
rect 1475 5759 2187 5760
rect 2294 5759 2307 5760
rect 2300 5761 3466 5762
rect 2300 5763 2313 5764
rect 2306 5765 2319 5766
rect 2312 5767 2325 5768
rect 2318 5769 2331 5770
rect 2324 5771 2349 5772
rect 2330 5773 2355 5774
rect 2333 5775 2358 5776
rect 2336 5777 3355 5778
rect 2336 5779 2367 5780
rect 2348 5781 2379 5782
rect 2354 5783 2361 5784
rect 2360 5785 2385 5786
rect 2366 5787 2397 5788
rect 2378 5789 2403 5790
rect 2384 5791 3331 5792
rect 2396 5793 2415 5794
rect 2402 5795 2427 5796
rect 2408 5797 2415 5798
rect 2408 5799 3406 5800
rect 2420 5801 3452 5802
rect 2222 5803 3452 5804
rect 2192 5805 2223 5806
rect 1478 5807 2193 5808
rect 2420 5807 2439 5808
rect 2426 5809 2451 5810
rect 2438 5811 2457 5812
rect 2450 5813 2469 5814
rect 2456 5815 2475 5816
rect 2468 5817 3324 5818
rect 2474 5819 2493 5820
rect 2486 5821 3321 5822
rect 2486 5823 3396 5824
rect 2492 5825 2505 5826
rect 2504 5827 2517 5828
rect 2516 5829 2529 5830
rect 2528 5831 2541 5832
rect 2540 5833 2553 5834
rect 2591 5833 2880 5834
rect 2594 5835 2619 5836
rect 2606 5837 2619 5838
rect 2606 5839 2649 5840
rect 2648 5841 2667 5842
rect 2672 5841 2679 5842
rect 2678 5843 2685 5844
rect 2684 5845 2691 5846
rect 2690 5847 2703 5848
rect 2696 5849 3366 5850
rect 2696 5851 2709 5852
rect 2702 5853 2715 5854
rect 2708 5855 2721 5856
rect 2714 5857 3469 5858
rect 2720 5859 2727 5860
rect 2726 5861 3408 5862
rect 2756 5863 2763 5864
rect 2762 5865 2775 5866
rect 2768 5867 2823 5868
rect 2774 5869 3404 5870
rect 2780 5871 3448 5872
rect 2432 5873 3449 5874
rect 2432 5875 2445 5876
rect 2444 5877 2463 5878
rect 2462 5879 2481 5880
rect 2480 5881 2499 5882
rect 2498 5883 2511 5884
rect 2510 5885 2523 5886
rect 2522 5887 2535 5888
rect 2534 5889 2547 5890
rect 2546 5891 2559 5892
rect 2558 5893 2565 5894
rect 2564 5895 2571 5896
rect 2570 5897 2577 5898
rect 1516 5899 2577 5900
rect 2786 5899 3430 5900
rect 2786 5901 2799 5902
rect 2792 5903 3445 5904
rect 2792 5905 2805 5906
rect 1512 5907 2805 5908
rect 1513 5909 1905 5910
rect 1904 5911 1935 5912
rect 1916 5913 1935 5914
rect 1892 5915 1917 5916
rect 1491 5917 1893 5918
rect 1492 5919 2601 5920
rect 2600 5921 2613 5922
rect 2612 5923 2625 5924
rect 2624 5925 2661 5926
rect 1538 5927 2661 5928
rect 2798 5927 2817 5928
rect 2801 5929 3024 5930
rect 2807 5931 2826 5932
rect 2810 5933 3401 5934
rect 2810 5935 2829 5936
rect 2816 5937 2835 5938
rect 2822 5939 2841 5940
rect 2828 5941 2847 5942
rect 2834 5943 2853 5944
rect 2840 5945 2859 5946
rect 2846 5947 2865 5948
rect 2852 5949 2871 5950
rect 2858 5951 3027 5952
rect 2864 5953 2883 5954
rect 2870 5955 2889 5956
rect 2876 5957 2895 5958
rect 2882 5959 2901 5960
rect 2888 5961 2964 5962
rect 2900 5963 2913 5964
rect 2906 5965 3352 5966
rect 2912 5967 2919 5968
rect 2918 5969 2925 5970
rect 2924 5971 2931 5972
rect 2930 5973 2937 5974
rect 2936 5975 2943 5976
rect 2942 5977 2973 5978
rect 2948 5979 3445 5980
rect 2948 5981 2955 5982
rect 2954 5983 2961 5984
rect 2960 5985 2967 5986
rect 2966 5987 3033 5988
rect 2972 5989 2979 5990
rect 2975 5991 2982 5992
rect 2978 5993 2985 5994
rect 2984 5995 2991 5996
rect 2990 5997 3394 5998
rect 2996 5999 3045 6000
rect 3011 6001 3036 6002
rect 3020 6003 3063 6004
rect 3026 6005 3069 6006
rect 3044 6007 3075 6008
rect 3062 6009 3111 6010
rect 3068 6011 3096 6012
rect 3074 6013 3093 6014
rect 3086 6015 3129 6016
rect 3092 6017 3117 6018
rect 3098 6019 3135 6020
rect 3104 6021 3111 6022
rect 3104 6023 3141 6024
rect 3107 6025 3114 6026
rect 3134 6025 3183 6026
rect 3140 6027 3189 6028
rect 3152 6029 3423 6030
rect 2126 6031 3424 6032
rect 2096 6033 2127 6034
rect 2096 6035 2151 6036
rect 2138 6037 2151 6038
rect 2138 6039 2163 6040
rect 2162 6041 2169 6042
rect 2168 6043 2175 6044
rect 1447 6045 2175 6046
rect 1448 6047 2553 6048
rect 3146 6047 3153 6048
rect 3146 6049 3195 6050
rect 3158 6051 3403 6052
rect 3158 6053 3207 6054
rect 3164 6055 3283 6056
rect 3164 6057 3201 6058
rect 3176 6059 3225 6060
rect 3182 6061 3231 6062
rect 3188 6063 3431 6064
rect 3200 6065 3249 6066
rect 3203 6067 3252 6068
rect 3206 6069 3219 6070
rect 3209 6071 3222 6072
rect 3218 6073 3261 6074
rect 3221 6075 3264 6076
rect 3224 6077 3267 6078
rect 3230 6079 3273 6080
rect 2588 6081 3273 6082
rect 2588 6083 2733 6084
rect 2732 6085 2739 6086
rect 2738 6087 2745 6088
rect 2744 6089 2751 6090
rect 3233 6089 3276 6090
rect 1640 6091 3276 6092
rect 1634 6093 1641 6094
rect 3242 6093 3285 6094
rect 3248 6095 3291 6096
rect 3260 6097 3309 6098
rect 3263 6099 3312 6100
rect 3266 6101 3315 6102
rect 3285 6103 3334 6104
rect 3291 6105 3340 6106
rect 2030 6107 3340 6108
rect 3296 6109 3399 6110
rect 3309 6111 3358 6112
rect 2066 6113 3359 6114
rect 3315 6115 3385 6116
rect 3321 6117 3370 6118
rect 2666 6119 3369 6120
rect 3324 6121 3373 6122
rect 3342 6123 3382 6124
rect 3345 6125 3388 6126
rect 3348 6127 3391 6128
rect 3371 6129 3414 6130
rect 3374 6131 3417 6132
rect 3377 6133 3435 6134
rect 3389 6135 3420 6136
rect 2342 6137 3421 6138
rect 2342 6139 2373 6140
rect 2372 6141 3427 6142
rect 3236 6143 3428 6144
rect 3236 6145 3279 6146
rect 3116 6147 3280 6148
rect 3410 6147 3459 6148
rect 3414 6149 3439 6150
rect 3392 6151 3438 6152
rect 3417 6153 3442 6154
rect 3014 6155 3442 6156
rect 3014 6157 3039 6158
rect 3038 6159 3051 6160
rect 3050 6161 3057 6162
rect 3056 6163 3081 6164
rect 3080 6165 3123 6166
rect 3122 6167 3171 6168
rect 3170 6169 3213 6170
rect 1417 6178 1851 6179
rect 1417 6180 1514 6181
rect 1420 6182 2187 6183
rect 1420 6184 1669 6185
rect 1424 6186 1813 6187
rect 1424 6188 1605 6189
rect 1427 6190 1483 6191
rect 1427 6192 1599 6193
rect 1431 6194 1675 6195
rect 1431 6196 1693 6197
rect 1434 6198 1731 6199
rect 1434 6200 1442 6201
rect 1438 6202 2167 6203
rect 1438 6204 1687 6205
rect 1441 6206 1743 6207
rect 1448 6208 2289 6209
rect 1448 6210 2845 6211
rect 1457 6212 1476 6213
rect 1457 6214 1464 6215
rect 1463 6216 1470 6217
rect 1469 6218 2808 6219
rect 1472 6220 2637 6221
rect 1476 6222 1747 6223
rect 1478 6224 2439 6225
rect 1479 6226 1629 6227
rect 1485 6228 2523 6229
rect 1489 6230 2547 6231
rect 1492 6232 1767 6233
rect 1494 6234 1502 6235
rect 1500 6236 1645 6237
rect 1503 6238 1701 6239
rect 1512 6240 1548 6241
rect 1516 6242 1890 6243
rect 1515 6244 2181 6245
rect 1518 6246 1551 6247
rect 1525 6248 1677 6249
rect 1524 6250 1557 6251
rect 1528 6252 2097 6253
rect 1532 6254 3012 6255
rect 1539 6256 1771 6257
rect 1542 6258 1581 6259
rect 1554 6260 1593 6261
rect 1560 6262 1611 6263
rect 1566 6264 1617 6265
rect 1572 6266 1623 6267
rect 1584 6268 2727 6269
rect 1587 6270 2805 6271
rect 1596 6272 1647 6273
rect 1608 6274 2649 6275
rect 1611 6276 2341 6277
rect 1614 6278 1665 6279
rect 1620 6280 1683 6281
rect 1626 6282 1689 6283
rect 1632 6284 1695 6285
rect 1652 6286 2034 6287
rect 1656 6288 1713 6289
rect 1662 6290 1725 6291
rect 1680 6292 1737 6293
rect 1698 6294 1719 6295
rect 1710 6296 1755 6297
rect 1716 6298 1797 6299
rect 1722 6300 1791 6301
rect 1728 6302 2565 6303
rect 1734 6304 1761 6305
rect 1740 6306 2475 6307
rect 1752 6308 2457 6309
rect 1758 6310 1773 6311
rect 1764 6312 1779 6313
rect 1776 6314 2361 6315
rect 1782 6316 1785 6317
rect 1788 6316 2463 6317
rect 1794 6318 2589 6319
rect 1800 6320 1869 6321
rect 1802 6322 1837 6323
rect 1806 6324 1809 6325
rect 1814 6324 1819 6325
rect 1820 6324 1843 6325
rect 1824 6326 2293 6327
rect 1826 6328 1849 6329
rect 1827 6330 2541 6331
rect 1829 6332 1852 6333
rect 1830 6334 1833 6335
rect 1838 6334 1855 6335
rect 1844 6336 1891 6337
rect 1856 6338 1879 6339
rect 1860 6340 2799 6341
rect 1862 6342 1885 6343
rect 1866 6344 2217 6345
rect 1872 6346 2223 6347
rect 1874 6348 2017 6349
rect 1880 6350 2089 6351
rect 1886 6352 3452 6353
rect 1568 6354 1888 6355
rect 1892 6354 1951 6355
rect 1896 6356 1917 6357
rect 1898 6358 1909 6359
rect 1902 6360 1911 6361
rect 1904 6362 1939 6363
rect 1905 6364 1920 6365
rect 1914 6366 1941 6367
rect 1920 6368 1923 6369
rect 1928 6368 2083 6369
rect 1932 6370 1935 6371
rect 1944 6370 1947 6371
rect 1956 6370 1959 6371
rect 1962 6370 1971 6371
rect 1964 6372 1981 6373
rect 1974 6374 1995 6375
rect 1976 6376 2065 6377
rect 1982 6378 1993 6379
rect 1986 6380 2001 6381
rect 1998 6382 2019 6383
rect 1925 6384 2020 6385
rect 1445 6386 1927 6387
rect 1445 6388 1953 6389
rect 2004 6388 2007 6389
rect 2010 6388 2013 6389
rect 2022 6388 2025 6389
rect 2028 6388 2049 6389
rect 2030 6390 2235 6391
rect 2034 6392 2073 6393
rect 2036 6394 2071 6395
rect 2040 6396 2061 6397
rect 2042 6398 2053 6399
rect 2046 6400 2055 6401
rect 2058 6400 3362 6401
rect 2066 6402 3403 6403
rect 2076 6404 2091 6405
rect 1967 6406 2092 6407
rect 1968 6408 1989 6409
rect 2078 6408 3228 6409
rect 2084 6410 2161 6411
rect 2094 6412 2103 6413
rect 2100 6414 2109 6415
rect 2106 6416 2115 6417
rect 2112 6418 2127 6419
rect 2118 6420 2145 6421
rect 2120 6422 3290 6423
rect 2124 6424 3424 6425
rect 2130 6426 2133 6427
rect 2136 6426 2193 6427
rect 2138 6428 2173 6429
rect 2142 6430 2157 6431
rect 2148 6432 2151 6433
rect 2154 6432 2163 6433
rect 2168 6432 2179 6433
rect 2174 6434 2185 6435
rect 2181 6436 2568 6437
rect 2190 6438 2205 6439
rect 2196 6440 2325 6441
rect 2198 6442 2215 6443
rect 2202 6444 2319 6445
rect 2208 6446 2211 6447
rect 2220 6446 2229 6447
rect 2223 6448 2592 6449
rect 2226 6450 2295 6451
rect 2232 6452 2301 6453
rect 2238 6454 2355 6455
rect 2240 6456 2269 6457
rect 2244 6458 2265 6459
rect 2246 6460 2263 6461
rect 2250 6462 2253 6463
rect 2256 6462 2259 6463
rect 2270 6462 2275 6463
rect 2276 6462 2287 6463
rect 2282 6464 2299 6465
rect 2304 6464 2331 6465
rect 2306 6466 2311 6467
rect 2307 6468 2334 6469
rect 2312 6470 2317 6471
rect 2322 6470 2391 6471
rect 2328 6472 3406 6473
rect 2334 6474 2415 6475
rect 2336 6476 2347 6477
rect 2337 6478 2802 6479
rect 2342 6480 3445 6481
rect 2348 6482 2353 6483
rect 2358 6482 2661 6483
rect 2364 6484 2409 6485
rect 2366 6486 2377 6487
rect 2370 6488 2421 6489
rect 2372 6490 2395 6491
rect 2378 6492 2383 6493
rect 2384 6492 3269 6493
rect 2396 6494 2407 6495
rect 2400 6496 2403 6497
rect 2412 6496 3421 6497
rect 2418 6498 3301 6499
rect 2424 6500 2451 6501
rect 2426 6502 2431 6503
rect 1640 6504 2428 6505
rect 2432 6504 2437 6505
rect 2442 6504 2481 6505
rect 2444 6506 2449 6507
rect 2454 6506 2469 6507
rect 2460 6508 2709 6509
rect 2466 6510 2859 6511
rect 2472 6512 2487 6513
rect 2478 6514 2625 6515
rect 2484 6516 2583 6517
rect 2490 6518 2505 6519
rect 2492 6520 3396 6521
rect 2496 6522 2511 6523
rect 2498 6524 3399 6525
rect 2502 6526 2553 6527
rect 2508 6528 2529 6529
rect 2514 6530 2559 6531
rect 2516 6532 2521 6533
rect 2526 6532 2571 6533
rect 2532 6534 2577 6535
rect 2534 6536 3352 6537
rect 2538 6538 3276 6539
rect 2544 6540 2823 6541
rect 2550 6542 2763 6543
rect 2556 6544 2601 6545
rect 2562 6546 3167 6547
rect 2568 6548 2607 6549
rect 2574 6550 2619 6551
rect 2580 6552 2943 6553
rect 2586 6554 2631 6555
rect 2592 6556 2643 6557
rect 2594 6558 3157 6559
rect 2598 6560 2655 6561
rect 2604 6562 2667 6563
rect 2610 6564 2703 6565
rect 2616 6566 2673 6567
rect 2622 6568 2679 6569
rect 2628 6570 2685 6571
rect 2634 6572 2691 6573
rect 2640 6574 3359 6575
rect 2646 6576 2697 6577
rect 2652 6578 3366 6579
rect 2658 6580 3369 6581
rect 2664 6582 2715 6583
rect 2670 6584 2721 6585
rect 2676 6586 2733 6587
rect 2682 6588 2739 6589
rect 2688 6590 2745 6591
rect 2706 6592 2775 6593
rect 2712 6594 2865 6595
rect 2718 6596 2871 6597
rect 2724 6598 2787 6599
rect 2730 6600 2793 6601
rect 2736 6602 2811 6603
rect 2742 6604 2817 6605
rect 2748 6606 2829 6607
rect 2754 6608 2835 6609
rect 2766 6610 2841 6611
rect 2772 6612 2847 6613
rect 2778 6614 2901 6615
rect 2784 6616 2907 6617
rect 2790 6618 2913 6619
rect 1535 6620 2914 6621
rect 1536 6622 2769 6623
rect 2796 6622 2877 6623
rect 2802 6624 2883 6625
rect 2808 6626 2889 6627
rect 2820 6628 2919 6629
rect 2826 6630 2925 6631
rect 2832 6632 2931 6633
rect 2838 6634 2937 6635
rect 2850 6636 2949 6637
rect 2856 6638 2955 6639
rect 2859 6640 2958 6641
rect 2862 6642 2961 6643
rect 2868 6644 2967 6645
rect 2874 6646 2973 6647
rect 2877 6648 3297 6649
rect 2880 6650 2979 6651
rect 2886 6652 2991 6653
rect 2892 6654 3003 6655
rect 2898 6656 2997 6657
rect 2904 6658 3015 6659
rect 1748 6660 3016 6661
rect 2910 6662 3009 6663
rect 2916 6664 3021 6665
rect 2922 6666 3027 6667
rect 2928 6668 3442 6669
rect 2940 6670 3045 6671
rect 2946 6672 3057 6673
rect 2952 6674 3051 6675
rect 2958 6676 3039 6677
rect 2964 6678 3069 6679
rect 2970 6680 3075 6681
rect 2975 6682 3294 6683
rect 2976 6684 3063 6685
rect 2982 6686 3081 6687
rect 2988 6688 3087 6689
rect 2994 6690 3093 6691
rect 3000 6692 3099 6693
rect 3006 6694 3105 6695
rect 3012 6696 3111 6697
rect 3018 6698 3117 6699
rect 2852 6700 3118 6701
rect 3024 6702 3123 6703
rect 3036 6704 3240 6705
rect 3048 6706 3135 6707
rect 3054 6708 3153 6709
rect 3060 6710 3165 6711
rect 3066 6712 3171 6713
rect 3078 6714 3207 6715
rect 3081 6716 3210 6717
rect 3090 6718 3177 6719
rect 3102 6720 3189 6721
rect 3105 6722 3183 6723
rect 3108 6724 3219 6725
rect 3111 6726 3222 6727
rect 3113 6728 3355 6729
rect 3114 6730 3225 6731
rect 2780 6732 3225 6733
rect 3120 6734 3231 6735
rect 3123 6736 3234 6737
rect 3126 6738 3237 6739
rect 3030 6740 3237 6741
rect 3132 6742 3249 6743
rect 3140 6744 3280 6745
rect 3144 6746 3261 6747
rect 2756 6748 3262 6749
rect 3146 6750 3283 6751
rect 3147 6752 3264 6753
rect 2700 6754 3265 6755
rect 3150 6756 3267 6757
rect 3158 6758 3234 6759
rect 2984 6760 3160 6761
rect 3163 6760 3304 6761
rect 3169 6762 3286 6763
rect 2280 6764 3287 6765
rect 3181 6766 3310 6767
rect 3187 6768 3316 6769
rect 3193 6770 3322 6771
rect 3196 6772 3325 6773
rect 3200 6774 3431 6775
rect 1544 6776 3200 6777
rect 3203 6776 3428 6777
rect 2612 6778 3203 6779
rect 3211 6778 3340 6779
rect 3214 6780 3343 6781
rect 3217 6782 3349 6783
rect 3220 6784 3346 6785
rect 3230 6786 3372 6787
rect 3242 6788 3273 6789
rect 2388 6790 3272 6791
rect 3243 6792 3292 6793
rect 3246 6794 3375 6795
rect 3255 6796 3393 6797
rect 3258 6798 3378 6799
rect 3280 6800 3415 6801
rect 3283 6802 3418 6803
rect 3389 6804 3438 6805
rect 3434 6806 3449 6807
rect 1427 6815 1555 6816
rect 1434 6817 1531 6818
rect 1438 6819 1669 6820
rect 1441 6821 1663 6822
rect 1445 6823 2065 6824
rect 1448 6825 1852 6826
rect 1454 6827 1915 6828
rect 1472 6829 1921 6830
rect 1476 6831 2167 6832
rect 1417 6833 1476 6834
rect 1479 6833 2227 6834
rect 1478 6835 2161 6836
rect 1482 6837 2491 6838
rect 1503 6839 1615 6840
rect 1512 6841 2155 6842
rect 1512 6843 2224 6844
rect 1536 6845 2011 6846
rect 1524 6847 1537 6848
rect 1518 6849 1525 6850
rect 1542 6849 1555 6850
rect 1548 6851 2497 6852
rect 1551 6853 1993 6854
rect 1566 6855 1579 6856
rect 1424 6857 1567 6858
rect 1599 6857 2107 6858
rect 1608 6859 1612 6860
rect 1596 6861 1609 6862
rect 1596 6863 1957 6864
rect 1469 6865 1957 6866
rect 1463 6867 1470 6868
rect 1457 6869 1464 6870
rect 1620 6869 1639 6870
rect 1620 6871 2791 6872
rect 1623 6873 2095 6874
rect 1632 6875 1651 6876
rect 1644 6877 1663 6878
rect 1626 6879 1645 6880
rect 1500 6881 1627 6882
rect 1494 6883 1501 6884
rect 1698 6883 1705 6884
rect 1692 6885 1699 6886
rect 1431 6887 1693 6888
rect 1430 6889 1765 6890
rect 1749 6891 2485 6892
rect 1764 6893 1771 6894
rect 1433 6895 1771 6896
rect 1836 6895 3328 6896
rect 1836 6897 1873 6898
rect 1740 6899 1873 6900
rect 1423 6901 1741 6902
rect 1866 6901 1915 6902
rect 1806 6903 1867 6904
rect 1788 6905 1807 6906
rect 1776 6907 1789 6908
rect 1758 6909 1777 6910
rect 1746 6911 1759 6912
rect 1887 6911 1960 6912
rect 1905 6913 1972 6914
rect 1656 6915 1906 6916
rect 1920 6915 2443 6916
rect 1950 6917 1993 6918
rect 1878 6919 1951 6920
rect 1728 6921 1879 6922
rect 1728 6923 1735 6924
rect 1426 6925 1735 6926
rect 1980 6925 2011 6926
rect 1938 6927 1981 6928
rect 1884 6929 1939 6930
rect 1884 6931 3203 6932
rect 2001 6933 2020 6934
rect 2025 6933 2308 6934
rect 2034 6935 2107 6936
rect 1962 6937 2035 6938
rect 1902 6939 1963 6940
rect 1848 6941 1903 6942
rect 1812 6943 1849 6944
rect 1800 6945 1813 6946
rect 1800 6947 3157 6948
rect 2043 6949 2092 6950
rect 2058 6951 2155 6952
rect 1974 6953 2059 6954
rect 1974 6955 2017 6956
rect 1944 6957 2017 6958
rect 1944 6959 2137 6960
rect 2040 6961 2137 6962
rect 2040 6963 2089 6964
rect 2064 6965 3190 6966
rect 2070 6967 2095 6968
rect 1986 6969 2071 6970
rect 1908 6971 1987 6972
rect 1437 6973 1909 6974
rect 2100 6973 2167 6974
rect 2004 6975 2101 6976
rect 1932 6977 2005 6978
rect 1890 6979 1933 6980
rect 1854 6981 1891 6982
rect 1440 6983 1855 6984
rect 2112 6983 3287 6984
rect 2022 6985 2113 6986
rect 1451 6987 2023 6988
rect 2130 6987 2161 6988
rect 2046 6989 2131 6990
rect 1420 6991 2047 6992
rect 2181 6991 2194 6992
rect 2184 6993 2227 6994
rect 1485 6995 2185 6996
rect 2235 6995 3237 6996
rect 2280 6997 3267 6998
rect 2280 6999 2323 7000
rect 2286 7001 2323 7002
rect 2250 7003 2287 7004
rect 2190 7005 2251 7006
rect 2178 7007 2191 7008
rect 2178 7009 3290 7010
rect 2310 7011 3332 7012
rect 2262 7013 2311 7014
rect 2214 7015 2263 7016
rect 1515 7017 2215 7018
rect 2316 7017 3335 7018
rect 2274 7019 2317 7020
rect 2274 7021 2299 7022
rect 2244 7023 2299 7024
rect 2232 7025 2245 7026
rect 2220 7027 2233 7028
rect 2142 7029 2221 7030
rect 2052 7031 2143 7032
rect 1968 7033 2053 7034
rect 1896 7035 1969 7036
rect 1842 7037 1897 7038
rect 1842 7039 2305 7040
rect 2268 7041 2305 7042
rect 2268 7043 2869 7044
rect 2337 7045 2770 7046
rect 2358 7047 3200 7048
rect 2340 7049 2359 7050
rect 1827 7051 2341 7052
rect 2391 7051 2428 7052
rect 2406 7053 2443 7054
rect 2376 7055 2407 7056
rect 2352 7057 2377 7058
rect 2328 7059 2353 7060
rect 2292 7061 2329 7062
rect 2256 7063 2293 7064
rect 2238 7065 2257 7066
rect 2208 7067 2239 7068
rect 2118 7069 2209 7070
rect 2118 7071 2203 7072
rect 2124 7073 2203 7074
rect 2028 7075 2125 7076
rect 2028 7077 2083 7078
rect 1998 7079 2083 7080
rect 1926 7081 1999 7082
rect 1926 7083 3301 7084
rect 2448 7085 3277 7086
rect 2418 7087 2449 7088
rect 2394 7089 2419 7090
rect 2364 7091 2395 7092
rect 2364 7093 2371 7094
rect 2346 7095 2371 7096
rect 2334 7097 2347 7098
rect 1824 7099 2335 7100
rect 1824 7101 1831 7102
rect 1521 7103 1831 7104
rect 2472 7103 2491 7104
rect 2454 7105 2473 7106
rect 2436 7107 2455 7108
rect 2412 7109 2437 7110
rect 2382 7111 2413 7112
rect 2382 7113 3304 7114
rect 2478 7115 3160 7116
rect 2478 7117 2521 7118
rect 2484 7119 3274 7120
rect 2496 7121 2539 7122
rect 2502 7123 2521 7124
rect 1584 7125 2503 7126
rect 1572 7127 1585 7128
rect 1560 7129 1573 7130
rect 2526 7129 2539 7130
rect 2526 7131 2563 7132
rect 2466 7133 2563 7134
rect 1746 7135 2467 7136
rect 2568 7135 3164 7136
rect 2568 7137 3289 7138
rect 2574 7139 3286 7140
rect 2556 7141 2575 7142
rect 1587 7143 2557 7144
rect 2616 7143 3303 7144
rect 2616 7145 2629 7146
rect 2628 7147 2647 7148
rect 2646 7149 2665 7150
rect 2664 7151 2683 7152
rect 2676 7153 3269 7154
rect 2676 7155 3318 7156
rect 2694 7157 3265 7158
rect 2712 7159 2791 7160
rect 2712 7161 2725 7162
rect 2706 7163 2725 7164
rect 2706 7165 3321 7166
rect 2760 7167 3118 7168
rect 2838 7169 2869 7170
rect 1447 7171 2839 7172
rect 2859 7171 2890 7172
rect 2862 7173 3297 7174
rect 2832 7175 2863 7176
rect 2778 7177 2833 7178
rect 2772 7179 2779 7180
rect 2766 7181 2773 7182
rect 1860 7183 2767 7184
rect 1818 7185 1861 7186
rect 1518 7187 1819 7188
rect 2877 7187 2908 7188
rect 2886 7189 3225 7190
rect 2856 7191 2887 7192
rect 2826 7193 2857 7194
rect 2718 7195 2827 7196
rect 2544 7197 2719 7198
rect 2532 7199 2545 7200
rect 2508 7201 2533 7202
rect 2508 7203 2551 7204
rect 1444 7205 2551 7206
rect 2895 7205 2914 7206
rect 2904 7207 2935 7208
rect 2874 7209 2905 7210
rect 2844 7211 2875 7212
rect 2784 7213 2845 7214
rect 2580 7215 2785 7216
rect 2580 7217 2593 7218
rect 2592 7219 2599 7220
rect 2598 7221 2611 7222
rect 2610 7223 2623 7224
rect 2622 7225 2641 7226
rect 2640 7227 2653 7228
rect 2652 7229 2671 7230
rect 2670 7231 2701 7232
rect 2700 7233 2731 7234
rect 2730 7235 2737 7236
rect 2736 7237 2743 7238
rect 1539 7239 2743 7240
rect 2940 7239 3296 7240
rect 2898 7241 2941 7242
rect 2892 7243 2899 7244
rect 2892 7245 2911 7246
rect 2880 7247 2911 7248
rect 2850 7249 2881 7250
rect 2820 7251 2851 7252
rect 2802 7253 2821 7254
rect 2796 7255 2803 7256
rect 2796 7257 3262 7258
rect 2964 7259 2992 7260
rect 2946 7261 2965 7262
rect 2916 7263 2947 7264
rect 2916 7265 3263 7266
rect 3006 7267 3043 7268
rect 3006 7269 3013 7270
rect 2982 7271 3013 7272
rect 3009 7273 3016 7274
rect 3030 7273 3073 7274
rect 3030 7275 3300 7276
rect 3036 7277 3142 7278
rect 3000 7279 3037 7280
rect 2958 7281 3001 7282
rect 3048 7281 3085 7282
rect 2976 7283 3049 7284
rect 2922 7285 2977 7286
rect 3066 7285 3097 7286
rect 3024 7287 3067 7288
rect 2994 7289 3025 7290
rect 2994 7291 3082 7292
rect 3078 7293 3157 7294
rect 3105 7295 3136 7296
rect 3108 7297 3139 7298
rect 3111 7299 3240 7300
rect 3123 7301 3154 7302
rect 3132 7303 3163 7304
rect 3102 7305 3133 7306
rect 3102 7307 3234 7308
rect 3144 7309 3175 7310
rect 3147 7311 3178 7312
rect 3159 7313 3228 7314
rect 3166 7315 3312 7316
rect 3169 7317 3200 7318
rect 3181 7319 3224 7320
rect 3150 7321 3181 7322
rect 3120 7323 3151 7324
rect 3090 7325 3121 7326
rect 3060 7327 3091 7328
rect 3054 7329 3061 7330
rect 3018 7331 3055 7332
rect 2988 7333 3019 7334
rect 2970 7335 2989 7336
rect 2952 7337 2971 7338
rect 2928 7339 2953 7340
rect 3193 7339 3236 7340
rect 2922 7341 3194 7342
rect 3196 7341 3239 7342
rect 2928 7343 3197 7344
rect 3205 7343 3244 7344
rect 3114 7345 3245 7346
rect 3211 7347 3254 7348
rect 3217 7349 3242 7350
rect 3220 7351 3270 7352
rect 3255 7353 3325 7354
rect 3214 7355 3257 7356
rect 3258 7355 3272 7356
rect 3126 7357 3260 7358
rect 3280 7357 3294 7358
rect 2958 7359 3293 7360
rect 3230 7361 3280 7362
rect 3187 7363 3230 7364
rect 2088 7365 3187 7366
rect 3283 7365 3315 7366
rect 3246 7367 3283 7368
rect 1423 7376 1729 7377
rect 1423 7378 1849 7379
rect 1430 7380 1777 7381
rect 1433 7382 1645 7383
rect 1437 7384 1464 7385
rect 1438 7386 1987 7387
rect 1444 7388 1470 7389
rect 1445 7390 1573 7391
rect 1447 7392 2761 7393
rect 1449 7394 1537 7395
rect 1451 7396 2107 7397
rect 1452 7398 1531 7399
rect 1454 7400 1795 7401
rect 1461 7402 1729 7403
rect 1464 7404 1807 7405
rect 1468 7406 1753 7407
rect 1475 7408 1572 7409
rect 1478 7410 2191 7411
rect 1480 7412 1501 7413
rect 1482 7414 1981 7415
rect 1485 7416 2896 7417
rect 1492 7418 3082 7419
rect 1504 7420 1513 7421
rect 1510 7422 1555 7423
rect 1442 7424 1554 7425
rect 1513 7426 2215 7427
rect 1518 7428 2995 7429
rect 1517 7430 1639 7431
rect 1521 7432 1525 7433
rect 1523 7434 1621 7435
rect 1551 7436 2533 7437
rect 1559 7438 1579 7439
rect 1580 7438 2881 7439
rect 1589 7440 1609 7441
rect 1599 7442 2161 7443
rect 1602 7444 2299 7445
rect 1605 7446 2257 7447
rect 1614 7448 1627 7449
rect 1623 7450 2479 7451
rect 1626 7452 1663 7453
rect 1644 7454 3001 7455
rect 1656 7456 2269 7457
rect 1662 7458 2563 7459
rect 1520 7460 2563 7461
rect 1668 7462 1717 7463
rect 1692 7464 1753 7465
rect 1710 7466 2368 7467
rect 1686 7468 1711 7469
rect 1650 7470 1687 7471
rect 1650 7472 3007 7473
rect 1716 7474 3091 7475
rect 1746 7476 2635 7477
rect 1746 7478 2917 7479
rect 1749 7480 2911 7481
rect 1776 7482 2785 7483
rect 1782 7484 1849 7485
rect 1782 7486 2869 7487
rect 1794 7488 2863 7489
rect 1806 7490 2719 7491
rect 1824 7492 1987 7493
rect 1722 7494 1825 7495
rect 1722 7496 2941 7497
rect 1896 7498 2107 7499
rect 1788 7500 1897 7501
rect 1471 7502 1789 7503
rect 1905 7502 2116 7503
rect 1959 7504 2284 7505
rect 1974 7506 2161 7507
rect 1974 7508 2833 7509
rect 1980 7510 2851 7511
rect 2001 7512 2278 7513
rect 2016 7514 2299 7515
rect 2016 7516 2467 7517
rect 2025 7518 2314 7519
rect 2028 7520 2257 7521
rect 2028 7522 2737 7523
rect 2043 7524 2290 7525
rect 2100 7526 3185 7527
rect 2100 7528 2389 7529
rect 2088 7530 2389 7531
rect 1890 7532 2089 7533
rect 1764 7534 1891 7535
rect 2190 7534 2359 7535
rect 2064 7536 2359 7537
rect 2064 7538 2641 7539
rect 2193 7540 2296 7541
rect 2208 7542 2479 7543
rect 1950 7544 2209 7545
rect 1812 7546 1951 7547
rect 1812 7548 1879 7549
rect 1818 7550 1879 7551
rect 1548 7552 1819 7553
rect 1547 7554 1567 7555
rect 1565 7556 1585 7557
rect 2214 7556 2551 7557
rect 2235 7558 2356 7559
rect 1971 7560 2236 7561
rect 2238 7560 2467 7561
rect 1992 7562 2239 7563
rect 1836 7564 1993 7565
rect 1598 7566 1837 7567
rect 2244 7566 3187 7567
rect 1440 7568 2245 7569
rect 2268 7568 2275 7569
rect 1998 7570 2275 7571
rect 1842 7572 1999 7573
rect 1758 7574 1843 7575
rect 1698 7576 1759 7577
rect 1698 7578 1705 7579
rect 2286 7578 2533 7579
rect 2004 7580 2287 7581
rect 2004 7582 2725 7583
rect 2316 7584 3190 7585
rect 2316 7586 2353 7587
rect 2052 7588 2353 7589
rect 1854 7590 2053 7591
rect 1426 7592 1855 7593
rect 1426 7594 1867 7595
rect 1740 7596 1867 7597
rect 1680 7598 1741 7599
rect 1680 7600 2893 7601
rect 2337 7602 2392 7603
rect 2361 7604 2770 7605
rect 2406 7606 3277 7607
rect 2166 7608 2407 7609
rect 2166 7610 2281 7611
rect 2280 7612 3188 7613
rect 2412 7614 3213 7615
rect 2124 7616 2413 7617
rect 1926 7618 2125 7619
rect 1926 7620 2557 7621
rect 2394 7622 2557 7623
rect 2130 7624 2395 7625
rect 2076 7626 2131 7627
rect 1914 7628 2077 7629
rect 1914 7630 2743 7631
rect 2454 7632 2551 7633
rect 2322 7634 2455 7635
rect 2034 7636 2323 7637
rect 2034 7638 3171 7639
rect 2460 7640 3267 7641
rect 2172 7642 2461 7643
rect 1938 7644 2173 7645
rect 1938 7646 2791 7647
rect 2472 7648 3263 7649
rect 2202 7650 2473 7651
rect 1956 7652 2203 7653
rect 1920 7654 1957 7655
rect 1920 7656 2503 7657
rect 2340 7658 2503 7659
rect 2046 7660 2341 7661
rect 1435 7662 2047 7663
rect 2490 7662 2641 7663
rect 2262 7664 2491 7665
rect 2040 7666 2263 7667
rect 2040 7668 2527 7669
rect 2508 7670 3167 7671
rect 2304 7672 2509 7673
rect 2094 7674 2305 7675
rect 1908 7676 2095 7677
rect 1770 7678 1909 7679
rect 1770 7680 2875 7681
rect 2514 7682 3145 7683
rect 2514 7684 2545 7685
rect 2310 7686 2545 7687
rect 2022 7688 2311 7689
rect 2022 7690 2497 7691
rect 2250 7692 2497 7693
rect 2010 7694 2251 7695
rect 2010 7696 2839 7697
rect 2526 7698 3270 7699
rect 2538 7700 2635 7701
rect 2292 7702 2539 7703
rect 2184 7704 2293 7705
rect 2184 7706 2233 7707
rect 1968 7708 2233 7709
rect 1968 7710 3274 7711
rect 2610 7712 3300 7713
rect 2424 7714 2611 7715
rect 2136 7716 2425 7717
rect 2118 7718 2137 7719
rect 2118 7720 2365 7721
rect 1596 7722 2365 7723
rect 1595 7724 2833 7725
rect 2616 7726 3303 7727
rect 2436 7728 2617 7729
rect 2196 7730 2437 7731
rect 2196 7732 2581 7733
rect 2370 7734 2581 7735
rect 2646 7734 2725 7735
rect 2664 7736 2737 7737
rect 2568 7738 2665 7739
rect 2568 7740 3328 7741
rect 2670 7742 2743 7743
rect 2670 7744 3289 7745
rect 2682 7746 3325 7747
rect 2688 7748 3321 7749
rect 2574 7750 2689 7751
rect 2520 7752 2575 7753
rect 2484 7754 2521 7755
rect 2220 7756 2485 7757
rect 2148 7758 2221 7759
rect 1932 7760 2149 7761
rect 1932 7762 2401 7763
rect 2142 7764 2401 7765
rect 2142 7766 3335 7767
rect 2694 7768 3148 7769
rect 2604 7770 2695 7771
rect 2604 7772 3210 7773
rect 2700 7774 2719 7775
rect 2622 7776 2701 7777
rect 2442 7778 2623 7779
rect 2334 7780 2443 7781
rect 2058 7782 2335 7783
rect 1860 7784 2059 7785
rect 1734 7786 1861 7787
rect 1674 7788 1735 7789
rect 1577 7790 1675 7791
rect 2706 7790 2761 7791
rect 2628 7792 2707 7793
rect 2448 7794 2629 7795
rect 2178 7796 2449 7797
rect 2178 7798 2347 7799
rect 2070 7800 2347 7801
rect 1884 7802 2071 7803
rect 1800 7804 1885 7805
rect 1800 7806 2857 7807
rect 2754 7808 3016 7809
rect 2784 7810 2845 7811
rect 2790 7812 2797 7813
rect 2772 7814 2797 7815
rect 2748 7816 2773 7817
rect 2676 7818 2749 7819
rect 2586 7820 2677 7821
rect 2376 7822 2587 7823
rect 2112 7824 2377 7825
rect 1902 7826 2113 7827
rect 1830 7828 1903 7829
rect 1830 7830 1873 7831
rect 1872 7832 2767 7833
rect 2712 7834 2767 7835
rect 2658 7836 2713 7837
rect 2592 7838 2659 7839
rect 2418 7840 2593 7841
rect 2328 7842 2419 7843
rect 2226 7844 2329 7845
rect 1962 7846 2227 7847
rect 1962 7848 3332 7849
rect 2814 7850 2821 7851
rect 2835 7850 3010 7851
rect 2838 7852 2947 7853
rect 2844 7854 2977 7855
rect 2850 7856 2899 7857
rect 2856 7858 2923 7859
rect 2862 7860 2887 7861
rect 2865 7862 2890 7863
rect 2868 7864 2929 7865
rect 2874 7866 3097 7867
rect 2880 7868 2905 7869
rect 2883 7870 2908 7871
rect 2886 7872 3130 7873
rect 2892 7874 3157 7875
rect 2895 7876 3160 7877
rect 2898 7878 3013 7879
rect 2904 7880 2959 7881
rect 2910 7882 2953 7883
rect 2916 7884 3296 7885
rect 2922 7886 2971 7887
rect 2928 7888 3019 7889
rect 2934 7890 3197 7891
rect 2940 7892 2989 7893
rect 2943 7894 2992 7895
rect 2946 7896 3031 7897
rect 2952 7898 3260 7899
rect 2958 7900 3025 7901
rect 2964 7902 3293 7903
rect 2964 7904 3318 7905
rect 2970 7906 3037 7907
rect 2976 7908 3043 7909
rect 2982 7910 3067 7911
rect 2370 7912 3067 7913
rect 2988 7914 3073 7915
rect 2994 7916 3142 7917
rect 3000 7918 3085 7919
rect 3006 7920 3151 7921
rect 3009 7922 3055 7923
rect 3012 7924 3245 7925
rect 3018 7926 3103 7927
rect 3030 7928 3139 7929
rect 3033 7930 3070 7931
rect 3036 7932 3121 7933
rect 3048 7934 3127 7935
rect 3048 7936 3133 7937
rect 3051 7938 3136 7939
rect 3054 7940 3163 7941
rect 3060 7942 3164 7943
rect 3060 7944 3178 7945
rect 3063 7946 3175 7947
rect 2730 7948 3174 7949
rect 2652 7950 2731 7951
rect 2652 7952 3203 7953
rect 3072 7954 3181 7955
rect 2646 7956 3181 7957
rect 3078 7958 3154 7959
rect 3084 7960 3200 7961
rect 3096 7962 3206 7963
rect 2382 7964 3206 7965
rect 2082 7966 2383 7967
rect 2082 7968 2599 7969
rect 2430 7970 2599 7971
rect 2154 7972 2431 7973
rect 1944 7974 2155 7975
rect 1944 7976 2827 7977
rect 2808 7978 2827 7979
rect 2802 7980 2809 7981
rect 2778 7982 2803 7983
rect 3108 7982 3224 7983
rect 3114 7984 3230 7985
rect 3120 7986 3236 7987
rect 3123 7988 3239 7989
rect 3138 7990 3254 7991
rect 3141 7992 3152 7993
rect 3154 7992 3257 7993
rect 3157 7994 3280 7995
rect 3160 7996 3283 7997
rect 3177 7998 3242 7999
rect 3193 8000 3286 8001
rect 3196 8002 3312 8003
rect 3199 8004 3315 8005
rect 1423 8013 1441 8014
rect 1423 8015 2209 8016
rect 1426 8017 2047 8018
rect 1430 8019 1489 8020
rect 1433 8021 1493 8022
rect 1438 8023 1927 8024
rect 1445 8025 2290 8026
rect 1444 8027 2323 8028
rect 1452 8029 1524 8030
rect 1454 8031 1891 8032
rect 1461 8033 1831 8034
rect 1464 8035 1813 8036
rect 1463 8037 1897 8038
rect 1437 8039 1897 8040
rect 1466 8041 1813 8042
rect 1468 8043 1548 8044
rect 1471 8045 1576 8046
rect 1480 8047 1495 8048
rect 1504 8047 1507 8048
rect 1510 8047 2371 8048
rect 1520 8049 2359 8050
rect 1524 8051 1765 8052
rect 1527 8053 1915 8054
rect 1548 8055 1554 8056
rect 1554 8057 1560 8058
rect 1560 8059 1566 8060
rect 1566 8061 1572 8062
rect 1572 8063 1651 8064
rect 1577 8065 3052 8066
rect 1584 8067 1590 8068
rect 1590 8069 1627 8070
rect 1593 8071 3055 8072
rect 1595 8073 1801 8074
rect 1598 8075 1795 8076
rect 1602 8077 2455 8078
rect 1602 8079 1615 8080
rect 1614 8081 1675 8082
rect 1620 8083 1687 8084
rect 1638 8085 1699 8086
rect 1650 8087 1735 8088
rect 1656 8089 1693 8090
rect 1656 8091 1741 8092
rect 1662 8093 1699 8094
rect 1662 8095 1669 8096
rect 1668 8097 1753 8098
rect 1674 8099 1759 8100
rect 1686 8101 1729 8102
rect 1704 8103 1789 8104
rect 1716 8105 2779 8106
rect 1716 8107 1777 8108
rect 1722 8109 2746 8110
rect 1722 8111 1807 8112
rect 1451 8113 1807 8114
rect 1728 8115 1819 8116
rect 1734 8117 1825 8118
rect 1740 8119 1783 8120
rect 1752 8121 1843 8122
rect 1758 8123 1849 8124
rect 1776 8125 1855 8126
rect 1782 8127 1861 8128
rect 1788 8129 1867 8130
rect 1794 8131 1903 8132
rect 1800 8133 1885 8134
rect 1818 8135 1879 8136
rect 1824 8137 1921 8138
rect 1830 8139 1945 8140
rect 1842 8141 1909 8142
rect 1836 8143 1909 8144
rect 1836 8145 1933 8146
rect 1848 8147 1975 8148
rect 1854 8149 1981 8150
rect 1860 8151 2011 8152
rect 1866 8153 2785 8154
rect 1878 8155 1963 8156
rect 1884 8157 1969 8158
rect 1890 8159 1951 8160
rect 1902 8161 2005 8162
rect 1473 8163 2005 8164
rect 1914 8165 2773 8166
rect 1926 8167 2035 8168
rect 1932 8169 3185 8170
rect 1944 8171 1993 8172
rect 1950 8173 1999 8174
rect 1962 8175 2017 8176
rect 1968 8177 2023 8178
rect 1974 8179 2761 8180
rect 1980 8181 2041 8182
rect 1992 8183 2053 8184
rect 1998 8185 2059 8186
rect 2010 8187 2083 8188
rect 2016 8189 2071 8190
rect 2022 8191 2077 8192
rect 2028 8193 3171 8194
rect 2028 8195 2683 8196
rect 2034 8197 2101 8198
rect 2040 8199 2089 8200
rect 2046 8201 2107 8202
rect 2052 8203 2113 8204
rect 2055 8205 2116 8206
rect 2058 8207 2095 8208
rect 2064 8209 3042 8210
rect 2064 8211 2119 8212
rect 1447 8213 2119 8214
rect 2070 8215 2143 8216
rect 2076 8217 2125 8218
rect 2082 8219 2131 8220
rect 2088 8221 2137 8222
rect 2094 8223 2155 8224
rect 2100 8225 2149 8226
rect 2106 8227 2179 8228
rect 2112 8229 2161 8230
rect 1580 8231 2161 8232
rect 2124 8233 2197 8234
rect 2130 8235 2185 8236
rect 2136 8237 3024 8238
rect 2142 8239 2191 8240
rect 1426 8241 2191 8242
rect 2148 8243 2173 8244
rect 2154 8245 2653 8246
rect 2166 8247 3203 8248
rect 2166 8249 2269 8250
rect 2172 8251 2215 8252
rect 1435 8253 2215 8254
rect 2178 8255 2521 8256
rect 2184 8257 2203 8258
rect 2196 8259 2221 8260
rect 2202 8261 2515 8262
rect 2208 8263 2293 8264
rect 2220 8265 2227 8266
rect 2226 8267 2233 8268
rect 2229 8269 2236 8270
rect 2232 8271 2239 8272
rect 2238 8273 2245 8274
rect 2244 8275 2251 8276
rect 2250 8277 2257 8278
rect 2256 8279 2263 8280
rect 2262 8281 2503 8282
rect 2268 8283 2275 8284
rect 2271 8285 2278 8286
rect 1442 8287 2278 8288
rect 2274 8289 2287 8290
rect 2280 8291 2287 8292
rect 1515 8293 2281 8294
rect 2283 8293 2290 8294
rect 2292 8293 2305 8294
rect 2298 8295 2305 8296
rect 2298 8297 2419 8298
rect 2313 8299 2332 8300
rect 2316 8301 3070 8302
rect 2316 8303 2365 8304
rect 2319 8305 3076 8306
rect 2322 8307 2443 8308
rect 1605 8309 2443 8310
rect 2337 8311 2350 8312
rect 2295 8313 2338 8314
rect 2346 8313 2359 8314
rect 2334 8315 2347 8316
rect 1470 8317 2335 8318
rect 2352 8317 2365 8318
rect 2340 8319 2353 8320
rect 2340 8321 2377 8322
rect 2370 8323 2395 8324
rect 2376 8325 2401 8326
rect 2382 8327 2395 8328
rect 2382 8329 2551 8330
rect 2400 8331 2491 8332
rect 2418 8333 2431 8334
rect 2424 8335 2431 8336
rect 2412 8337 2425 8338
rect 2412 8339 3148 8340
rect 2454 8341 2467 8342
rect 2466 8343 2557 8344
rect 2490 8345 2509 8346
rect 2496 8347 2957 8348
rect 2496 8349 2563 8350
rect 2502 8351 2575 8352
rect 2508 8353 2527 8354
rect 2514 8355 2569 8356
rect 2520 8357 2533 8358
rect 2526 8359 2539 8360
rect 2532 8361 2599 8362
rect 2538 8363 3181 8364
rect 2544 8365 3021 8366
rect 2544 8367 2593 8368
rect 2550 8369 2617 8370
rect 2556 8371 2611 8372
rect 2562 8373 2581 8374
rect 2568 8375 2587 8376
rect 2574 8377 2623 8378
rect 2586 8379 2605 8380
rect 2592 8381 2629 8382
rect 2604 8383 2641 8384
rect 2610 8385 2647 8386
rect 2616 8387 2659 8388
rect 2622 8389 2671 8390
rect 2628 8391 2665 8392
rect 2640 8393 2695 8394
rect 2646 8395 2701 8396
rect 2652 8397 2707 8398
rect 2658 8399 2737 8400
rect 2664 8401 2743 8402
rect 1746 8403 2743 8404
rect 1746 8405 1873 8406
rect 1872 8407 1957 8408
rect 1956 8409 2719 8410
rect 2670 8411 2725 8412
rect 2682 8413 2749 8414
rect 2694 8415 2797 8416
rect 2700 8417 2803 8418
rect 2706 8419 2809 8420
rect 2724 8421 2827 8422
rect 2733 8423 2836 8424
rect 2736 8425 2851 8426
rect 1517 8427 2851 8428
rect 1449 8429 1519 8430
rect 2748 8429 2863 8430
rect 2751 8431 2866 8432
rect 2754 8433 2869 8434
rect 2769 8435 3210 8436
rect 2772 8437 2845 8438
rect 2775 8439 2839 8440
rect 2784 8441 2887 8442
rect 2796 8443 2911 8444
rect 2802 8445 3127 8446
rect 2808 8447 2923 8448
rect 2826 8449 2941 8450
rect 2829 8451 2944 8452
rect 2832 8453 3174 8454
rect 2832 8455 2971 8456
rect 2838 8457 2947 8458
rect 2856 8459 3067 8460
rect 2856 8461 2977 8462
rect 2862 8463 2875 8464
rect 2874 8465 3001 8466
rect 2883 8467 3206 8468
rect 2898 8469 3167 8470
rect 2898 8471 3013 8472
rect 2598 8473 3012 8474
rect 2901 8475 3016 8476
rect 2910 8477 3019 8478
rect 2916 8479 3178 8480
rect 2916 8481 3034 8482
rect 2712 8483 3035 8484
rect 2712 8485 2815 8486
rect 2814 8487 2929 8488
rect 2919 8489 2995 8490
rect 2928 8491 3049 8492
rect 2931 8493 2965 8494
rect 2934 8495 3064 8496
rect 2937 8497 2950 8498
rect 2940 8499 3073 8500
rect 2730 8501 3073 8502
rect 1644 8503 2731 8504
rect 1644 8505 1711 8506
rect 1680 8507 1711 8508
rect 1680 8509 2368 8510
rect 2355 8511 2368 8512
rect 2946 8511 3061 8512
rect 2952 8513 3069 8514
rect 2406 8515 2954 8516
rect 2388 8517 2407 8518
rect 2388 8519 2437 8520
rect 2436 8521 3145 8522
rect 2958 8523 3066 8524
rect 2959 8525 3085 8526
rect 2971 8527 3124 8528
rect 2986 8529 3002 8530
rect 2995 8531 3152 8532
rect 2998 8533 3142 8534
rect 3004 8535 3121 8536
rect 3006 8537 3082 8538
rect 2982 8539 3083 8540
rect 3009 8541 3130 8542
rect 2634 8543 3009 8544
rect 2634 8545 2677 8546
rect 1770 8547 2677 8548
rect 1770 8549 1939 8550
rect 1938 8551 1987 8552
rect 1986 8553 2767 8554
rect 2766 8555 2881 8556
rect 2880 8557 2989 8558
rect 3014 8557 3158 8558
rect 3017 8559 3161 8560
rect 3027 8561 3097 8562
rect 3036 8563 3213 8564
rect 2983 8565 3038 8566
rect 3044 8565 3115 8566
rect 3047 8567 3200 8568
rect 3059 8569 3079 8570
rect 2688 8571 3080 8572
rect 2688 8573 2791 8574
rect 2790 8575 2905 8576
rect 2904 8577 3164 8578
rect 3062 8579 3197 8580
rect 3108 8581 3188 8582
rect 3138 8583 3155 8584
rect 1423 8592 2185 8593
rect 1423 8594 2005 8595
rect 1426 8596 1681 8597
rect 1426 8598 1999 8599
rect 1430 8600 2189 8601
rect 1430 8602 2227 8603
rect 1433 8604 2230 8605
rect 1437 8606 2233 8607
rect 1440 8608 1445 8609
rect 1444 8610 1657 8611
rect 1447 8612 1759 8613
rect 1433 8614 1448 8615
rect 1451 8614 1693 8615
rect 1451 8616 1771 8617
rect 1454 8618 1694 8619
rect 1454 8620 1777 8621
rect 1461 8622 2734 8623
rect 1466 8624 1801 8625
rect 1470 8626 2359 8627
rect 1470 8628 1939 8629
rect 1473 8630 1940 8631
rect 1473 8632 2245 8633
rect 1458 8634 2246 8635
rect 1494 8636 1501 8637
rect 1488 8638 1495 8639
rect 1512 8638 1981 8639
rect 1506 8640 1513 8641
rect 1506 8642 3038 8643
rect 1515 8644 1535 8645
rect 1524 8646 1747 8647
rect 1531 8648 1963 8649
rect 1543 8650 1567 8651
rect 1552 8652 1885 8653
rect 1560 8654 1568 8655
rect 1554 8656 1562 8657
rect 1584 8656 1598 8657
rect 1588 8658 1628 8659
rect 1602 8660 1610 8661
rect 1620 8660 2267 8661
rect 1614 8662 1622 8663
rect 1644 8662 1658 8663
rect 1638 8664 1646 8665
rect 1674 8664 1682 8665
rect 1668 8666 1676 8667
rect 1662 8668 1670 8669
rect 1650 8670 1664 8671
rect 1585 8672 1652 8673
rect 1722 8672 1748 8673
rect 1723 8674 1735 8675
rect 1716 8676 1736 8677
rect 1717 8678 1729 8679
rect 1729 8680 2731 8681
rect 1740 8682 1802 8683
rect 1741 8684 1753 8685
rect 1527 8686 1754 8687
rect 1527 8688 2290 8689
rect 1759 8690 1783 8691
rect 1764 8692 1772 8693
rect 1765 8694 1789 8695
rect 1463 8696 1790 8697
rect 1777 8698 1795 8699
rect 1783 8700 1807 8701
rect 1795 8702 1819 8703
rect 1807 8704 1825 8705
rect 1819 8706 1831 8707
rect 1825 8708 1855 8709
rect 1831 8710 1909 8711
rect 1848 8712 2976 8713
rect 1849 8714 1867 8715
rect 1855 8716 1879 8717
rect 1867 8718 1897 8719
rect 1879 8720 1903 8721
rect 1894 8722 1915 8723
rect 1897 8724 2677 8725
rect 1903 8726 1927 8727
rect 1909 8728 1933 8729
rect 1915 8730 1945 8731
rect 1921 8732 1951 8733
rect 1927 8734 1957 8735
rect 1933 8736 1975 8737
rect 1945 8738 1969 8739
rect 1951 8740 2011 8741
rect 1957 8742 1993 8743
rect 1963 8744 2029 8745
rect 1969 8746 2017 8747
rect 1975 8748 2023 8749
rect 1981 8750 2924 8751
rect 1993 8752 2065 8753
rect 1572 8754 2066 8755
rect 1548 8756 1574 8757
rect 1549 8758 1813 8759
rect 1813 8760 1843 8761
rect 1843 8762 1861 8763
rect 1861 8764 1891 8765
rect 1999 8764 2041 8765
rect 2005 8766 2047 8767
rect 2011 8768 2053 8769
rect 2014 8770 2056 8771
rect 2017 8772 2059 8773
rect 2023 8774 2035 8775
rect 2029 8776 2107 8777
rect 2032 8778 2362 8779
rect 2035 8780 2077 8781
rect 2041 8782 2083 8783
rect 2047 8784 2095 8785
rect 2053 8786 2101 8787
rect 2059 8788 2089 8789
rect 2070 8790 2102 8791
rect 2071 8792 2113 8793
rect 2077 8794 2119 8795
rect 2083 8796 2647 8797
rect 2089 8798 2131 8799
rect 2095 8800 2137 8801
rect 1440 8802 2138 8803
rect 2107 8804 2143 8805
rect 2113 8806 2161 8807
rect 2119 8808 2167 8809
rect 2124 8810 2132 8811
rect 2125 8812 2149 8813
rect 2143 8814 2179 8815
rect 2149 8816 2617 8817
rect 2161 8818 2197 8819
rect 2167 8820 2191 8821
rect 2179 8822 2323 8823
rect 2185 8824 2215 8825
rect 2191 8826 2209 8827
rect 2197 8828 2257 8829
rect 2202 8830 3012 8831
rect 2203 8832 2281 8833
rect 2209 8834 2299 8835
rect 2215 8836 2467 8837
rect 2227 8838 2311 8839
rect 2233 8840 2293 8841
rect 1593 8842 2294 8843
rect 2250 8844 3045 8845
rect 2251 8846 2269 8847
rect 2254 8848 2272 8849
rect 2257 8850 2275 8851
rect 2260 8852 2278 8853
rect 2262 8854 2853 8855
rect 2263 8856 2287 8857
rect 2269 8858 2503 8859
rect 2275 8860 2443 8861
rect 2281 8862 2317 8863
rect 1575 8864 2318 8865
rect 2287 8866 2305 8867
rect 2299 8868 2957 8869
rect 2305 8870 2335 8871
rect 2308 8872 2338 8873
rect 2311 8874 2329 8875
rect 2314 8876 2332 8877
rect 2319 8878 2357 8879
rect 2323 8880 2347 8881
rect 2326 8882 2350 8883
rect 2329 8884 2341 8885
rect 2335 8886 2353 8887
rect 2341 8888 2365 8889
rect 2344 8890 2368 8891
rect 2347 8892 2389 8893
rect 2353 8894 2962 8895
rect 2359 8896 2371 8897
rect 2365 8898 2377 8899
rect 2371 8900 2395 8901
rect 2377 8902 2491 8903
rect 2389 8904 2455 8905
rect 2395 8906 2413 8907
rect 2400 8908 2954 8909
rect 2401 8910 2419 8911
rect 2413 8912 2431 8913
rect 2419 8914 2437 8915
rect 2431 8916 2449 8917
rect 2437 8918 2461 8919
rect 2443 8920 2515 8921
rect 2449 8922 2509 8923
rect 2455 8924 2485 8925
rect 2461 8926 2473 8927
rect 2467 8928 2479 8929
rect 2473 8930 2545 8931
rect 2479 8932 2533 8933
rect 2485 8934 2551 8935
rect 2491 8936 2521 8937
rect 2496 8938 3009 8939
rect 2497 8940 2527 8941
rect 2503 8942 2539 8943
rect 2509 8944 2557 8945
rect 2515 8946 2593 8947
rect 2521 8948 2563 8949
rect 2527 8950 2569 8951
rect 2533 8952 2599 8953
rect 2536 8954 2902 8955
rect 2539 8956 2770 8957
rect 2545 8958 2587 8959
rect 2551 8960 2605 8961
rect 2557 8962 2611 8963
rect 2563 8964 2623 8965
rect 2569 8966 2629 8967
rect 2574 8968 3035 8969
rect 2575 8970 2635 8971
rect 2581 8972 2653 8973
rect 2593 8974 2665 8975
rect 2605 8976 3080 8977
rect 2611 8978 2671 8979
rect 2617 8980 2801 8981
rect 2620 8982 2896 8983
rect 2623 8984 2689 8985
rect 2629 8986 2695 8987
rect 2635 8988 2701 8989
rect 2653 8990 2752 8991
rect 2656 8992 2725 8993
rect 2658 8994 3073 8995
rect 2659 8996 2849 8997
rect 2665 8998 2737 8999
rect 2671 9000 2743 9001
rect 2677 9002 2755 9003
rect 2695 9004 2767 9005
rect 2698 9006 3083 9007
rect 2701 9008 2773 9009
rect 2704 9010 2776 9011
rect 2719 9012 2797 9013
rect 2722 9014 2902 9015
rect 2725 9016 2863 9017
rect 2731 9018 2969 9019
rect 2737 9020 2809 9021
rect 2743 9022 2785 9023
rect 2761 9024 2827 9025
rect 2764 9026 2830 9027
rect 2767 9028 2833 9029
rect 2773 9030 2851 9031
rect 2785 9032 2803 9033
rect 2797 9034 2893 9035
rect 2818 9036 2920 9037
rect 2332 9038 2921 9039
rect 2821 9040 2905 9041
rect 2682 9042 2905 9043
rect 2683 9044 2746 9045
rect 2827 9044 2911 9045
rect 2833 9046 2950 9047
rect 2836 9048 2938 9049
rect 2790 9050 2938 9051
rect 2838 9052 3066 9053
rect 2839 9054 2941 9055
rect 2845 9056 3076 9057
rect 2856 9058 2892 9059
rect 2220 9060 2856 9061
rect 2221 9062 2239 9063
rect 1524 9064 2240 9065
rect 2858 9064 2960 9065
rect 2748 9066 2959 9067
rect 2749 9068 2815 9069
rect 2815 9070 3031 9071
rect 2870 9072 2972 9073
rect 2712 9074 2973 9075
rect 2880 9076 3021 9077
rect 2882 9078 3002 9079
rect 2885 9080 2987 9081
rect 2888 9082 2996 9083
rect 2894 9084 2899 9085
rect 1836 9086 2898 9087
rect 1437 9088 1838 9089
rect 2907 9088 3015 9089
rect 2910 9090 3018 9091
rect 2913 9092 3024 9093
rect 2916 9094 3028 9095
rect 2154 9096 2917 9097
rect 2155 9098 2173 9099
rect 2173 9100 2383 9101
rect 2383 9102 2407 9103
rect 2407 9104 2425 9105
rect 1590 9106 2426 9107
rect 2928 9106 3042 9107
rect 1986 9108 2928 9109
rect 1987 9110 2641 9111
rect 2641 9112 2707 9113
rect 2707 9114 2779 9115
rect 2931 9114 3069 9115
rect 2587 9116 2931 9117
rect 2934 9116 2947 9117
rect 2874 9118 2935 9119
rect 2940 9118 3048 9119
rect 2952 9120 3060 9121
rect 2955 9122 3063 9123
rect 2965 9124 2999 9125
rect 2983 9126 3005 9127
rect 1426 9135 1958 9136
rect 1426 9137 2264 9138
rect 1430 9139 1784 9140
rect 1430 9141 2186 9142
rect 1437 9143 2261 9144
rect 1440 9145 1814 9146
rect 1444 9147 2522 9148
rect 1444 9149 2258 9150
rect 1451 9151 2618 9152
rect 1458 9153 2594 9154
rect 1458 9155 2210 9156
rect 1461 9157 2306 9158
rect 1461 9159 1796 9160
rect 1470 9161 1535 9162
rect 1470 9163 2060 9164
rect 1473 9165 2342 9166
rect 1473 9167 2042 9168
rect 1531 9169 1892 9170
rect 1531 9171 2126 9172
rect 1534 9173 1574 9174
rect 1537 9175 1562 9176
rect 1543 9177 1556 9178
rect 1543 9179 1568 9180
rect 1549 9181 1874 9182
rect 1552 9183 1598 9184
rect 1564 9185 1700 9186
rect 1576 9187 2856 9188
rect 1585 9189 2549 9190
rect 1588 9191 2333 9192
rect 1603 9193 1658 9194
rect 1609 9195 1634 9196
rect 1609 9197 1664 9198
rect 1437 9199 1664 9200
rect 1615 9201 1646 9202
rect 1621 9203 1859 9204
rect 1621 9205 1676 9206
rect 1627 9207 2522 9208
rect 1627 9209 1682 9210
rect 1639 9211 1694 9212
rect 1645 9213 1688 9214
rect 1657 9215 1718 9216
rect 1675 9217 1766 9218
rect 1681 9219 1724 9220
rect 1687 9221 1742 9222
rect 1693 9223 1712 9224
rect 1423 9225 1712 9226
rect 1423 9227 2294 9228
rect 1717 9229 2006 9230
rect 1723 9231 2012 9232
rect 1726 9233 2015 9234
rect 1741 9235 2000 9236
rect 1747 9237 2258 9238
rect 1747 9239 2054 9240
rect 1765 9241 2066 9242
rect 1777 9243 2210 9244
rect 1777 9245 2138 9246
rect 1783 9247 1916 9248
rect 1795 9249 2168 9250
rect 1798 9251 2267 9252
rect 1813 9253 2192 9254
rect 1825 9255 2342 9256
rect 1825 9257 2090 9258
rect 1846 9259 2255 9260
rect 1852 9261 2189 9262
rect 1873 9263 2312 9264
rect 1885 9265 2336 9266
rect 1888 9267 2345 9268
rect 1894 9269 2387 9270
rect 1903 9271 2898 9272
rect 1524 9273 1904 9274
rect 1440 9275 1525 9276
rect 1915 9275 2372 9276
rect 1927 9277 2931 9278
rect 1927 9279 2384 9280
rect 1933 9281 2928 9282
rect 1933 9283 2234 9284
rect 1957 9285 2408 9286
rect 1999 9287 2348 9288
rect 2005 9289 2438 9290
rect 1735 9291 2438 9292
rect 1735 9293 2018 9294
rect 2011 9295 2300 9296
rect 2017 9297 2432 9298
rect 2023 9299 2192 9300
rect 1433 9301 2024 9302
rect 2032 9301 2417 9302
rect 2041 9303 2462 9304
rect 2053 9305 2676 9306
rect 2059 9307 2114 9308
rect 2029 9309 2114 9310
rect 2029 9311 2390 9312
rect 1849 9313 2390 9314
rect 1849 9315 2962 9316
rect 2065 9317 2450 9318
rect 1897 9319 2450 9320
rect 1897 9321 2324 9322
rect 1819 9323 2324 9324
rect 1819 9325 2198 9326
rect 1789 9327 2198 9328
rect 1789 9329 2048 9330
rect 2083 9329 2735 9330
rect 2083 9331 2492 9332
rect 2089 9333 2498 9334
rect 2098 9335 2456 9336
rect 2101 9337 2917 9338
rect 1969 9339 2102 9340
rect 1969 9341 2120 9342
rect 2119 9343 2528 9344
rect 2125 9345 2510 9346
rect 2131 9347 2914 9348
rect 2095 9349 2132 9350
rect 2095 9351 2504 9352
rect 2137 9353 2546 9354
rect 1651 9355 2546 9356
rect 1651 9357 1670 9358
rect 1669 9359 1760 9360
rect 1759 9361 2072 9362
rect 2071 9363 2444 9364
rect 1573 9365 2444 9366
rect 2143 9367 2627 9368
rect 2143 9369 2474 9370
rect 2149 9371 2921 9372
rect 2107 9373 2150 9374
rect 1939 9375 2108 9376
rect 1939 9377 2228 9378
rect 1945 9379 2228 9380
rect 1945 9381 2330 9382
rect 1951 9383 2330 9384
rect 1951 9385 2180 9386
rect 1993 9387 2180 9388
rect 1993 9389 2396 9390
rect 1843 9391 2396 9392
rect 1843 9393 2252 9394
rect 1771 9395 2252 9396
rect 1454 9397 1772 9398
rect 1454 9399 1501 9400
rect 1451 9401 1501 9402
rect 2161 9401 2779 9402
rect 1921 9403 2162 9404
rect 1921 9405 2240 9406
rect 1561 9407 2240 9408
rect 2164 9409 2315 9410
rect 2167 9411 2516 9412
rect 2173 9413 2186 9414
rect 1837 9415 2174 9416
rect 1837 9417 2246 9418
rect 2200 9419 2309 9420
rect 2212 9421 2327 9422
rect 2215 9423 2902 9424
rect 1855 9425 2216 9426
rect 2233 9425 2270 9426
rect 2155 9427 2270 9428
rect 2155 9429 2426 9430
rect 2245 9431 2534 9432
rect 2293 9433 2564 9434
rect 2299 9435 2570 9436
rect 2305 9437 2576 9438
rect 2311 9439 2716 9440
rect 2317 9441 2895 9442
rect 1801 9443 2318 9444
rect 1433 9445 1802 9446
rect 2335 9445 2582 9446
rect 2347 9447 2612 9448
rect 2356 9449 2471 9450
rect 2359 9451 2669 9452
rect 1831 9453 2360 9454
rect 1831 9455 2222 9456
rect 1753 9457 2222 9458
rect 1753 9459 2078 9460
rect 1527 9461 2078 9462
rect 1527 9463 2786 9464
rect 2371 9465 2588 9466
rect 2383 9467 2537 9468
rect 2407 9469 2636 9470
rect 2419 9471 2712 9472
rect 2419 9473 2624 9474
rect 2425 9475 2642 9476
rect 2431 9477 2905 9478
rect 2455 9479 2660 9480
rect 2461 9481 2849 9482
rect 2467 9483 2973 9484
rect 1705 9485 2468 9486
rect 1705 9487 1868 9488
rect 1867 9489 2288 9490
rect 2473 9489 2696 9490
rect 2476 9491 2699 9492
rect 2485 9493 2742 9494
rect 2485 9495 2672 9496
rect 2497 9497 2720 9498
rect 1963 9499 2719 9500
rect 1963 9501 2282 9502
rect 1981 9503 2282 9504
rect 1447 9505 1982 9506
rect 1447 9507 1856 9508
rect 2500 9507 2723 9508
rect 2515 9509 2702 9510
rect 2518 9511 2705 9512
rect 2527 9513 2732 9514
rect 2263 9515 2731 9516
rect 2533 9517 2966 9518
rect 2539 9519 2853 9520
rect 1729 9521 2540 9522
rect 1729 9523 1862 9524
rect 1861 9525 2036 9526
rect 2035 9527 2378 9528
rect 1909 9529 2378 9530
rect 1909 9531 2354 9532
rect 1879 9533 2354 9534
rect 1879 9535 2204 9536
rect 2551 9535 2673 9536
rect 2551 9537 2752 9538
rect 2557 9539 2728 9540
rect 2563 9541 2762 9542
rect 2566 9543 2765 9544
rect 2569 9545 2750 9546
rect 2575 9547 2768 9548
rect 2581 9549 2774 9550
rect 2593 9551 2744 9552
rect 2479 9553 2745 9554
rect 2479 9555 2678 9556
rect 2599 9557 2708 9558
rect 2401 9559 2709 9560
rect 2401 9561 2630 9562
rect 2605 9563 2749 9564
rect 2605 9565 2726 9566
rect 2611 9567 2801 9568
rect 2614 9569 2684 9570
rect 2620 9571 2798 9572
rect 2635 9573 2816 9574
rect 2638 9575 2819 9576
rect 2641 9577 2822 9578
rect 2647 9579 2828 9580
rect 2653 9581 2938 9582
rect 2653 9583 2834 9584
rect 2656 9585 2935 9586
rect 2656 9587 2837 9588
rect 2659 9589 2840 9590
rect 2665 9591 2846 9592
rect 2365 9593 2666 9594
rect 2678 9593 2871 9594
rect 2696 9595 2883 9596
rect 2699 9597 2886 9598
rect 2702 9599 2889 9600
rect 2705 9601 2892 9602
rect 2721 9603 2908 9604
rect 2724 9605 2911 9606
rect 2737 9607 2969 9608
rect 1987 9609 2738 9610
rect 1987 9611 2276 9612
rect 1807 9613 2276 9614
rect 1807 9615 1976 9616
rect 1975 9617 2414 9618
rect 2413 9619 2624 9620
rect 2754 9619 2941 9620
rect 2760 9621 2956 9622
rect 2772 9623 2959 9624
rect 2775 9625 2953 9626
rect 2781 9627 2976 9628
rect 2858 9629 2924 9630
rect 1423 9638 1519 9639
rect 1423 9640 1616 9641
rect 1426 9642 1832 9643
rect 1426 9644 2264 9645
rect 1430 9646 1778 9647
rect 1430 9648 2060 9649
rect 1433 9650 2528 9651
rect 1433 9652 2276 9653
rect 1437 9654 1604 9655
rect 1437 9656 1634 9657
rect 1440 9658 1603 9659
rect 1440 9660 2700 9661
rect 1444 9662 1712 9663
rect 1444 9664 2213 9665
rect 1447 9666 1699 9667
rect 1447 9668 1610 9669
rect 1451 9670 1900 9671
rect 1454 9672 2165 9673
rect 1456 9674 1880 9675
rect 1458 9676 1538 9677
rect 1459 9678 2099 9679
rect 1463 9680 1640 9681
rect 1466 9682 1646 9683
rect 1473 9684 1862 9685
rect 1481 9686 1495 9687
rect 1487 9688 1501 9689
rect 1493 9690 1513 9691
rect 1496 9692 1507 9693
rect 1499 9694 1544 9695
rect 1511 9696 2387 9697
rect 1518 9698 2414 9699
rect 1524 9700 2546 9701
rect 1527 9702 1633 9703
rect 1566 9704 1628 9705
rect 1573 9706 2450 9707
rect 1572 9708 1627 9709
rect 1578 9710 1652 9711
rect 1590 9712 1658 9713
rect 1521 9714 1657 9715
rect 1596 9716 1682 9717
rect 1611 9718 2066 9719
rect 1614 9720 1670 9721
rect 1638 9722 1688 9723
rect 1644 9724 1772 9725
rect 1650 9726 2198 9727
rect 1663 9728 2666 9729
rect 1662 9730 1730 9731
rect 1668 9732 1706 9733
rect 1680 9734 1784 9735
rect 1686 9736 2162 9737
rect 1693 9738 2634 9739
rect 1692 9740 2108 9741
rect 1704 9742 1802 9743
rect 1710 9744 2174 9745
rect 1726 9746 1744 9747
rect 1728 9748 2719 9749
rect 1753 9750 1777 9751
rect 1747 9752 1753 9753
rect 1741 9754 1747 9755
rect 1723 9756 1741 9757
rect 1722 9758 1808 9759
rect 1759 9760 1771 9761
rect 1735 9762 1759 9763
rect 1717 9764 1735 9765
rect 1716 9766 2102 9767
rect 1798 9768 1828 9769
rect 1800 9770 2180 9771
rect 1806 9772 2078 9773
rect 1830 9774 1970 9775
rect 1843 9776 1861 9777
rect 1819 9778 1843 9779
rect 1461 9780 1819 9781
rect 1846 9780 1864 9781
rect 1858 9782 1870 9783
rect 1867 9784 1879 9785
rect 1855 9786 1867 9787
rect 1837 9788 1855 9789
rect 1836 9790 2054 9791
rect 1888 9792 1924 9793
rect 1852 9794 1888 9795
rect 1851 9796 2201 9797
rect 1921 9798 2617 9799
rect 1885 9800 1921 9801
rect 1849 9802 1885 9803
rect 1813 9804 1849 9805
rect 1812 9806 1826 9807
rect 1795 9808 1825 9809
rect 1789 9810 1795 9811
rect 1470 9812 1789 9813
rect 1968 9812 2114 9813
rect 1981 9814 2709 9815
rect 1980 9816 2012 9817
rect 1987 9818 2053 9819
rect 1957 9820 1987 9821
rect 1927 9822 1957 9823
rect 1903 9824 1927 9825
rect 1902 9826 2024 9827
rect 1993 9828 2011 9829
rect 1992 9830 2712 9831
rect 2005 9832 2023 9833
rect 1951 9834 2005 9835
rect 1915 9836 1951 9837
rect 1897 9838 1915 9839
rect 1873 9840 1897 9841
rect 1531 9842 1873 9843
rect 2029 9842 2047 9843
rect 2035 9844 2059 9845
rect 2041 9846 2110 9847
rect 2017 9848 2041 9849
rect 1999 9850 2017 9851
rect 1975 9852 1999 9853
rect 1963 9854 1975 9855
rect 1945 9856 1963 9857
rect 1939 9858 1945 9859
rect 1909 9860 1939 9861
rect 1891 9862 1909 9863
rect 1534 9864 1891 9865
rect 2071 9864 2113 9865
rect 2070 9866 2192 9867
rect 2073 9868 2210 9869
rect 2076 9870 2132 9871
rect 2083 9872 2620 9873
rect 2082 9874 2669 9875
rect 2095 9876 2107 9877
rect 2089 9878 2095 9879
rect 2088 9880 2150 9881
rect 2100 9882 2673 9883
rect 2125 9884 2752 9885
rect 2124 9886 2216 9887
rect 2130 9888 2252 9889
rect 2133 9890 2417 9891
rect 2148 9892 2240 9893
rect 2155 9894 2742 9895
rect 2137 9896 2155 9897
rect 2119 9898 2137 9899
rect 2118 9900 2651 9901
rect 2160 9902 2186 9903
rect 1564 9904 2185 9905
rect 2167 9906 2173 9907
rect 1561 9908 2167 9909
rect 1560 9910 1622 9911
rect 1620 9912 1676 9913
rect 1608 9914 1675 9915
rect 2178 9914 2228 9915
rect 2190 9916 2318 9917
rect 2196 9918 2234 9919
rect 2202 9920 2246 9921
rect 2208 9922 2324 9923
rect 2214 9924 2282 9925
rect 2221 9926 2624 9927
rect 2034 9928 2624 9929
rect 2220 9930 2342 9931
rect 2226 9932 2294 9933
rect 2232 9934 2306 9935
rect 2238 9936 2631 9937
rect 2250 9938 2336 9939
rect 2257 9940 2782 9941
rect 2256 9942 2360 9943
rect 1514 9944 2359 9945
rect 2262 9946 2438 9947
rect 2269 9948 2728 9949
rect 2268 9950 2348 9951
rect 2274 9952 2608 9953
rect 2280 9954 2372 9955
rect 2286 9956 2396 9957
rect 2299 9958 2554 9959
rect 2298 9960 2384 9961
rect 2301 9962 2354 9963
rect 2304 9964 2378 9965
rect 2311 9966 2627 9967
rect 2310 9968 2444 9969
rect 2316 9970 2426 9971
rect 2322 9972 2420 9973
rect 2329 9974 2735 9975
rect 1576 9976 2329 9977
rect 1575 9978 2432 9979
rect 2334 9980 2402 9981
rect 2346 9982 2456 9983
rect 2352 9984 2462 9985
rect 2364 9986 2480 9987
rect 2370 9988 2486 9989
rect 2382 9990 2474 9991
rect 2385 9992 2477 9993
rect 2394 9994 2498 9995
rect 2397 9996 2408 9997
rect 2400 9998 2584 9999
rect 2412 10000 2534 10001
rect 2418 10002 2516 10003
rect 2421 10004 2519 10005
rect 2424 10006 2468 10007
rect 2427 10008 2471 10009
rect 2430 10010 2552 10011
rect 2028 10012 2551 10013
rect 2442 10014 2564 10015
rect 2445 10016 2567 10017
rect 2454 10018 2549 10019
rect 2457 10020 2540 10021
rect 2460 10022 2570 10023
rect 2466 10024 2576 10025
rect 2472 10026 2738 10027
rect 2478 10028 2582 10029
rect 2490 10030 2594 10031
rect 2496 10032 2600 10033
rect 2500 10034 2644 10035
rect 2502 10036 2569 10037
rect 2508 10038 2572 10039
rect 2526 10040 2612 10041
rect 2529 10042 2615 10043
rect 2532 10044 2636 10045
rect 2535 10046 2639 10047
rect 2544 10048 2648 10049
rect 2521 10050 2647 10051
rect 2556 10052 2657 10053
rect 2559 10054 2606 10055
rect 2389 10056 2605 10057
rect 2388 10058 2581 10059
rect 2574 10060 2660 10061
rect 2592 10062 2697 10063
rect 2595 10064 2679 10065
rect 2598 10066 2725 10067
rect 2601 10068 2779 10069
rect 2610 10070 2703 10071
rect 2613 10072 2706 10073
rect 2626 10074 2684 10075
rect 2637 10076 2642 10077
rect 2538 10078 2641 10079
rect 2656 10078 2755 10079
rect 2662 10080 2761 10081
rect 2668 10082 2776 10083
rect 2675 10084 2716 10085
rect 2680 10086 2773 10087
rect 2721 10088 2745 10089
rect 2730 10090 2749 10091
rect 1423 10099 1879 10100
rect 1426 10101 1645 10102
rect 1430 10103 2131 10104
rect 1429 10105 1789 10106
rect 1433 10107 1999 10108
rect 1432 10109 1603 10110
rect 1437 10111 1597 10112
rect 1436 10113 1744 10114
rect 1440 10115 1591 10116
rect 1439 10117 1561 10118
rect 1447 10119 1795 10120
rect 1446 10121 1900 10122
rect 1459 10123 2389 10124
rect 1463 10125 2455 10126
rect 1462 10127 1627 10128
rect 1466 10129 2329 10130
rect 1465 10131 1675 10132
rect 1481 10133 2031 10134
rect 1480 10135 1500 10136
rect 1487 10137 2043 10138
rect 1486 10139 1975 10140
rect 1489 10141 1957 10142
rect 1493 10143 2067 10144
rect 1496 10145 1924 10146
rect 1498 10147 2299 10148
rect 1501 10149 2353 10150
rect 1505 10151 1927 10152
rect 1508 10153 2163 10154
rect 1511 10155 1801 10156
rect 1514 10157 2071 10158
rect 1518 10159 1596 10160
rect 1521 10161 1888 10162
rect 1523 10163 1612 10164
rect 1535 10165 1579 10166
rect 1541 10167 1555 10168
rect 1553 10169 2527 10170
rect 1556 10171 2199 10172
rect 1566 10173 1578 10174
rect 1568 10175 2137 10176
rect 1572 10177 2359 10178
rect 1458 10179 1572 10180
rect 1575 10179 2425 10180
rect 1583 10181 1729 10182
rect 1589 10183 2263 10184
rect 1601 10185 1657 10186
rect 1620 10187 1644 10188
rect 1619 10189 1639 10190
rect 1614 10191 1638 10192
rect 1613 10193 1633 10194
rect 1650 10193 1656 10194
rect 1649 10195 2257 10196
rect 1664 10197 2191 10198
rect 1673 10199 2209 10200
rect 1680 10201 2388 10202
rect 1679 10203 2221 10204
rect 1686 10205 1728 10206
rect 1722 10207 1782 10208
rect 1721 10209 2125 10210
rect 1734 10211 1809 10212
rect 1733 10213 2167 10214
rect 1787 10215 2275 10216
rect 1793 10217 2347 10218
rect 1827 10219 1941 10220
rect 1832 10221 2371 10222
rect 1836 10223 1878 10224
rect 1764 10225 1836 10226
rect 1698 10227 1764 10228
rect 1697 10229 2185 10230
rect 1848 10231 1956 10232
rect 1776 10233 1848 10234
rect 1716 10235 1776 10236
rect 1668 10237 1716 10238
rect 1851 10237 1959 10238
rect 1854 10239 1974 10240
rect 1853 10241 2179 10242
rect 1863 10243 1983 10244
rect 1869 10245 2013 10246
rect 1920 10247 2064 10248
rect 1925 10249 2197 10250
rect 1932 10251 2620 10252
rect 1931 10253 2029 10254
rect 1884 10255 2028 10256
rect 1883 10257 1903 10258
rect 1901 10259 2077 10260
rect 1938 10261 2076 10262
rect 1824 10263 1938 10264
rect 1752 10265 1824 10266
rect 1444 10267 1752 10268
rect 1443 10269 2089 10270
rect 1950 10271 2223 10272
rect 1872 10273 1950 10274
rect 1812 10275 1872 10276
rect 1746 10277 1812 10278
rect 1704 10279 1746 10280
rect 1703 10281 2149 10282
rect 1952 10283 2134 10284
rect 1997 10285 2053 10286
rect 1914 10287 2052 10288
rect 1818 10289 1914 10290
rect 1758 10291 1818 10292
rect 1757 10293 2319 10294
rect 2016 10295 2088 10296
rect 1908 10297 2016 10298
rect 1907 10299 2551 10300
rect 2024 10301 2530 10302
rect 2034 10303 2136 10304
rect 2033 10305 2203 10306
rect 2040 10307 2627 10308
rect 1896 10309 2040 10310
rect 1895 10311 2317 10312
rect 2046 10313 2205 10314
rect 1608 10315 2046 10316
rect 1565 10317 1608 10318
rect 2054 10317 2074 10318
rect 2058 10319 2617 10320
rect 1962 10321 2058 10322
rect 1842 10323 1962 10324
rect 1770 10325 1842 10326
rect 1769 10327 2316 10328
rect 2060 10329 2311 10330
rect 2069 10331 2101 10332
rect 2078 10333 2428 10334
rect 2082 10335 2148 10336
rect 2081 10337 2113 10338
rect 2010 10339 2112 10340
rect 1456 10341 2010 10342
rect 1455 10343 1626 10344
rect 2094 10343 2166 10344
rect 2093 10345 2220 10346
rect 2106 10347 2651 10348
rect 1992 10349 2106 10350
rect 1991 10351 2624 10352
rect 2118 10353 2124 10354
rect 1986 10355 2118 10356
rect 1866 10357 1986 10358
rect 1806 10359 1866 10360
rect 1740 10361 1806 10362
rect 1692 10363 1740 10364
rect 1691 10365 1711 10366
rect 1662 10367 1710 10368
rect 2129 10367 2161 10368
rect 2154 10369 2187 10370
rect 2153 10371 2391 10372
rect 2159 10373 2215 10374
rect 2168 10375 2323 10376
rect 2172 10377 2631 10378
rect 2174 10379 2227 10380
rect 2180 10381 2233 10382
rect 2192 10383 2251 10384
rect 2201 10385 2401 10386
rect 2207 10387 2305 10388
rect 2225 10389 2269 10390
rect 2231 10391 2503 10392
rect 2238 10393 2425 10394
rect 2243 10395 2461 10396
rect 2249 10397 2383 10398
rect 2252 10399 2386 10400
rect 2255 10401 2435 10402
rect 2261 10403 2463 10404
rect 2267 10405 2413 10406
rect 2273 10407 2473 10408
rect 2286 10409 2608 10410
rect 2291 10411 2443 10412
rect 2294 10413 2446 10414
rect 2022 10415 2446 10416
rect 1980 10417 2022 10418
rect 1860 10419 1980 10420
rect 1859 10421 1969 10422
rect 1967 10423 2005 10424
rect 1944 10425 2004 10426
rect 1890 10427 1944 10428
rect 1830 10429 1890 10430
rect 2297 10429 2479 10430
rect 2301 10431 2554 10432
rect 2309 10433 2557 10434
rect 2312 10435 2509 10436
rect 2321 10437 2406 10438
rect 2334 10439 2453 10440
rect 2333 10441 2533 10442
rect 2336 10443 2536 10444
rect 2339 10445 2641 10446
rect 2345 10447 2409 10448
rect 2351 10449 2439 10450
rect 2357 10451 2442 10452
rect 2364 10453 2644 10454
rect 2369 10455 2575 10456
rect 2375 10457 2634 10458
rect 2381 10459 2599 10460
rect 2384 10461 2602 10462
rect 2394 10463 2647 10464
rect 2397 10465 2456 10466
rect 2399 10467 2593 10468
rect 2402 10469 2596 10470
rect 2411 10471 2611 10472
rect 2414 10473 2614 10474
rect 2418 10475 2584 10476
rect 2109 10477 2418 10478
rect 2421 10477 2581 10478
rect 2280 10479 2421 10480
rect 2279 10481 2431 10482
rect 2427 10483 2539 10484
rect 2431 10485 2467 10486
rect 2448 10487 2605 10488
rect 2457 10489 2569 10490
rect 2459 10491 2497 10492
rect 2465 10493 2657 10494
rect 2471 10495 2663 10496
rect 2477 10497 2669 10498
rect 2490 10499 2654 10500
rect 2489 10501 2681 10502
rect 2492 10503 2684 10504
rect 2544 10505 2638 10506
rect 2559 10507 2572 10508
rect 1429 10516 1536 10517
rect 1432 10518 2028 10519
rect 1436 10520 1770 10521
rect 1439 10522 1665 10523
rect 1441 10524 1650 10525
rect 1443 10526 2010 10527
rect 1444 10528 1481 10529
rect 1448 10530 1734 10531
rect 1451 10532 1782 10533
rect 1455 10534 1620 10535
rect 1455 10536 1746 10537
rect 1458 10538 1614 10539
rect 1465 10540 1692 10541
rect 1467 10542 1535 10543
rect 1470 10544 2031 10545
rect 1479 10546 1884 10547
rect 1482 10548 1820 10549
rect 1486 10550 2412 10551
rect 1486 10552 1959 10553
rect 1489 10554 1890 10555
rect 1489 10556 1566 10557
rect 1498 10558 2016 10559
rect 1498 10560 1953 10561
rect 1505 10562 1986 10563
rect 1504 10564 1542 10565
rect 1510 10566 1634 10567
rect 1523 10568 1529 10569
rect 1462 10570 1523 10571
rect 1537 10570 1964 10571
rect 1553 10572 1902 10573
rect 1552 10574 2435 10575
rect 1556 10576 2181 10577
rect 1558 10578 2046 10579
rect 1561 10580 1758 10581
rect 1568 10582 2346 10583
rect 1577 10584 1778 10585
rect 1576 10586 1833 10587
rect 1612 10588 1638 10589
rect 1618 10590 1644 10591
rect 1630 10592 2022 10593
rect 1651 10594 1674 10595
rect 1655 10596 2220 10597
rect 1654 10598 2232 10599
rect 1660 10600 1794 10601
rect 1666 10602 2316 10603
rect 1672 10604 1710 10605
rect 1684 10606 1704 10607
rect 1446 10608 1703 10609
rect 1690 10610 1752 10611
rect 1708 10612 1764 10613
rect 1727 10614 2391 10615
rect 1697 10616 1727 10617
rect 1732 10616 1776 10617
rect 1735 10618 2043 10619
rect 1750 10620 1806 10621
rect 1753 10622 1809 10623
rect 1756 10624 1812 10625
rect 1762 10626 1818 10627
rect 1774 10628 1824 10629
rect 1780 10630 2202 10631
rect 1789 10632 1842 10633
rect 1795 10634 1848 10635
rect 1801 10636 1854 10637
rect 1807 10638 1866 10639
rect 1813 10640 1878 10641
rect 1831 10642 2169 10643
rect 1835 10644 1889 10645
rect 1843 10646 1926 10647
rect 1849 10648 1938 10649
rect 1852 10650 1941 10651
rect 1855 10652 1914 10653
rect 1859 10654 2177 10655
rect 1861 10656 1992 10657
rect 1867 10658 2034 10659
rect 1871 10660 2102 10661
rect 1873 10662 1962 10663
rect 1876 10664 2013 10665
rect 1879 10666 1974 10667
rect 1885 10668 1980 10669
rect 1891 10670 1956 10671
rect 1895 10672 2132 10673
rect 1739 10674 1895 10675
rect 1738 10676 1788 10677
rect 1897 10676 2160 10677
rect 1903 10678 1944 10679
rect 1907 10680 2425 10681
rect 1458 10682 1907 10683
rect 1909 10682 2004 10683
rect 1915 10684 1932 10685
rect 1921 10686 1968 10687
rect 1924 10688 2025 10689
rect 1927 10690 2052 10691
rect 1930 10692 2055 10693
rect 1936 10694 2313 10695
rect 1939 10696 2064 10697
rect 1942 10698 2067 10699
rect 1945 10700 2058 10701
rect 1501 10702 2057 10703
rect 1949 10704 2197 10705
rect 1679 10706 1949 10707
rect 1678 10708 1716 10709
rect 1508 10710 1715 10711
rect 1951 10710 2076 10711
rect 1954 10712 2079 10713
rect 1957 10714 2180 10715
rect 1969 10716 2094 10717
rect 1972 10718 2310 10719
rect 1975 10720 2082 10721
rect 1982 10722 2456 10723
rect 1981 10724 2124 10725
rect 1987 10726 2070 10727
rect 1993 10728 2118 10729
rect 1997 10730 2099 10731
rect 1999 10732 2112 10733
rect 2002 10734 2163 10735
rect 2005 10736 2428 10737
rect 2011 10738 2136 10739
rect 2017 10740 2148 10741
rect 2029 10742 2142 10743
rect 2039 10744 2141 10745
rect 2041 10746 2193 10747
rect 2047 10748 2199 10749
rect 2060 10750 2421 10751
rect 2062 10752 2208 10753
rect 2068 10754 2253 10755
rect 2071 10756 2187 10757
rect 1601 10758 2187 10759
rect 1600 10760 1626 10761
rect 1607 10762 1625 10763
rect 1595 10764 1607 10765
rect 1589 10766 1595 10767
rect 1583 10768 1589 10769
rect 1571 10770 1583 10771
rect 2074 10770 2274 10771
rect 2080 10772 2453 10773
rect 2083 10774 2166 10775
rect 2087 10776 2449 10777
rect 2086 10778 2244 10779
rect 2092 10780 2415 10781
rect 2095 10782 2298 10783
rect 2105 10784 2144 10785
rect 2110 10786 2280 10787
rect 2122 10788 2292 10789
rect 2125 10790 2295 10791
rect 2129 10792 2203 10793
rect 2128 10794 2334 10795
rect 2134 10796 2340 10797
rect 2146 10798 2352 10799
rect 2153 10800 2191 10801
rect 2158 10802 2400 10803
rect 2161 10804 2322 10805
rect 2164 10806 2337 10807
rect 2167 10808 2194 10809
rect 2170 10810 2382 10811
rect 2174 10812 2200 10813
rect 2173 10814 2358 10815
rect 2183 10816 2403 10817
rect 2204 10818 2388 10819
rect 2205 10820 2439 10821
rect 2208 10822 2466 10823
rect 2220 10824 2490 10825
rect 2222 10826 2250 10827
rect 2223 10828 2493 10829
rect 2225 10830 2463 10831
rect 2226 10832 2472 10833
rect 2229 10834 2478 10835
rect 2255 10836 2418 10837
rect 2261 10838 2432 10839
rect 2267 10840 2460 10841
rect 2318 10842 2446 10843
rect 2369 10844 2406 10845
rect 2375 10846 2409 10847
rect 2384 10848 2442 10849
rect 1423 10857 1715 10858
rect 1426 10859 1601 10860
rect 1430 10861 1874 10862
rect 1433 10863 1922 10864
rect 1437 10865 1796 10866
rect 1441 10867 1607 10868
rect 1440 10869 1754 10870
rect 1444 10871 1683 10872
rect 1444 10873 1529 10874
rect 1451 10875 1733 10876
rect 1450 10877 1904 10878
rect 1453 10879 2030 10880
rect 1458 10881 1895 10882
rect 1448 10883 1460 10884
rect 1447 10885 1523 10886
rect 1462 10887 1685 10888
rect 1467 10889 1652 10890
rect 1470 10891 1949 10892
rect 1477 10893 2102 10894
rect 1479 10895 1814 10896
rect 1482 10897 1808 10898
rect 1486 10899 1721 10900
rect 1489 10901 1778 10902
rect 1489 10903 1928 10904
rect 1496 10905 1511 10906
rect 1498 10907 1509 10908
rect 1499 10909 1505 10910
rect 1511 10909 1907 10910
rect 1514 10911 1553 10912
rect 1520 10913 1589 10914
rect 1526 10915 1595 10916
rect 1532 10917 1613 10918
rect 1537 10919 1952 10920
rect 1538 10921 1619 10922
rect 1544 10923 1625 10924
rect 1550 10925 1583 10926
rect 1558 10927 1925 10928
rect 1561 10929 1767 10930
rect 1568 10931 1661 10932
rect 1586 10933 1673 10934
rect 1592 10935 1679 10936
rect 1595 10937 1877 10938
rect 1598 10939 1709 10940
rect 1604 10941 1866 10942
rect 1622 10943 1751 10944
rect 1625 10945 1757 10946
rect 1630 10947 2162 10948
rect 1631 10949 1763 10950
rect 1576 10951 1764 10952
rect 1577 10953 1955 10954
rect 1633 10955 2042 10956
rect 1534 10957 1635 10958
rect 1637 10957 1691 10958
rect 1643 10959 1703 10960
rect 1661 10961 1739 10962
rect 1673 10963 1781 10964
rect 1455 10965 1782 10966
rect 1456 10967 1736 10968
rect 1676 10969 2144 10970
rect 1688 10971 1832 10972
rect 1694 10973 1850 10974
rect 1697 10975 1853 10976
rect 1712 10977 1892 10978
rect 1715 10979 1856 10980
rect 1724 10981 1880 10982
rect 1726 10983 1951 10984
rect 1730 10985 1886 10986
rect 1733 10987 1889 10988
rect 1736 10989 1898 10990
rect 1742 10991 1844 10992
rect 1748 10993 1910 10994
rect 1654 10995 1911 10996
rect 1655 10997 1790 10998
rect 1754 10999 1868 11000
rect 1760 11001 1916 11002
rect 1769 11003 1940 11004
rect 1666 11005 1940 11006
rect 1772 11007 1943 11008
rect 1774 11009 2180 11010
rect 1492 11011 1776 11012
rect 1778 11011 1931 11012
rect 1787 11013 1921 11014
rect 1790 11015 2003 11016
rect 1793 11017 1964 11018
rect 1799 11019 1970 11020
rect 1801 11021 1954 11022
rect 1805 11023 2184 11024
rect 1811 11025 1976 11026
rect 1817 11027 1982 11028
rect 1819 11029 2141 11030
rect 1823 11031 1988 11032
rect 1829 11033 2012 11034
rect 1835 11035 2006 11036
rect 1841 11037 2200 11038
rect 1847 11039 2057 11040
rect 1859 11041 2048 11042
rect 1861 11043 1914 11044
rect 1574 11045 1863 11046
rect 1868 11045 2072 11046
rect 1877 11047 2093 11048
rect 1880 11049 2096 11050
rect 1883 11051 1973 11052
rect 1886 11053 1937 11054
rect 1889 11055 2129 11056
rect 1892 11057 2132 11058
rect 1895 11059 2123 11060
rect 1904 11061 2159 11062
rect 1907 11063 2168 11064
rect 1917 11065 1958 11066
rect 1923 11067 2171 11068
rect 1926 11069 2147 11070
rect 1929 11071 2087 11072
rect 1932 11073 2075 11074
rect 1936 11075 1946 11076
rect 1853 11077 1947 11078
rect 1943 11079 2063 11080
rect 1956 11081 2111 11082
rect 1959 11083 2126 11084
rect 1993 11085 2177 11086
rect 1999 11087 2187 11088
rect 2017 11089 2194 11090
rect 2068 11091 2099 11092
rect 2080 11093 2206 11094
rect 2083 11095 2197 11096
rect 2134 11097 2203 11098
rect 2164 11099 2209 11100
rect 2173 11101 2191 11102
rect 2220 11101 2230 11102
rect 2223 11103 2227 11104
rect 1423 11112 1605 11113
rect 1426 11114 1599 11115
rect 1430 11116 1535 11117
rect 1429 11118 1632 11119
rect 1433 11120 1749 11121
rect 1432 11122 1764 11123
rect 1437 11124 1656 11125
rect 1436 11126 1773 11127
rect 1440 11128 1734 11129
rect 1439 11130 1539 11131
rect 1444 11132 1478 11133
rect 1443 11134 1533 11135
rect 1447 11136 1596 11137
rect 1446 11138 1593 11139
rect 1450 11140 1623 11141
rect 1450 11142 1716 11143
rect 1453 11144 1713 11145
rect 1453 11146 1788 11147
rect 1459 11148 1644 11149
rect 1462 11150 1638 11151
rect 1465 11152 1695 11153
rect 1468 11154 1626 11155
rect 1471 11156 1635 11157
rect 1474 11158 1587 11159
rect 1483 11160 1731 11161
rect 1486 11162 1725 11163
rect 1489 11164 1884 11165
rect 1489 11166 1698 11167
rect 1492 11168 1836 11169
rect 1492 11170 1918 11171
rect 1496 11172 1509 11173
rect 1495 11174 1779 11175
rect 1499 11176 1512 11177
rect 1498 11178 1770 11179
rect 1501 11180 1545 11181
rect 1504 11182 1527 11183
rect 1507 11184 1521 11185
rect 1514 11186 1520 11187
rect 1513 11188 1551 11189
rect 1525 11190 1761 11191
rect 1546 11192 1908 11193
rect 1555 11194 1830 11195
rect 1561 11196 1755 11197
rect 1564 11198 1791 11199
rect 1568 11200 1604 11201
rect 1574 11202 1586 11203
rect 1573 11204 1824 11205
rect 1577 11206 1589 11207
rect 1576 11208 1794 11209
rect 1579 11210 1887 11211
rect 1582 11212 1800 11213
rect 1597 11214 1893 11215
rect 1600 11216 1677 11217
rect 1606 11218 1806 11219
rect 1609 11220 1737 11221
rect 1612 11222 1662 11223
rect 1616 11224 1818 11225
rect 1619 11226 1812 11227
rect 1623 11228 1689 11229
rect 1626 11230 1683 11231
rect 1629 11232 1776 11233
rect 1632 11234 1869 11235
rect 1673 11236 1954 11237
rect 1742 11238 1914 11239
rect 1766 11240 1866 11241
rect 1781 11242 1947 11243
rect 1841 11244 1940 11245
rect 1847 11246 1944 11247
rect 1853 11248 1863 11249
rect 1859 11250 1951 11251
rect 1877 11252 1933 11253
rect 1880 11254 1930 11255
rect 1889 11256 1911 11257
rect 1895 11258 1957 11259
rect 1904 11260 1921 11261
rect 1923 11260 1960 11261
rect 1926 11262 1937 11263
rect 1429 11271 1469 11272
rect 1432 11273 1472 11274
rect 1436 11275 1484 11276
rect 1439 11277 1487 11278
rect 1443 11279 1457 11280
rect 1446 11281 1475 11282
rect 1450 11283 1556 11284
rect 1453 11285 1526 11286
rect 1465 11287 1630 11288
rect 1477 11289 1520 11290
rect 1480 11291 1535 11292
rect 1489 11293 1499 11294
rect 1489 11295 1586 11296
rect 1492 11297 1496 11298
rect 1492 11299 1589 11300
rect 1501 11301 1508 11302
rect 1504 11303 1514 11304
rect 1546 11303 1604 11304
rect 1561 11305 1633 11306
rect 1564 11307 1610 11308
rect 1573 11309 1620 11310
rect 1576 11311 1617 11312
rect 1579 11313 1613 11314
rect 1582 11315 1607 11316
rect 1597 11317 1627 11318
rect 1600 11319 1624 11320
rect 1477 11328 1493 11329
rect 1480 11330 1490 11331
<< metal2 >>
rect 1423 683 1424 733
rect 1561 683 1562 733
rect 1426 685 1427 733
rect 1594 685 1595 733
rect 1430 687 1431 733
rect 1437 687 1438 733
rect 1433 689 1434 733
rect 1449 689 1450 733
rect 1440 691 1441 733
rect 1458 691 1459 733
rect 1443 693 1444 733
rect 1486 693 1487 733
rect 1446 695 1447 733
rect 1489 695 1490 733
rect 1452 697 1453 733
rect 1597 697 1598 733
rect 1455 699 1456 733
rect 1492 699 1493 733
rect 1461 701 1462 733
rect 1498 701 1499 733
rect 1464 703 1465 733
rect 1567 703 1568 733
rect 1468 705 1469 733
rect 1516 705 1517 733
rect 1471 707 1472 733
rect 1555 707 1556 733
rect 1495 709 1496 733
rect 1629 709 1630 733
rect 1507 711 1508 733
rect 1519 711 1520 733
rect 1510 713 1511 733
rect 1513 713 1514 733
rect 1525 713 1526 733
rect 1600 713 1601 733
rect 1543 715 1544 733
rect 1606 715 1607 733
rect 1546 717 1547 733
rect 1549 717 1550 733
rect 1552 717 1553 733
rect 1618 717 1619 733
rect 1558 719 1559 733
rect 1636 719 1637 733
rect 1564 721 1565 733
rect 1632 721 1633 733
rect 1579 723 1580 733
rect 1639 723 1640 733
rect 1582 725 1583 733
rect 1622 725 1623 733
rect 1603 727 1604 733
rect 1609 727 1610 733
rect 1612 727 1613 733
rect 1625 727 1626 733
rect 1615 729 1616 733
rect 1642 729 1643 733
rect 1423 737 1424 740
rect 1682 739 1683 902
rect 1423 741 1424 902
rect 1685 741 1686 902
rect 1426 737 1427 744
rect 1721 743 1722 902
rect 1426 745 1427 902
rect 1724 745 1725 902
rect 1430 737 1431 748
rect 1709 747 1710 902
rect 1430 749 1431 902
rect 1679 749 1680 902
rect 1433 737 1434 752
rect 1649 751 1650 902
rect 1433 753 1434 902
rect 1667 753 1668 902
rect 1437 737 1438 756
rect 1589 755 1590 902
rect 1436 757 1437 902
rect 2029 757 2030 902
rect 1440 737 1441 760
rect 1688 759 1689 902
rect 1439 761 1440 902
rect 1805 761 1806 902
rect 1443 737 1444 764
rect 1715 763 1716 902
rect 1443 765 1444 902
rect 1706 765 1707 902
rect 1446 737 1447 768
rect 1922 767 1923 902
rect 1446 769 1447 902
rect 1634 769 1635 902
rect 1455 737 1456 772
rect 1961 771 1962 902
rect 1464 737 1465 774
rect 1895 773 1896 902
rect 1465 775 1466 902
rect 1661 775 1662 902
rect 1468 737 1469 778
rect 1733 777 1734 902
rect 1471 737 1472 780
rect 1781 779 1782 902
rect 1474 781 1475 902
rect 1964 781 1965 902
rect 1481 783 1482 902
rect 1541 783 1542 902
rect 1484 785 1485 902
rect 1535 785 1536 902
rect 1486 737 1487 788
rect 1703 787 1704 902
rect 1489 737 1490 790
rect 1697 789 1698 902
rect 1505 791 1506 902
rect 1597 737 1598 792
rect 1507 737 1508 794
rect 1817 793 1818 902
rect 1510 737 1511 796
rect 1745 795 1746 902
rect 1511 797 1512 902
rect 1513 737 1514 798
rect 1516 737 1517 798
rect 1727 797 1728 902
rect 1477 799 1478 902
rect 1517 799 1518 902
rect 1519 737 1520 800
rect 1793 799 1794 902
rect 1523 801 1524 902
rect 1582 737 1583 802
rect 1525 737 1526 804
rect 1763 803 1764 902
rect 1543 737 1544 806
rect 1999 805 2000 902
rect 1546 737 1547 808
rect 1832 807 1833 902
rect 1547 809 1548 902
rect 1889 809 1890 902
rect 1552 737 1553 812
rect 1877 811 1878 902
rect 1555 737 1556 814
rect 1751 813 1752 902
rect 1558 737 1559 816
rect 1928 815 1929 902
rect 1561 737 1562 818
rect 1955 817 1956 902
rect 1564 737 1565 820
rect 1757 819 1758 902
rect 1567 737 1568 822
rect 1835 821 1836 902
rect 1549 737 1550 824
rect 1568 823 1569 902
rect 1550 825 1551 902
rect 1739 825 1740 902
rect 1571 827 1572 902
rect 1639 737 1640 828
rect 1579 737 1580 830
rect 1841 829 1842 902
rect 1594 737 1595 832
rect 1820 831 1821 902
rect 1458 737 1459 834
rect 1595 833 1596 902
rect 1600 737 1601 834
rect 1958 833 1959 902
rect 1601 835 1602 902
rect 1603 737 1604 836
rect 1606 737 1607 836
rect 1907 835 1908 902
rect 1609 737 1610 838
rect 1910 837 1911 902
rect 1612 737 1613 840
rect 1937 839 1938 902
rect 1615 737 1616 842
rect 1916 841 1917 902
rect 1449 737 1450 844
rect 1616 843 1617 902
rect 1450 845 1451 902
rect 1610 845 1611 902
rect 1618 737 1619 846
rect 1986 845 1987 902
rect 1452 737 1453 848
rect 1619 847 1620 902
rect 1453 849 1454 902
rect 1604 849 1605 902
rect 1622 737 1623 850
rect 2012 849 2013 902
rect 1625 737 1626 852
rect 1799 851 1800 902
rect 1492 737 1493 854
rect 1625 853 1626 902
rect 1493 855 1494 902
rect 1952 855 1953 902
rect 1629 737 1630 858
rect 1691 857 1692 902
rect 1632 737 1633 860
rect 1769 859 1770 902
rect 1495 737 1496 862
rect 1631 861 1632 902
rect 1496 863 1497 902
rect 1829 863 1830 902
rect 1636 737 1637 866
rect 1736 865 1737 902
rect 1498 737 1499 868
rect 1637 867 1638 902
rect 1642 737 1643 868
rect 2009 867 2010 902
rect 1461 737 1462 870
rect 1643 869 1644 902
rect 1462 871 1463 902
rect 1931 871 1932 902
rect 1655 873 1656 902
rect 2032 873 2033 902
rect 1673 875 1674 902
rect 1996 875 1997 902
rect 1775 877 1776 902
rect 1967 877 1968 902
rect 1787 879 1788 902
rect 1971 879 1972 902
rect 1811 881 1812 902
rect 2015 881 2016 902
rect 1847 883 1848 902
rect 1992 883 1993 902
rect 1853 885 1854 902
rect 1989 885 1990 902
rect 1859 887 1860 902
rect 2022 887 2023 902
rect 1913 889 1914 902
rect 1919 889 1920 902
rect 1925 889 1926 902
rect 2036 889 2037 902
rect 1934 891 1935 902
rect 2039 891 2040 902
rect 1940 893 1941 902
rect 2018 893 2019 902
rect 1943 895 1944 902
rect 2006 895 2007 902
rect 1974 897 1975 902
rect 2025 897 2026 902
rect 1977 899 1978 902
rect 2003 899 2004 902
rect 1417 908 1418 1183
rect 1556 908 1557 1183
rect 1430 906 1431 911
rect 1643 906 1644 911
rect 1443 906 1444 913
rect 1901 912 1902 1183
rect 1448 914 1449 1183
rect 2288 914 2289 1183
rect 1450 906 1451 917
rect 2219 916 2220 1183
rect 1455 918 1456 1183
rect 1574 918 1575 1183
rect 1459 920 1460 1183
rect 1631 906 1632 921
rect 1474 906 1475 923
rect 1526 922 1527 1183
rect 1477 906 1478 925
rect 1511 906 1512 925
rect 1481 906 1482 927
rect 2063 926 2064 1183
rect 1484 906 1485 929
rect 2213 928 2214 1183
rect 1483 930 1484 1183
rect 1568 906 1569 931
rect 1486 932 1487 1183
rect 1943 906 1944 933
rect 1490 934 1491 1183
rect 1853 906 1854 935
rect 1493 906 1494 937
rect 2159 936 2160 1183
rect 1474 938 1475 1183
rect 1493 938 1494 1183
rect 1502 938 1503 1183
rect 2240 938 2241 1183
rect 1505 906 1506 941
rect 1514 940 1515 1183
rect 1505 942 1506 1183
rect 2237 942 2238 1183
rect 1517 906 1518 945
rect 1532 944 1533 1183
rect 1520 946 1521 1183
rect 1523 906 1524 947
rect 1535 906 1536 947
rect 2111 946 2112 1183
rect 1541 906 1542 949
rect 2129 948 2130 1183
rect 1547 906 1548 951
rect 1910 906 1911 951
rect 1550 906 1551 953
rect 2183 952 2184 1183
rect 1420 954 1421 1183
rect 1550 954 1551 1183
rect 1586 954 1587 1183
rect 1616 906 1617 955
rect 1592 956 1593 1183
rect 2276 956 2277 1183
rect 1601 906 1602 959
rect 1712 958 1713 1183
rect 1589 906 1590 961
rect 1601 960 1602 1183
rect 1496 906 1497 963
rect 1589 962 1590 1183
rect 1607 962 1608 1183
rect 1673 906 1674 963
rect 1613 964 1614 1183
rect 1679 906 1680 965
rect 1595 906 1596 967
rect 1679 966 1680 1183
rect 1595 968 1596 1183
rect 2282 968 2283 1183
rect 1619 906 1620 971
rect 1883 970 1884 1183
rect 1619 972 1620 1183
rect 1685 906 1686 973
rect 1439 906 1440 975
rect 1685 974 1686 1183
rect 1438 976 1439 1183
rect 1568 976 1569 1183
rect 1625 906 1626 977
rect 2345 976 2346 1183
rect 1625 978 1626 1183
rect 1703 906 1704 979
rect 1423 906 1424 981
rect 1703 980 1704 1183
rect 1424 982 1425 1183
rect 1979 982 1980 1183
rect 1631 984 1632 1183
rect 1721 906 1722 985
rect 1637 906 1638 987
rect 2048 986 2049 1183
rect 1471 988 1472 1183
rect 1637 988 1638 1183
rect 1643 988 1644 1183
rect 1697 906 1698 989
rect 1649 906 1650 991
rect 1673 990 1674 1183
rect 1649 992 1650 1183
rect 1667 906 1668 993
rect 1667 994 1668 1183
rect 2374 994 2375 1183
rect 1676 996 1677 1183
rect 1682 906 1683 997
rect 1691 906 1692 997
rect 1865 996 1866 1183
rect 1697 998 1698 1183
rect 1769 906 1770 999
rect 1709 906 1710 1001
rect 1871 1000 1872 1183
rect 1436 906 1437 1003
rect 1709 1002 1710 1183
rect 1721 1002 1722 1183
rect 1757 906 1758 1003
rect 1724 906 1725 1005
rect 2045 1004 2046 1183
rect 1739 906 1740 1007
rect 2177 1006 2178 1183
rect 1727 906 1728 1009
rect 1739 1008 1740 1183
rect 1727 1010 1728 1183
rect 2424 1010 2425 1183
rect 1745 906 1746 1013
rect 2093 1012 2094 1183
rect 1431 1014 1432 1183
rect 1745 1014 1746 1183
rect 1751 906 1752 1015
rect 1823 1014 1824 1183
rect 1733 906 1734 1017
rect 1751 1016 1752 1183
rect 1688 906 1689 1019
rect 1733 1018 1734 1183
rect 1757 1018 1758 1183
rect 1775 906 1776 1019
rect 1465 906 1466 1021
rect 1775 1020 1776 1183
rect 1769 1022 1770 1183
rect 2015 906 2016 1023
rect 1426 906 1427 1025
rect 2015 1024 2016 1183
rect 1427 1026 1428 1183
rect 1598 1026 1599 1183
rect 1781 906 1782 1027
rect 1853 1026 1854 1183
rect 1793 906 1794 1029
rect 2069 1028 2070 1183
rect 1793 1030 1794 1183
rect 2364 1030 2365 1183
rect 1817 906 1818 1033
rect 2087 1032 2088 1183
rect 1462 906 1463 1035
rect 1817 1034 1818 1183
rect 1462 1036 1463 1183
rect 2324 1036 2325 1183
rect 1820 906 1821 1039
rect 2216 1038 2217 1183
rect 1829 906 1830 1041
rect 2153 1040 2154 1183
rect 1763 906 1764 1043
rect 1829 1042 1830 1183
rect 1763 1044 1764 1183
rect 2371 1044 2372 1183
rect 1832 906 1833 1047
rect 2165 1046 2166 1183
rect 1835 906 1836 1049
rect 2141 1048 2142 1183
rect 1787 906 1788 1051
rect 1835 1050 1836 1183
rect 1787 1052 1788 1183
rect 1811 906 1812 1053
rect 1661 906 1662 1055
rect 1811 1054 1812 1183
rect 1859 906 1860 1055
rect 2051 1054 2052 1183
rect 1859 1056 1860 1183
rect 2022 906 2023 1057
rect 1706 906 1707 1059
rect 2021 1058 2022 1183
rect 1877 906 1878 1061
rect 2099 1060 2100 1183
rect 1805 906 1806 1063
rect 1877 1062 1878 1183
rect 1715 906 1716 1065
rect 1805 1064 1806 1183
rect 1715 1066 1716 1183
rect 2421 1066 2422 1183
rect 1889 906 1890 1069
rect 2171 1068 2172 1183
rect 1799 906 1800 1071
rect 1889 1070 1890 1183
rect 1799 1072 1800 1183
rect 2367 1072 2368 1183
rect 1895 906 1896 1075
rect 2081 1074 2082 1183
rect 1895 1076 1896 1183
rect 1967 906 1968 1077
rect 1907 906 1908 1079
rect 2321 1078 2322 1183
rect 1571 906 1572 1081
rect 1907 1080 1908 1183
rect 1913 906 1914 1081
rect 2442 1080 2443 1183
rect 1913 1082 1914 1183
rect 1928 906 1929 1083
rect 1916 906 1917 1085
rect 2105 1084 2106 1183
rect 1919 906 1920 1087
rect 2255 1086 2256 1183
rect 1655 906 1656 1089
rect 1919 1088 1920 1183
rect 1433 906 1434 1091
rect 1655 1090 1656 1183
rect 1434 1092 1435 1183
rect 2327 1092 2328 1183
rect 1922 906 1923 1095
rect 2252 1094 2253 1183
rect 1736 906 1737 1097
rect 1922 1096 1923 1183
rect 1441 1098 1442 1183
rect 1736 1098 1737 1183
rect 1925 906 1926 1099
rect 2291 1098 2292 1183
rect 1925 1100 1926 1183
rect 2029 906 2030 1101
rect 1931 906 1932 1103
rect 2438 1102 2439 1183
rect 1841 906 1842 1105
rect 1931 1104 1932 1183
rect 1841 1106 1842 1183
rect 2018 906 2019 1107
rect 1934 906 1935 1109
rect 1943 1108 1944 1183
rect 1937 906 1938 1111
rect 2330 1110 2331 1183
rect 1937 1112 1938 1183
rect 2032 906 2033 1113
rect 1446 906 1447 1115
rect 2033 1114 2034 1183
rect 1445 1116 1446 1183
rect 1661 1116 1662 1183
rect 1940 906 1941 1117
rect 2123 1116 2124 1183
rect 1952 906 1953 1119
rect 2339 1118 2340 1183
rect 1955 906 1956 1121
rect 2075 1120 2076 1183
rect 1610 906 1611 1123
rect 1955 1122 1956 1183
rect 1958 906 1959 1123
rect 2258 1122 2259 1183
rect 1961 906 1962 1125
rect 2195 1124 2196 1183
rect 1961 1126 1962 1183
rect 2389 1126 2390 1183
rect 1964 906 1965 1129
rect 2057 1128 2058 1183
rect 1974 906 1975 1131
rect 2294 1130 2295 1183
rect 1604 906 1605 1133
rect 1973 1132 1974 1183
rect 1977 906 1978 1133
rect 2333 1132 2334 1183
rect 1986 906 1987 1135
rect 2249 1134 2250 1183
rect 1847 906 1848 1137
rect 1985 1136 1986 1183
rect 1847 1138 1848 1183
rect 1971 906 1972 1139
rect 1992 906 1993 1139
rect 2027 1138 2028 1183
rect 1991 1140 1992 1183
rect 1999 906 2000 1141
rect 1996 906 1997 1143
rect 2234 1142 2235 1183
rect 1997 1144 1998 1183
rect 2348 1144 2349 1183
rect 2003 906 2004 1147
rect 2201 1146 2202 1183
rect 1989 906 1990 1149
rect 2003 1148 2004 1183
rect 2006 906 2007 1149
rect 2207 1148 2208 1183
rect 2009 906 2010 1151
rect 2358 1150 2359 1183
rect 1453 906 1454 1153
rect 2009 1152 2010 1183
rect 1452 1154 1453 1183
rect 1580 1154 1581 1183
rect 2012 906 2013 1155
rect 2361 1154 2362 1183
rect 1634 906 1635 1157
rect 2012 1156 2013 1183
rect 2025 906 2026 1157
rect 2117 1156 2118 1183
rect 2039 906 2040 1159
rect 2138 1158 2139 1183
rect 2036 906 2037 1161
rect 2039 1160 2040 1183
rect 2036 1162 2037 1183
rect 2431 1162 2432 1183
rect 2135 1164 2136 1183
rect 2435 1164 2436 1183
rect 2189 1166 2190 1183
rect 2445 1166 2446 1183
rect 2231 1168 2232 1183
rect 2428 1168 2429 1183
rect 2297 1170 2298 1183
rect 2352 1170 2353 1183
rect 2336 1172 2337 1183
rect 2392 1172 2393 1183
rect 2342 1174 2343 1183
rect 2355 1174 2356 1183
rect 2383 1174 2384 1183
rect 2410 1174 2411 1183
rect 2386 1176 2387 1183
rect 2407 1176 2408 1183
rect 2401 1178 2402 1183
rect 2417 1178 2418 1183
rect 2404 1180 2405 1183
rect 2414 1180 2415 1183
rect 1417 1187 1418 1190
rect 1589 1187 1590 1190
rect 1417 1191 1418 1572
rect 1967 1191 1968 1572
rect 1420 1187 1421 1194
rect 2066 1193 2067 1572
rect 1427 1187 1428 1196
rect 2282 1187 2283 1196
rect 1427 1197 1428 1572
rect 2060 1197 2061 1572
rect 1434 1187 1435 1200
rect 1739 1187 1740 1200
rect 1438 1187 1439 1202
rect 2054 1201 2055 1572
rect 1438 1203 1439 1572
rect 1655 1187 1656 1204
rect 1448 1187 1449 1206
rect 2583 1205 2584 1572
rect 1448 1207 1449 1572
rect 1835 1187 1836 1208
rect 1455 1187 1456 1210
rect 2036 1187 2037 1210
rect 1455 1211 1456 1572
rect 1571 1211 1572 1572
rect 1462 1187 1463 1214
rect 2078 1213 2079 1572
rect 1466 1215 1467 1572
rect 1631 1187 1632 1216
rect 1474 1187 1475 1218
rect 2252 1187 2253 1218
rect 1473 1219 1474 1572
rect 2156 1219 2157 1572
rect 1476 1221 1477 1572
rect 2669 1221 2670 1572
rect 1480 1223 1481 1572
rect 1520 1187 1521 1224
rect 1483 1187 1484 1226
rect 1901 1187 1902 1226
rect 1483 1227 1484 1572
rect 1589 1227 1590 1572
rect 1490 1187 1491 1230
rect 1973 1187 1974 1230
rect 1471 1187 1472 1232
rect 1973 1231 1974 1572
rect 1493 1187 1494 1234
rect 1835 1233 1836 1572
rect 1502 1187 1503 1236
rect 1886 1235 1887 1572
rect 1505 1187 1506 1238
rect 1592 1187 1593 1238
rect 1514 1187 1515 1240
rect 1583 1239 1584 1572
rect 1523 1241 1524 1572
rect 1676 1187 1677 1242
rect 1529 1243 1530 1572
rect 2549 1243 2550 1572
rect 1547 1245 1548 1572
rect 1922 1187 1923 1246
rect 1550 1187 1551 1248
rect 1970 1247 1971 1572
rect 1559 1249 1560 1572
rect 2352 1187 2353 1250
rect 1577 1251 1578 1572
rect 2324 1187 2325 1252
rect 1631 1253 1632 1572
rect 2237 1187 2238 1254
rect 1643 1187 1644 1256
rect 2421 1187 2422 1256
rect 1712 1187 1713 1258
rect 2102 1257 2103 1572
rect 1781 1259 1782 1572
rect 2015 1187 2016 1260
rect 1486 1187 1487 1262
rect 2015 1261 2016 1572
rect 1487 1263 1488 1572
rect 2057 1187 2058 1264
rect 1598 1187 1599 1266
rect 2057 1265 2058 1572
rect 1793 1187 1794 1268
rect 2225 1267 2226 1572
rect 1793 1269 1794 1572
rect 2189 1187 2190 1270
rect 1757 1187 1758 1272
rect 2189 1271 2190 1572
rect 1757 1273 1758 1572
rect 2021 1187 2022 1274
rect 1829 1187 1830 1276
rect 2367 1187 2368 1276
rect 1829 1277 1830 1572
rect 2087 1187 2088 1278
rect 1685 1187 1686 1280
rect 2087 1279 2088 1572
rect 1685 1281 1686 1572
rect 2213 1187 2214 1282
rect 1841 1187 1842 1284
rect 2642 1283 2643 1572
rect 1841 1285 1842 1572
rect 1955 1187 1956 1286
rect 1847 1187 1848 1288
rect 2243 1287 2244 1572
rect 1459 1187 1460 1290
rect 1847 1289 1848 1572
rect 1459 1291 1460 1572
rect 2063 1187 2064 1292
rect 1673 1187 1674 1294
rect 2063 1293 2064 1572
rect 1574 1187 1575 1296
rect 1673 1295 1674 1572
rect 1859 1187 1860 1296
rect 2237 1295 2238 1572
rect 1859 1297 1860 1572
rect 2009 1187 2010 1298
rect 1424 1187 1425 1300
rect 2009 1299 2010 1572
rect 1424 1301 1425 1572
rect 1499 1301 1500 1572
rect 1889 1187 1890 1302
rect 2374 1187 2375 1302
rect 1595 1187 1596 1304
rect 2375 1303 2376 1572
rect 1595 1305 1596 1572
rect 2276 1187 2277 1306
rect 1889 1307 1890 1572
rect 2099 1187 2100 1308
rect 1703 1187 1704 1310
rect 2099 1309 2100 1572
rect 1703 1311 1704 1572
rect 2111 1187 2112 1312
rect 1895 1187 1896 1314
rect 2213 1313 2214 1572
rect 1895 1315 1896 1572
rect 2048 1187 2049 1316
rect 1901 1317 1902 1572
rect 1919 1187 1920 1318
rect 1420 1319 1421 1572
rect 1919 1319 1920 1572
rect 1925 1187 1926 1320
rect 2285 1319 2286 1572
rect 1865 1187 1866 1322
rect 1925 1321 1926 1572
rect 1865 1323 1866 1572
rect 2093 1187 2094 1324
rect 1637 1187 1638 1326
rect 2093 1325 2094 1572
rect 1452 1187 1453 1328
rect 1637 1327 1638 1572
rect 1452 1329 1453 1572
rect 1907 1187 1908 1330
rect 1871 1187 1872 1332
rect 1907 1331 1908 1572
rect 1727 1187 1728 1334
rect 1871 1333 1872 1572
rect 1727 1335 1728 1572
rect 2153 1187 2154 1336
rect 1751 1187 1752 1338
rect 2153 1337 2154 1572
rect 1751 1339 1752 1572
rect 2033 1187 2034 1340
rect 1613 1187 1614 1342
rect 2033 1341 2034 1572
rect 1613 1343 1614 1572
rect 2240 1187 2241 1344
rect 1931 1187 1932 1346
rect 2279 1345 2280 1572
rect 1931 1347 1932 1572
rect 2105 1187 2106 1348
rect 1943 1187 1944 1350
rect 2303 1349 2304 1572
rect 1943 1351 1944 1572
rect 2027 1187 2028 1352
rect 1949 1353 1950 1572
rect 2543 1353 2544 1572
rect 1985 1187 1986 1356
rect 2027 1355 2028 1572
rect 1763 1187 1764 1358
rect 1985 1357 1986 1572
rect 1763 1359 1764 1572
rect 2177 1187 2178 1360
rect 1715 1187 1716 1362
rect 2177 1361 2178 1572
rect 1715 1363 1716 1572
rect 2219 1187 2220 1364
rect 1787 1187 1788 1366
rect 2219 1365 2220 1572
rect 1431 1187 1432 1368
rect 1787 1367 1788 1572
rect 1431 1369 1432 1572
rect 1505 1369 1506 1572
rect 1991 1187 1992 1370
rect 2315 1369 2316 1572
rect 1991 1371 1992 1572
rect 2635 1371 2636 1572
rect 2003 1187 2004 1374
rect 2111 1373 2112 1572
rect 1775 1187 1776 1376
rect 2003 1375 2004 1572
rect 1775 1377 1776 1572
rect 2183 1187 2184 1378
rect 2012 1187 2013 1380
rect 2024 1379 2025 1572
rect 2045 1187 2046 1380
rect 2108 1379 2109 1572
rect 1607 1187 1608 1382
rect 2045 1381 2046 1572
rect 2105 1381 2106 1572
rect 2371 1187 2372 1382
rect 2117 1187 2118 1384
rect 2381 1383 2382 1572
rect 1805 1187 1806 1386
rect 2117 1385 2118 1572
rect 1805 1387 1806 1572
rect 2069 1187 2070 1388
rect 1709 1187 1710 1390
rect 2069 1389 2070 1572
rect 1709 1391 1710 1572
rect 2129 1187 2130 1392
rect 2051 1187 2052 1394
rect 2129 1393 2130 1572
rect 1619 1187 1620 1396
rect 2051 1395 2052 1572
rect 1526 1187 1527 1398
rect 1619 1397 1620 1572
rect 2123 1187 2124 1398
rect 2351 1397 2352 1572
rect 1661 1187 1662 1400
rect 2123 1399 2124 1572
rect 1556 1187 1557 1402
rect 1661 1401 1662 1572
rect 2135 1187 2136 1402
rect 2420 1401 2421 1572
rect 1667 1187 1668 1404
rect 2135 1403 2136 1572
rect 1568 1187 1569 1406
rect 1667 1405 1668 1572
rect 2138 1187 2139 1406
rect 2309 1405 2310 1572
rect 2141 1187 2142 1408
rect 2369 1407 2370 1572
rect 1913 1187 1914 1410
rect 2141 1409 2142 1572
rect 1586 1187 1587 1412
rect 1913 1411 1914 1572
rect 2183 1411 2184 1572
rect 2392 1187 2393 1412
rect 2195 1187 2196 1414
rect 2453 1413 2454 1572
rect 1769 1187 1770 1416
rect 2195 1415 2196 1572
rect 1462 1417 1463 1572
rect 1769 1417 1770 1572
rect 2198 1417 2199 1572
rect 2216 1187 2217 1418
rect 2204 1419 2205 1572
rect 2255 1187 2256 1420
rect 1961 1187 1962 1422
rect 2255 1421 2256 1572
rect 1961 1423 1962 1572
rect 2540 1423 2541 1572
rect 2207 1187 2208 1426
rect 2447 1425 2448 1572
rect 1877 1187 1878 1428
rect 2207 1427 2208 1572
rect 1877 1429 1878 1572
rect 1883 1187 1884 1430
rect 1490 1431 1491 1572
rect 1883 1431 1884 1572
rect 2231 1187 2232 1432
rect 2477 1431 2478 1572
rect 1799 1187 1800 1434
rect 2231 1433 2232 1572
rect 2249 1187 2250 1434
rect 2501 1433 2502 1572
rect 1853 1187 1854 1436
rect 2249 1435 2250 1572
rect 2258 1187 2259 1436
rect 2507 1435 2508 1572
rect 2261 1437 2262 1572
rect 2336 1187 2337 1438
rect 2267 1439 2268 1572
rect 2639 1439 2640 1572
rect 2273 1441 2274 1572
rect 2389 1187 2390 1442
rect 2288 1187 2289 1444
rect 2495 1443 2496 1572
rect 2291 1187 2292 1446
rect 2498 1445 2499 1572
rect 2291 1447 2292 1572
rect 2632 1447 2633 1572
rect 2294 1187 2295 1450
rect 2537 1449 2538 1572
rect 2297 1187 2298 1452
rect 2513 1451 2514 1572
rect 1937 1187 1938 1454
rect 2297 1453 2298 1572
rect 1817 1187 1818 1456
rect 1937 1455 1938 1572
rect 1679 1187 1680 1458
rect 1817 1457 1818 1572
rect 1580 1187 1581 1460
rect 1679 1459 1680 1572
rect 2321 1187 2322 1460
rect 2378 1459 2379 1572
rect 1997 1187 1998 1462
rect 2321 1461 2322 1572
rect 1979 1187 1980 1464
rect 1997 1463 1998 1572
rect 1811 1187 1812 1466
rect 1979 1465 1980 1572
rect 1601 1187 1602 1468
rect 1811 1467 1812 1572
rect 1441 1187 1442 1470
rect 1601 1469 1602 1572
rect 1441 1471 1442 1572
rect 1955 1471 1956 1572
rect 2327 1187 2328 1472
rect 2564 1471 2565 1572
rect 2327 1473 2328 1572
rect 2703 1473 2704 1572
rect 2330 1187 2331 1476
rect 2465 1475 2466 1572
rect 2333 1187 2334 1478
rect 2570 1477 2571 1572
rect 2075 1187 2076 1480
rect 2333 1479 2334 1572
rect 1625 1187 1626 1482
rect 2075 1481 2076 1572
rect 1532 1187 1533 1484
rect 1625 1483 1626 1572
rect 1532 1485 1533 1572
rect 2147 1485 2148 1572
rect 2339 1187 2340 1486
rect 2546 1485 2547 1572
rect 2039 1187 2040 1488
rect 2339 1487 2340 1572
rect 1649 1187 1650 1490
rect 2039 1489 2040 1572
rect 1649 1491 1650 1572
rect 1736 1187 1737 1492
rect 2342 1187 2343 1492
rect 2519 1491 2520 1572
rect 2345 1187 2346 1494
rect 2687 1493 2688 1572
rect 2345 1495 2346 1572
rect 2579 1495 2580 1572
rect 2348 1187 2349 1498
rect 2573 1497 2574 1572
rect 2355 1187 2356 1500
rect 2525 1499 2526 1572
rect 2358 1187 2359 1502
rect 2595 1501 2596 1572
rect 1469 1503 1470 1572
rect 2357 1503 2358 1572
rect 2361 1187 2362 1504
rect 2531 1503 2532 1572
rect 2364 1187 2365 1506
rect 2424 1187 2425 1506
rect 2081 1187 2082 1508
rect 2363 1507 2364 1572
rect 1445 1187 1446 1510
rect 2081 1509 2082 1572
rect 1445 1511 1446 1572
rect 2021 1511 2022 1572
rect 2234 1187 2235 1512
rect 2423 1511 2424 1572
rect 2383 1187 2384 1514
rect 2435 1187 2436 1514
rect 2386 1187 2387 1516
rect 2607 1515 2608 1572
rect 2393 1517 2394 1572
rect 2700 1517 2701 1572
rect 2399 1519 2400 1572
rect 2445 1187 2446 1520
rect 2401 1187 2402 1522
rect 2651 1521 2652 1572
rect 2404 1187 2405 1524
rect 2645 1523 2646 1572
rect 2405 1525 2406 1572
rect 2710 1525 2711 1572
rect 2407 1187 2408 1528
rect 2622 1527 2623 1572
rect 2410 1187 2411 1530
rect 2619 1529 2620 1572
rect 2414 1187 2415 1532
rect 2666 1531 2667 1572
rect 2417 1187 2418 1534
rect 2663 1533 2664 1572
rect 2417 1535 2418 1572
rect 2714 1535 2715 1572
rect 2428 1187 2429 1538
rect 2483 1537 2484 1572
rect 2431 1187 2432 1540
rect 2486 1539 2487 1572
rect 2438 1187 2439 1542
rect 2707 1541 2708 1572
rect 2442 1187 2443 1544
rect 2504 1543 2505 1572
rect 2201 1187 2202 1546
rect 2441 1545 2442 1572
rect 1823 1187 1824 1548
rect 2201 1547 2202 1572
rect 1733 1187 1734 1550
rect 1823 1549 1824 1572
rect 1733 1551 1734 1572
rect 2159 1187 2160 1552
rect 1697 1187 1698 1554
rect 2159 1553 2160 1572
rect 1434 1555 1435 1572
rect 1697 1555 1698 1572
rect 2459 1555 2460 1572
rect 2672 1555 2673 1572
rect 2489 1557 2490 1572
rect 2586 1557 2587 1572
rect 2558 1559 2559 1572
rect 2723 1559 2724 1572
rect 2561 1561 2562 1572
rect 2720 1561 2721 1572
rect 2576 1563 2577 1572
rect 2717 1563 2718 1572
rect 2601 1565 2602 1572
rect 2628 1565 2629 1572
rect 2604 1567 2605 1572
rect 2625 1567 2626 1572
rect 2675 1567 2676 1572
rect 2693 1567 2694 1572
rect 2690 1569 2691 1572
rect 2696 1569 2697 1572
rect 1424 1576 1425 1579
rect 1517 1578 1518 2029
rect 1417 1576 1418 1581
rect 1424 1580 1425 2029
rect 1427 1576 1428 1581
rect 2174 1580 2175 2029
rect 1431 1576 1432 1583
rect 2045 1576 2046 1583
rect 1445 1576 1446 1585
rect 1931 1576 1932 1585
rect 1448 1576 1449 1587
rect 1469 1576 1470 1587
rect 1448 1588 1449 2029
rect 1619 1576 1620 1589
rect 1452 1576 1453 1591
rect 1787 1576 1788 1591
rect 1452 1592 1453 2029
rect 1865 1576 1866 1593
rect 1455 1576 1456 1595
rect 1781 1576 1782 1595
rect 1466 1576 1467 1597
rect 2318 1596 2319 2029
rect 1476 1576 1477 1599
rect 2246 1598 2247 2029
rect 1469 1600 1470 2029
rect 1476 1600 1477 2029
rect 1483 1576 1484 1601
rect 1583 1576 1584 1601
rect 1485 1602 1486 2029
rect 2123 1576 2124 1603
rect 1487 1576 1488 1605
rect 1883 1576 1884 1605
rect 1502 1606 1503 2029
rect 2369 1576 2370 1607
rect 1505 1576 1506 1609
rect 1541 1608 1542 2029
rect 1532 1576 1533 1611
rect 2900 1610 2901 2029
rect 1565 1612 1566 2029
rect 2078 1576 2079 1613
rect 1577 1576 1578 1615
rect 1607 1614 1608 2029
rect 1547 1576 1548 1617
rect 1577 1616 1578 2029
rect 1473 1576 1474 1619
rect 1547 1618 1548 2029
rect 1473 1620 1474 2029
rect 2525 1576 2526 1621
rect 1625 1576 1626 1623
rect 1655 1622 1656 2029
rect 1480 1576 1481 1625
rect 1625 1624 1626 2029
rect 1643 1624 1644 2029
rect 1886 1576 1887 1625
rect 1661 1576 1662 1627
rect 1691 1626 1692 2029
rect 1631 1576 1632 1629
rect 1661 1628 1662 2029
rect 1589 1576 1590 1631
rect 1631 1630 1632 2029
rect 1679 1576 1680 1631
rect 2778 1630 2779 2029
rect 1667 1576 1668 1633
rect 1679 1632 1680 2029
rect 1709 1576 1710 1633
rect 1739 1632 1740 2029
rect 1685 1576 1686 1635
rect 1709 1634 1710 2029
rect 1745 1576 1746 1635
rect 1781 1634 1782 2029
rect 1715 1576 1716 1637
rect 1745 1636 1746 2029
rect 1751 1576 1752 1637
rect 1799 1636 1800 2029
rect 1721 1576 1722 1639
rect 1751 1638 1752 2029
rect 1703 1576 1704 1641
rect 1721 1640 1722 2029
rect 1673 1576 1674 1643
rect 1703 1642 1704 2029
rect 1649 1576 1650 1645
rect 1673 1644 1674 2029
rect 1613 1576 1614 1647
rect 1649 1646 1650 2029
rect 1571 1576 1572 1649
rect 1613 1648 1614 2029
rect 1571 1650 1572 2029
rect 2156 1576 2157 1651
rect 1763 1576 1764 1653
rect 1787 1652 1788 2029
rect 1727 1576 1728 1655
rect 1763 1654 1764 2029
rect 1697 1576 1698 1657
rect 1727 1656 1728 2029
rect 1637 1576 1638 1659
rect 1697 1658 1698 2029
rect 1595 1576 1596 1661
rect 1637 1660 1638 2029
rect 1559 1576 1560 1663
rect 1595 1662 1596 2029
rect 1523 1576 1524 1665
rect 1559 1664 1560 2029
rect 1523 1666 1524 2029
rect 2060 1576 2061 1667
rect 1805 1576 1806 1669
rect 1883 1668 1884 2029
rect 1434 1576 1435 1671
rect 1805 1670 1806 2029
rect 1817 1576 1818 1671
rect 1853 1670 1854 2029
rect 1775 1576 1776 1673
rect 1817 1672 1818 2029
rect 1601 1576 1602 1675
rect 1775 1674 1776 2029
rect 1835 1576 1836 1675
rect 1865 1674 1866 2029
rect 1835 1676 1836 2029
rect 2867 1676 2868 2029
rect 1889 1576 1890 1679
rect 2826 1678 2827 2029
rect 1841 1576 1842 1681
rect 1889 1680 1890 2029
rect 1841 1682 1842 2029
rect 2635 1576 2636 1683
rect 1931 1684 1932 2029
rect 2291 1576 2292 1685
rect 1943 1576 1944 1687
rect 2543 1576 2544 1687
rect 1895 1576 1896 1689
rect 1943 1688 1944 2029
rect 1970 1576 1971 1689
rect 2072 1688 2073 2029
rect 1973 1576 1974 1691
rect 2045 1690 2046 2029
rect 1793 1576 1794 1693
rect 1973 1692 1974 2029
rect 1455 1694 1456 2029
rect 1793 1694 1794 2029
rect 1991 1576 1992 1695
rect 2771 1694 2772 2029
rect 1937 1576 1938 1697
rect 1991 1696 1992 2029
rect 1490 1576 1491 1699
rect 1937 1698 1938 2029
rect 2021 1576 2022 1699
rect 2123 1698 2124 2029
rect 1979 1576 1980 1701
rect 2021 1700 2022 2029
rect 1417 1702 1418 2029
rect 1979 1702 1980 2029
rect 2054 1576 2055 1703
rect 2168 1702 2169 2029
rect 2066 1576 2067 1705
rect 2162 1704 2163 2029
rect 2108 1576 2109 1707
rect 2222 1706 2223 2029
rect 2177 1576 2178 1709
rect 2291 1708 2292 2029
rect 1441 1576 1442 1711
rect 2177 1710 2178 2029
rect 1441 1712 1442 2029
rect 1847 1576 1848 1713
rect 1811 1576 1812 1715
rect 1847 1714 1848 2029
rect 1757 1576 1758 1717
rect 1811 1716 1812 2029
rect 2198 1576 2199 1717
rect 2324 1716 2325 2029
rect 2102 1576 2103 1719
rect 2198 1718 2199 2029
rect 2204 1576 2205 1719
rect 2270 1718 2271 2029
rect 1529 1576 1530 1721
rect 2204 1720 2205 2029
rect 1499 1576 1500 1723
rect 1529 1722 1530 2029
rect 1499 1724 1500 2029
rect 2741 1724 2742 2029
rect 2243 1576 2244 1727
rect 2369 1726 2370 2029
rect 2153 1576 2154 1729
rect 2243 1728 2244 2029
rect 2033 1576 2034 1731
rect 2153 1730 2154 2029
rect 1955 1576 1956 1733
rect 2033 1732 2034 2029
rect 1907 1576 1908 1735
rect 1955 1734 1956 2029
rect 1859 1576 1860 1737
rect 1907 1736 1908 2029
rect 1823 1576 1824 1739
rect 1859 1738 1860 2029
rect 1459 1576 1460 1741
rect 1823 1740 1824 2029
rect 1459 1742 1460 2029
rect 2126 1742 2127 2029
rect 2261 1576 2262 1743
rect 2411 1742 2412 2029
rect 2147 1576 2148 1745
rect 2261 1744 2262 2029
rect 2063 1576 2064 1747
rect 2147 1746 2148 2029
rect 1420 1576 1421 1749
rect 2063 1748 2064 2029
rect 1420 1750 1421 2029
rect 1913 1576 1914 1751
rect 1829 1576 1830 1753
rect 1913 1752 1914 2029
rect 1769 1576 1770 1755
rect 1829 1754 1830 2029
rect 1733 1576 1734 1757
rect 1769 1756 1770 2029
rect 1427 1758 1428 2029
rect 1733 1758 1734 2029
rect 2285 1576 2286 1759
rect 2429 1758 2430 2029
rect 2165 1576 2166 1761
rect 2285 1760 2286 2029
rect 2051 1576 2052 1763
rect 2165 1762 2166 2029
rect 1488 1764 1489 2029
rect 2051 1764 2052 2029
rect 2321 1576 2322 1765
rect 2435 1764 2436 2029
rect 1492 1766 1493 2029
rect 2321 1766 2322 2029
rect 2327 1576 2328 1767
rect 2471 1766 2472 2029
rect 2207 1576 2208 1769
rect 2327 1768 2328 2029
rect 2093 1576 2094 1771
rect 2207 1770 2208 2029
rect 2093 1772 2094 2029
rect 2840 1772 2841 2029
rect 2333 1576 2334 1775
rect 2579 1576 2580 1775
rect 2219 1576 2220 1777
rect 2333 1776 2334 2029
rect 2105 1576 2106 1779
rect 2219 1778 2220 2029
rect 1466 1780 1467 2029
rect 2105 1780 2106 2029
rect 2378 1576 2379 1781
rect 2492 1780 2493 2029
rect 2381 1576 2382 1783
rect 2525 1782 2526 2029
rect 2255 1576 2256 1785
rect 2381 1784 2382 2029
rect 2171 1576 2172 1787
rect 2255 1786 2256 2029
rect 2057 1576 2058 1789
rect 2171 1788 2172 2029
rect 1985 1576 1986 1791
rect 2057 1790 2058 2029
rect 1462 1576 1463 1793
rect 1985 1792 1986 2029
rect 1462 1794 1463 2029
rect 2024 1576 2025 1795
rect 2387 1794 2388 2029
rect 2775 1794 2776 2029
rect 2423 1576 2424 1797
rect 2579 1796 2580 2029
rect 2279 1576 2280 1799
rect 2423 1798 2424 2029
rect 2279 1800 2280 2029
rect 2768 1800 2769 2029
rect 2441 1576 2442 1803
rect 2707 1576 2708 1803
rect 2303 1576 2304 1805
rect 2441 1804 2442 2029
rect 2189 1576 2190 1807
rect 2303 1806 2304 2029
rect 2141 1576 2142 1809
rect 2189 1808 2190 2029
rect 2099 1576 2100 1811
rect 2141 1810 2142 2029
rect 2003 1576 2004 1813
rect 2099 1812 2100 2029
rect 1961 1576 1962 1815
rect 2003 1814 2004 2029
rect 1925 1576 1926 1817
rect 1961 1816 1962 2029
rect 1877 1576 1878 1819
rect 1925 1818 1926 2029
rect 1431 1820 1432 2029
rect 1877 1820 1878 2029
rect 2447 1576 2448 1821
rect 2555 1820 2556 2029
rect 2309 1576 2310 1823
rect 2447 1822 2448 2029
rect 2309 1824 2310 2029
rect 2918 1824 2919 2029
rect 2459 1576 2460 1827
rect 2615 1826 2616 2029
rect 2315 1576 2316 1829
rect 2459 1828 2460 2029
rect 2486 1576 2487 1829
rect 2630 1828 2631 2029
rect 2498 1576 2499 1831
rect 2583 1576 2584 1831
rect 2501 1576 2502 1833
rect 2654 1832 2655 2029
rect 2357 1576 2358 1835
rect 2501 1834 2502 2029
rect 2213 1576 2214 1837
rect 2357 1836 2358 2029
rect 2117 1576 2118 1839
rect 2213 1838 2214 2029
rect 2117 1840 2118 2029
rect 2393 1576 2394 1841
rect 2393 1842 2394 2029
rect 2639 1576 2640 1843
rect 2489 1576 2490 1845
rect 2639 1844 2640 2029
rect 2375 1576 2376 1847
rect 2489 1846 2490 2029
rect 2249 1576 2250 1849
rect 2375 1848 2376 2029
rect 2135 1576 2136 1851
rect 2249 1850 2250 2029
rect 2069 1576 2070 1853
rect 2135 1852 2136 2029
rect 1967 1576 1968 1855
rect 2069 1854 2070 2029
rect 1919 1576 1920 1857
rect 1967 1856 1968 2029
rect 1871 1576 1872 1859
rect 1919 1858 1920 2029
rect 1434 1860 1435 2029
rect 1871 1860 1872 2029
rect 2507 1576 2508 1861
rect 2657 1860 2658 2029
rect 2363 1576 2364 1863
rect 2507 1862 2508 2029
rect 2237 1576 2238 1865
rect 2363 1864 2364 2029
rect 2237 1866 2238 2029
rect 2642 1576 2643 1867
rect 2540 1576 2541 1869
rect 2672 1576 2673 1869
rect 2543 1870 2544 2029
rect 2907 1870 2908 2029
rect 2546 1576 2547 1873
rect 2744 1872 2745 2029
rect 2549 1576 2550 1875
rect 2747 1874 2748 2029
rect 2399 1576 2400 1877
rect 2549 1876 2550 2029
rect 2267 1576 2268 1879
rect 2399 1878 2400 2029
rect 2201 1576 2202 1881
rect 2267 1880 2268 2029
rect 2075 1576 2076 1883
rect 2201 1882 2202 2029
rect 2027 1576 2028 1885
rect 2075 1884 2076 2029
rect 2027 1886 2028 2029
rect 2837 1886 2838 2029
rect 2564 1576 2565 1889
rect 2756 1888 2757 2029
rect 2570 1576 2571 1891
rect 2830 1890 2831 2029
rect 2573 1576 2574 1893
rect 2632 1576 2633 1893
rect 2417 1576 2418 1895
rect 2573 1894 2574 2029
rect 2273 1576 2274 1897
rect 2417 1896 2418 2029
rect 2159 1576 2160 1899
rect 2273 1898 2274 2029
rect 2039 1576 2040 1901
rect 2159 1900 2160 2029
rect 1495 1902 1496 2029
rect 2039 1902 2040 2029
rect 2465 1576 2466 1903
rect 2633 1902 2634 2029
rect 2465 1904 2466 2029
rect 2870 1904 2871 2029
rect 2576 1576 2577 1907
rect 2911 1906 2912 2029
rect 2591 1908 2592 2029
rect 2669 1576 2670 1909
rect 2513 1576 2514 1911
rect 2669 1910 2670 2029
rect 2595 1576 2596 1913
rect 2787 1912 2788 2029
rect 2597 1914 2598 2029
rect 2823 1914 2824 2029
rect 2601 1576 2602 1917
rect 2820 1916 2821 2029
rect 2604 1576 2605 1919
rect 2781 1918 2782 2029
rect 2453 1576 2454 1921
rect 2603 1920 2604 2029
rect 2297 1576 2298 1923
rect 2453 1922 2454 2029
rect 2195 1576 2196 1925
rect 2297 1924 2298 2029
rect 2081 1576 2082 1927
rect 2195 1926 2196 2029
rect 2081 1928 2082 2029
rect 2111 1576 2112 1929
rect 2009 1576 2010 1931
rect 2111 1930 2112 2029
rect 2009 1932 2010 2029
rect 2129 1576 2130 1933
rect 2129 1934 2130 2029
rect 2904 1934 2905 2029
rect 2607 1576 2608 1937
rect 2799 1936 2800 2029
rect 2609 1938 2610 2029
rect 2717 1576 2718 1939
rect 2619 1576 2620 1941
rect 2811 1940 2812 2029
rect 2622 1576 2623 1943
rect 2814 1942 2815 2029
rect 2477 1576 2478 1945
rect 2621 1944 2622 2029
rect 2345 1576 2346 1947
rect 2477 1946 2478 2029
rect 2225 1576 2226 1949
rect 2345 1948 2346 2029
rect 2183 1576 2184 1951
rect 2225 1950 2226 2029
rect 2087 1576 2088 1953
rect 2183 1952 2184 2029
rect 2015 1576 2016 1955
rect 2087 1954 2088 2029
rect 1997 1576 1998 1957
rect 2015 1956 2016 2029
rect 1949 1576 1950 1959
rect 1997 1958 1998 2029
rect 1901 1576 1902 1961
rect 1949 1960 1950 2029
rect 1445 1962 1446 2029
rect 1901 1962 1902 2029
rect 2625 1576 2626 1963
rect 2817 1962 2818 2029
rect 2628 1576 2629 1965
rect 2925 1964 2926 2029
rect 2483 1576 2484 1967
rect 2627 1966 2628 2029
rect 2339 1576 2340 1969
rect 2483 1968 2484 2029
rect 2339 1970 2340 2029
rect 2703 1576 2704 1971
rect 2645 1576 2646 1973
rect 2843 1972 2844 2029
rect 2651 1576 2652 1975
rect 2849 1974 2850 2029
rect 2651 1976 2652 2029
rect 2928 1976 2929 2029
rect 2663 1576 2664 1979
rect 2861 1978 2862 2029
rect 2495 1576 2496 1981
rect 2663 1980 2664 2029
rect 2351 1576 2352 1983
rect 2495 1982 2496 2029
rect 2231 1576 2232 1985
rect 2351 1984 2352 2029
rect 2231 1986 2232 2029
rect 2708 1986 2709 2029
rect 2666 1576 2667 1989
rect 2864 1988 2865 2029
rect 2586 1576 2587 1991
rect 2666 1990 2667 2029
rect 2405 1576 2406 1993
rect 2585 1992 2586 2029
rect 2405 1994 2406 2029
rect 2921 1994 2922 2029
rect 2675 1576 2676 1997
rect 2873 1996 2874 2029
rect 2519 1576 2520 1999
rect 2675 1998 2676 2029
rect 2519 2000 2520 2029
rect 2897 2000 2898 2029
rect 2687 1576 2688 2003
rect 2696 1576 2697 2003
rect 2531 1576 2532 2005
rect 2696 2004 2697 2029
rect 2504 1576 2505 2007
rect 2531 2006 2532 2029
rect 2690 1576 2691 2007
rect 2894 2006 2895 2029
rect 2693 1576 2694 2009
rect 2891 2008 2892 2029
rect 2537 1576 2538 2011
rect 2693 2010 2694 2029
rect 1438 1576 1439 2013
rect 2537 2012 2538 2029
rect 1438 2014 1439 2029
rect 2315 2014 2316 2029
rect 2700 1576 2701 2015
rect 2702 2014 2703 2029
rect 2710 1576 2711 2015
rect 2879 2014 2880 2029
rect 1583 2016 1584 2029
rect 2711 2016 2712 2029
rect 2714 1576 2715 2017
rect 2765 2016 2766 2029
rect 2561 1576 2562 2019
rect 2714 2018 2715 2029
rect 2420 1576 2421 2021
rect 2561 2020 2562 2029
rect 2720 1576 2721 2021
rect 2726 2020 2727 2029
rect 2558 1576 2559 2023
rect 2720 2022 2721 2029
rect 2723 1576 2724 2023
rect 2882 2022 2883 2029
rect 2738 2024 2739 2029
rect 2914 2024 2915 2029
rect 2762 2026 2763 2029
rect 2833 2026 2834 2029
rect 1417 2033 1418 2036
rect 2103 2035 2104 2558
rect 1420 2033 1421 2038
rect 1989 2037 1990 2558
rect 1424 2033 1425 2040
rect 3018 2039 3019 2558
rect 1427 2033 1428 2042
rect 1899 2041 1900 2558
rect 1431 2033 1432 2044
rect 1490 2043 1491 2558
rect 1432 2045 1433 2558
rect 2337 2045 2338 2558
rect 1434 2033 1435 2048
rect 1865 2033 1866 2048
rect 1436 2049 1437 2558
rect 1959 2049 1960 2558
rect 1438 2033 1439 2052
rect 2165 2033 2166 2052
rect 1443 2053 1444 2558
rect 1853 2033 1854 2054
rect 1445 2033 1446 2056
rect 1689 2055 1690 2558
rect 1448 2033 1449 2058
rect 2198 2033 2199 2058
rect 1450 2059 1451 2558
rect 1733 2033 1734 2060
rect 1452 2033 1453 2062
rect 2174 2033 2175 2062
rect 1453 2063 1454 2558
rect 1779 2063 1780 2558
rect 1455 2033 1456 2066
rect 2289 2065 2290 2558
rect 1457 2067 1458 2558
rect 1821 2067 1822 2558
rect 1462 2033 1463 2070
rect 2708 2033 2709 2070
rect 1464 2071 1465 2558
rect 2199 2071 2200 2558
rect 1466 2033 1467 2074
rect 2099 2033 2100 2074
rect 1467 2075 1468 2558
rect 2057 2033 2058 2076
rect 1469 2033 1470 2078
rect 2097 2077 2098 2558
rect 1471 2079 1472 2558
rect 2121 2079 2122 2558
rect 1473 2033 1474 2082
rect 2021 2033 2022 2082
rect 1474 2083 1475 2558
rect 1673 2033 1674 2084
rect 1476 2033 1477 2086
rect 2151 2085 2152 2558
rect 1483 2087 1484 2558
rect 1803 2087 1804 2558
rect 1485 2033 1486 2090
rect 1587 2089 1588 2558
rect 1488 2033 1489 2092
rect 2379 2091 2380 2558
rect 1492 2033 1493 2094
rect 1931 2033 1932 2094
rect 1497 2095 1498 2558
rect 1607 2033 1608 2096
rect 1499 2033 1500 2098
rect 2013 2097 2014 2558
rect 1500 2099 1501 2558
rect 1611 2099 1612 2558
rect 1502 2033 1503 2102
rect 1977 2101 1978 2558
rect 1515 2103 1516 2558
rect 2126 2033 2127 2104
rect 1486 2105 1487 2558
rect 2127 2105 2128 2558
rect 1521 2107 1522 2558
rect 1547 2033 1548 2108
rect 1523 2033 1524 2110
rect 2778 2033 2779 2110
rect 1529 2033 1530 2112
rect 1533 2111 1534 2558
rect 1541 2033 1542 2112
rect 1551 2111 1552 2558
rect 1545 2113 1546 2558
rect 1565 2033 1566 2114
rect 1557 2115 1558 2558
rect 1571 2033 1572 2116
rect 1559 2033 1560 2118
rect 1569 2117 1570 2558
rect 1563 2119 1564 2558
rect 2162 2033 2163 2120
rect 1575 2121 1576 2558
rect 1577 2033 1578 2122
rect 1583 2033 1584 2122
rect 1599 2121 1600 2558
rect 1593 2123 1594 2558
rect 1595 2033 1596 2124
rect 1613 2033 1614 2124
rect 1629 2123 1630 2558
rect 1623 2125 1624 2558
rect 2318 2033 2319 2126
rect 1429 2127 1430 2558
rect 2319 2127 2320 2558
rect 1625 2033 1626 2130
rect 1641 2129 1642 2558
rect 1631 2033 1632 2132
rect 1647 2131 1648 2558
rect 1637 2033 1638 2134
rect 1653 2133 1654 2558
rect 1643 2033 1644 2136
rect 1659 2135 1660 2558
rect 1649 2033 1650 2138
rect 1671 2137 1672 2558
rect 1655 2033 1656 2140
rect 1683 2139 1684 2558
rect 1661 2033 1662 2142
rect 1665 2141 1666 2558
rect 1677 2141 1678 2558
rect 1775 2033 1776 2142
rect 1691 2033 1692 2144
rect 1737 2143 1738 2558
rect 1692 2145 1693 2558
rect 2019 2145 2020 2558
rect 1695 2147 1696 2558
rect 1709 2033 1710 2148
rect 1697 2033 1698 2150
rect 1719 2149 1720 2558
rect 1701 2151 1702 2558
rect 1721 2033 1722 2152
rect 1703 2033 1704 2154
rect 1725 2153 1726 2558
rect 1707 2155 1708 2558
rect 1739 2033 1740 2156
rect 1727 2033 1728 2158
rect 1773 2157 1774 2558
rect 1743 2159 1744 2558
rect 1745 2033 1746 2160
rect 1749 2159 1750 2558
rect 2222 2033 2223 2160
rect 1751 2033 1752 2162
rect 1785 2161 1786 2558
rect 1761 2163 1762 2558
rect 2669 2033 2670 2164
rect 1763 2033 1764 2166
rect 1809 2165 1810 2558
rect 1769 2033 1770 2168
rect 1815 2167 1816 2558
rect 1781 2033 1782 2170
rect 1827 2169 1828 2558
rect 1787 2033 1788 2172
rect 1851 2171 1852 2558
rect 1791 2173 1792 2558
rect 2666 2033 2667 2174
rect 1793 2033 1794 2176
rect 1833 2175 1834 2558
rect 1797 2177 1798 2558
rect 2633 2033 2634 2178
rect 1799 2033 1800 2180
rect 1839 2179 1840 2558
rect 1805 2033 1806 2182
rect 1869 2181 1870 2558
rect 1811 2033 1812 2184
rect 1845 2183 1846 2558
rect 1817 2033 1818 2186
rect 1875 2185 1876 2558
rect 1823 2033 1824 2188
rect 1857 2187 1858 2558
rect 1829 2033 1830 2190
rect 1863 2189 1864 2558
rect 1835 2033 1836 2192
rect 1881 2191 1882 2558
rect 1841 2033 1842 2194
rect 1887 2193 1888 2558
rect 1847 2033 1848 2196
rect 1935 2195 1936 2558
rect 1859 2033 1860 2198
rect 1941 2197 1942 2558
rect 1871 2033 1872 2200
rect 1953 2199 1954 2558
rect 1877 2033 1878 2202
rect 1965 2201 1966 2558
rect 1883 2033 1884 2204
rect 1911 2203 1912 2558
rect 1889 2033 1890 2206
rect 1929 2205 1930 2558
rect 1893 2207 1894 2558
rect 1973 2033 1974 2208
rect 1901 2033 1902 2210
rect 1983 2209 1984 2558
rect 1905 2211 1906 2558
rect 1985 2033 1986 2212
rect 1907 2033 1908 2214
rect 1947 2213 1948 2558
rect 1913 2033 1914 2216
rect 1923 2215 1924 2558
rect 1919 2033 1920 2218
rect 2007 2217 2008 2558
rect 1925 2033 1926 2220
rect 2001 2219 2002 2558
rect 1937 2033 1938 2222
rect 1995 2221 1996 2558
rect 1943 2033 1944 2224
rect 2055 2223 2056 2558
rect 1949 2033 1950 2226
rect 2025 2225 2026 2558
rect 1955 2033 1956 2228
rect 2067 2227 2068 2558
rect 1961 2033 1962 2230
rect 2079 2229 2080 2558
rect 1971 2231 1972 2558
rect 2117 2033 2118 2232
rect 1979 2033 1980 2234
rect 2109 2233 2110 2558
rect 1991 2033 1992 2236
rect 2115 2235 2116 2558
rect 1997 2033 1998 2238
rect 2043 2237 2044 2558
rect 2003 2033 2004 2240
rect 2049 2239 2050 2558
rect 2009 2033 2010 2242
rect 2031 2241 2032 2558
rect 2015 2033 2016 2244
rect 2145 2243 2146 2558
rect 2027 2033 2028 2246
rect 2157 2245 2158 2558
rect 2033 2033 2034 2248
rect 2163 2247 2164 2558
rect 2037 2249 2038 2558
rect 2093 2033 2094 2250
rect 2045 2033 2046 2252
rect 2175 2251 2176 2558
rect 2051 2033 2052 2254
rect 2181 2253 2182 2558
rect 2061 2255 2062 2558
rect 2639 2033 2640 2256
rect 2063 2033 2064 2258
rect 2187 2257 2188 2558
rect 2069 2033 2070 2260
rect 2193 2259 2194 2558
rect 2075 2033 2076 2262
rect 2577 2261 2578 2558
rect 2081 2033 2082 2264
rect 2601 2263 2602 2558
rect 2085 2265 2086 2558
rect 2477 2033 2478 2266
rect 2087 2033 2088 2268
rect 2217 2267 2218 2558
rect 2091 2269 2092 2558
rect 2768 2033 2769 2270
rect 2105 2033 2106 2272
rect 2229 2271 2230 2558
rect 2111 2033 2112 2274
rect 2235 2273 2236 2558
rect 2129 2033 2130 2276
rect 2241 2275 2242 2558
rect 2133 2277 2134 2558
rect 3012 2277 3013 2558
rect 2139 2279 2140 2558
rect 2471 2033 2472 2280
rect 2141 2033 2142 2282
rect 2277 2281 2278 2558
rect 2147 2033 2148 2284
rect 2916 2283 2917 2558
rect 2153 2033 2154 2286
rect 2295 2285 2296 2558
rect 2159 2033 2160 2288
rect 2301 2287 2302 2558
rect 2171 2033 2172 2290
rect 2313 2289 2314 2558
rect 2177 2033 2178 2292
rect 2283 2291 2284 2558
rect 2183 2033 2184 2294
rect 2307 2293 2308 2558
rect 2189 2033 2190 2296
rect 2967 2295 2968 2558
rect 2195 2033 2196 2298
rect 2771 2033 2772 2298
rect 2072 2033 2073 2300
rect 2196 2299 2197 2558
rect 1967 2033 1968 2302
rect 2073 2301 2074 2558
rect 2201 2033 2202 2302
rect 2331 2301 2332 2558
rect 2207 2033 2208 2304
rect 2355 2303 2356 2558
rect 2211 2305 2212 2558
rect 3118 2305 3119 2558
rect 2213 2033 2214 2308
rect 2265 2307 2266 2558
rect 2219 2033 2220 2310
rect 2367 2309 2368 2558
rect 2225 2033 2226 2312
rect 2253 2311 2254 2558
rect 2231 2033 2232 2314
rect 2343 2313 2344 2558
rect 2237 2033 2238 2316
rect 2511 2315 2512 2558
rect 2243 2033 2244 2318
rect 2373 2317 2374 2558
rect 2249 2033 2250 2320
rect 2711 2033 2712 2320
rect 1459 2033 1460 2322
rect 2250 2321 2251 2558
rect 1460 2323 1461 2558
rect 2168 2033 2169 2324
rect 2039 2033 2040 2326
rect 2169 2325 2170 2558
rect 2255 2033 2256 2326
rect 2391 2325 2392 2558
rect 2259 2327 2260 2558
rect 2381 2033 2382 2328
rect 2261 2033 2262 2330
rect 2397 2329 2398 2558
rect 2267 2033 2268 2332
rect 2361 2331 2362 2558
rect 2273 2033 2274 2334
rect 2415 2333 2416 2558
rect 2279 2033 2280 2336
rect 2427 2335 2428 2558
rect 2285 2033 2286 2338
rect 2421 2337 2422 2558
rect 2291 2033 2292 2340
rect 2904 2033 2905 2340
rect 2297 2033 2298 2342
rect 2403 2341 2404 2558
rect 2303 2033 2304 2344
rect 2439 2343 2440 2558
rect 2309 2033 2310 2346
rect 2451 2345 2452 2558
rect 2310 2347 2311 2558
rect 2918 2033 2919 2348
rect 2315 2033 2316 2350
rect 2433 2349 2434 2558
rect 1517 2033 1518 2352
rect 2316 2351 2317 2558
rect 2321 2033 2322 2352
rect 2457 2351 2458 2558
rect 1679 2033 1680 2354
rect 2322 2353 2323 2558
rect 2327 2033 2328 2354
rect 2385 2353 2386 2558
rect 2333 2033 2334 2356
rect 2475 2355 2476 2558
rect 2204 2033 2205 2358
rect 2334 2357 2335 2558
rect 1495 2033 1496 2360
rect 2205 2359 2206 2558
rect 2339 2033 2340 2360
rect 2481 2359 2482 2558
rect 1446 2361 1447 2558
rect 2340 2361 2341 2558
rect 2345 2033 2346 2362
rect 2469 2361 2470 2558
rect 2349 2363 2350 2558
rect 2411 2033 2412 2364
rect 2351 2033 2352 2366
rect 2487 2365 2488 2558
rect 2357 2033 2358 2368
rect 2463 2367 2464 2558
rect 2369 2033 2370 2370
rect 2499 2369 2500 2558
rect 1441 2033 1442 2372
rect 2370 2371 2371 2558
rect 2375 2033 2376 2372
rect 2505 2371 2506 2558
rect 2246 2033 2247 2374
rect 2376 2373 2377 2558
rect 2123 2033 2124 2376
rect 2247 2375 2248 2558
rect 2387 2033 2388 2376
rect 2541 2375 2542 2558
rect 2393 2033 2394 2378
rect 2529 2377 2530 2558
rect 2399 2033 2400 2380
rect 2535 2379 2536 2558
rect 2400 2381 2401 2558
rect 2492 2033 2493 2382
rect 2363 2033 2364 2384
rect 2493 2383 2494 2558
rect 2270 2033 2271 2386
rect 2364 2385 2365 2558
rect 2135 2033 2136 2388
rect 2271 2387 2272 2558
rect 2405 2033 2406 2388
rect 2523 2387 2524 2558
rect 2409 2389 2410 2558
rect 2775 2033 2776 2390
rect 2417 2033 2418 2392
rect 2553 2391 2554 2558
rect 2423 2033 2424 2394
rect 2565 2393 2566 2558
rect 2429 2033 2430 2396
rect 2571 2395 2572 2558
rect 2435 2033 2436 2398
rect 2870 2033 2871 2398
rect 2436 2399 2437 2558
rect 3114 2399 3115 2558
rect 2441 2033 2442 2402
rect 2583 2401 2584 2558
rect 2445 2403 2446 2558
rect 2840 2033 2841 2404
rect 1493 2405 1494 2558
rect 2841 2405 2842 2558
rect 2447 2033 2448 2408
rect 2589 2407 2590 2558
rect 2453 2033 2454 2410
rect 2595 2409 2596 2558
rect 2459 2033 2460 2412
rect 2607 2411 2608 2558
rect 2324 2033 2325 2414
rect 2460 2413 2461 2558
rect 2325 2415 2326 2558
rect 2823 2033 2824 2416
rect 2465 2033 2466 2418
rect 2837 2033 2838 2418
rect 2483 2033 2484 2420
rect 2613 2419 2614 2558
rect 2489 2033 2490 2422
rect 2826 2033 2827 2422
rect 2495 2033 2496 2424
rect 3015 2423 3016 2558
rect 2507 2033 2508 2426
rect 2661 2425 2662 2558
rect 2508 2427 2509 2558
rect 2663 2033 2664 2428
rect 2517 2429 2518 2558
rect 3057 2429 3058 2558
rect 2519 2033 2520 2432
rect 2673 2431 2674 2558
rect 2525 2033 2526 2434
rect 2679 2433 2680 2558
rect 2531 2033 2532 2436
rect 2691 2435 2692 2558
rect 2547 2437 2548 2558
rect 3054 2437 3055 2558
rect 2549 2033 2550 2440
rect 2709 2439 2710 2558
rect 2555 2033 2556 2442
rect 3024 2441 3025 2558
rect 2559 2443 2560 2558
rect 3128 2443 3129 2558
rect 2585 2033 2586 2446
rect 2751 2445 2752 2558
rect 2591 2033 2592 2448
rect 2769 2447 2770 2558
rect 2603 2033 2604 2450
rect 2775 2449 2776 2558
rect 2619 2451 2620 2558
rect 3064 2451 3065 2558
rect 2625 2453 2626 2558
rect 3061 2453 3062 2558
rect 2627 2033 2628 2456
rect 2793 2455 2794 2558
rect 2630 2033 2631 2458
rect 2796 2457 2797 2558
rect 2631 2459 2632 2558
rect 2900 2033 2901 2460
rect 2637 2461 2638 2558
rect 3121 2461 3122 2558
rect 2643 2463 2644 2558
rect 3107 2463 3108 2558
rect 2649 2465 2650 2558
rect 3104 2465 3105 2558
rect 2651 2033 2652 2468
rect 2823 2467 2824 2558
rect 2654 2033 2655 2470
rect 2925 2033 2926 2470
rect 2501 2033 2502 2472
rect 2655 2471 2656 2558
rect 2667 2471 2668 2558
rect 2897 2033 2898 2472
rect 2675 2033 2676 2474
rect 2835 2473 2836 2558
rect 2685 2475 2686 2558
rect 3111 2475 3112 2558
rect 2696 2033 2697 2478
rect 2886 2477 2887 2558
rect 2537 2033 2538 2480
rect 2697 2479 2698 2558
rect 2720 2033 2721 2480
rect 2898 2479 2899 2558
rect 2561 2033 2562 2482
rect 2721 2481 2722 2558
rect 2726 2033 2727 2482
rect 2904 2481 2905 2558
rect 2727 2483 2728 2558
rect 3027 2483 3028 2558
rect 2733 2485 2734 2558
rect 2867 2033 2868 2486
rect 2741 2033 2742 2488
rect 2868 2487 2869 2558
rect 2756 2033 2757 2490
rect 2946 2489 2947 2558
rect 2757 2491 2758 2558
rect 2907 2033 2908 2492
rect 2762 2033 2763 2494
rect 2952 2493 2953 2558
rect 2597 2033 2598 2496
rect 2763 2495 2764 2558
rect 2781 2033 2782 2496
rect 2970 2495 2971 2558
rect 2609 2033 2610 2498
rect 2781 2497 2782 2558
rect 2787 2033 2788 2498
rect 2982 2497 2983 2558
rect 2615 2033 2616 2500
rect 2787 2499 2788 2558
rect 2799 2033 2800 2500
rect 2988 2499 2989 2558
rect 1439 2501 1440 2558
rect 2799 2501 2800 2558
rect 2805 2501 2806 2558
rect 3125 2501 3126 2558
rect 2811 2033 2812 2504
rect 3000 2503 3001 2558
rect 2811 2505 2812 2558
rect 2964 2505 2965 2558
rect 2814 2033 2815 2508
rect 3003 2507 3004 2558
rect 2817 2033 2818 2510
rect 3006 2509 3007 2558
rect 2820 2033 2821 2512
rect 3009 2511 3010 2558
rect 2826 2513 2827 2558
rect 2928 2033 2929 2514
rect 2738 2033 2739 2516
rect 2928 2515 2929 2558
rect 2573 2033 2574 2518
rect 2739 2517 2740 2558
rect 2830 2033 2831 2518
rect 2919 2517 2920 2558
rect 2657 2033 2658 2520
rect 2829 2519 2830 2558
rect 2833 2033 2834 2520
rect 3021 2519 3022 2558
rect 2843 2033 2844 2522
rect 3030 2521 3031 2558
rect 2847 2523 2848 2558
rect 3100 2523 3101 2558
rect 2849 2033 2850 2526
rect 3036 2525 3037 2558
rect 2853 2527 2854 2558
rect 3097 2527 3098 2558
rect 2861 2033 2862 2530
rect 3048 2529 3049 2558
rect 2864 2033 2865 2532
rect 3051 2531 3052 2558
rect 2693 2033 2694 2534
rect 2865 2533 2866 2558
rect 2873 2033 2874 2534
rect 3079 2533 3080 2558
rect 2702 2033 2703 2536
rect 2874 2535 2875 2558
rect 2543 2033 2544 2538
rect 2703 2537 2704 2558
rect 2879 2033 2880 2538
rect 3076 2537 3077 2558
rect 2744 2033 2745 2540
rect 2880 2539 2881 2558
rect 2579 2033 2580 2542
rect 2745 2541 2746 2558
rect 2891 2033 2892 2542
rect 3091 2541 3092 2558
rect 2714 2033 2715 2544
rect 2892 2543 2893 2558
rect 2621 2033 2622 2546
rect 2715 2545 2716 2558
rect 2894 2033 2895 2546
rect 3094 2545 3095 2558
rect 2911 2033 2912 2548
rect 2943 2547 2944 2558
rect 2882 2033 2883 2550
rect 2910 2549 2911 2558
rect 2747 2033 2748 2552
rect 2883 2551 2884 2558
rect 2914 2033 2915 2552
rect 2940 2551 2941 2558
rect 2921 2033 2922 2554
rect 3073 2553 3074 2558
rect 2765 2033 2766 2556
rect 2922 2555 2923 2558
rect 1420 2564 1421 3127
rect 2259 2562 2260 2565
rect 1434 2566 1435 3127
rect 1604 2566 1605 3127
rect 1436 2562 1437 2569
rect 2151 2562 2152 2569
rect 1439 2562 1440 2571
rect 2319 2562 2320 2571
rect 1441 2572 1442 3127
rect 2177 2572 2178 3127
rect 1443 2562 1444 2575
rect 2307 2562 2308 2575
rect 1450 2562 1451 2577
rect 1773 2562 1774 2577
rect 1438 2578 1439 3127
rect 1450 2578 1451 3127
rect 1457 2562 1458 2579
rect 1947 2562 1948 2579
rect 1456 2580 1457 3127
rect 1641 2562 1642 2581
rect 1464 2562 1465 2583
rect 2181 2562 2182 2583
rect 1463 2584 1464 3127
rect 2322 2562 2323 2585
rect 1474 2562 1475 2587
rect 2115 2562 2116 2587
rect 1473 2588 1474 3127
rect 1863 2562 1864 2589
rect 1486 2562 1487 2591
rect 2793 2562 2794 2591
rect 1488 2592 1489 3127
rect 1923 2562 1924 2593
rect 1427 2594 1428 3127
rect 1922 2594 1923 3127
rect 1490 2562 1491 2597
rect 1839 2562 1840 2597
rect 1491 2598 1492 3127
rect 2049 2562 2050 2599
rect 1493 2562 1494 2601
rect 2858 2600 2859 3127
rect 1497 2562 1498 2603
rect 1593 2562 1594 2603
rect 1498 2604 1499 3127
rect 2048 2604 2049 3127
rect 1500 2562 1501 2607
rect 2400 2562 2401 2607
rect 1514 2608 1515 3127
rect 1515 2562 1516 2609
rect 1521 2562 1522 2609
rect 3114 2562 3115 2609
rect 1526 2610 1527 3127
rect 1545 2562 1546 2611
rect 1533 2562 1534 2613
rect 1538 2612 1539 3127
rect 1569 2562 1570 2613
rect 1580 2612 1581 3127
rect 1568 2614 1569 3127
rect 1575 2562 1576 2615
rect 1563 2562 1564 2617
rect 1574 2616 1575 3127
rect 1551 2562 1552 2619
rect 1562 2618 1563 3127
rect 1550 2620 1551 3127
rect 1557 2562 1558 2621
rect 1417 2622 1418 3127
rect 1556 2622 1557 3127
rect 1587 2562 1588 2623
rect 1592 2622 1593 3127
rect 1601 2622 1602 3127
rect 2984 2622 2985 3127
rect 1611 2562 1612 2625
rect 2441 2624 2442 3127
rect 1616 2626 1617 3127
rect 3164 2626 3165 3127
rect 1629 2562 1630 2629
rect 1634 2628 1635 3127
rect 1677 2562 1678 2629
rect 1766 2628 1767 3127
rect 1676 2630 1677 3127
rect 1683 2562 1684 2631
rect 1665 2562 1666 2633
rect 1682 2632 1683 3127
rect 1653 2562 1654 2635
rect 1664 2634 1665 3127
rect 1623 2562 1624 2637
rect 1652 2636 1653 3127
rect 1689 2562 1690 2637
rect 3030 2562 3031 2637
rect 1688 2638 1689 3127
rect 1719 2562 1720 2639
rect 1695 2562 1696 2641
rect 1712 2640 1713 3127
rect 1694 2642 1695 3127
rect 1725 2562 1726 2643
rect 1701 2562 1702 2645
rect 1724 2644 1725 3127
rect 1707 2562 1708 2647
rect 1730 2646 1731 3127
rect 1706 2648 1707 3127
rect 1737 2562 1738 2649
rect 1718 2650 1719 3127
rect 1749 2562 1750 2651
rect 1736 2652 1737 3127
rect 1743 2562 1744 2653
rect 1453 2562 1454 2655
rect 1742 2654 1743 3127
rect 1748 2654 1749 3127
rect 1779 2562 1780 2655
rect 1754 2656 1755 3127
rect 1785 2562 1786 2657
rect 1761 2562 1762 2659
rect 2990 2658 2991 3127
rect 1671 2562 1672 2661
rect 1760 2660 1761 3127
rect 1659 2562 1660 2663
rect 1670 2662 1671 3127
rect 1647 2562 1648 2665
rect 1658 2664 1659 3127
rect 1772 2664 1773 3127
rect 1833 2562 1834 2665
rect 1784 2666 1785 3127
rect 1845 2562 1846 2667
rect 1797 2562 1798 2669
rect 2912 2668 2913 3127
rect 1796 2670 1797 3127
rect 1857 2562 1858 2671
rect 1832 2672 1833 3127
rect 1851 2562 1852 2673
rect 1838 2674 1839 3127
rect 1875 2562 1876 2675
rect 1844 2676 1845 3127
rect 1971 2562 1972 2677
rect 1850 2678 1851 3127
rect 1881 2562 1882 2679
rect 1856 2680 1857 3127
rect 1899 2562 1900 2681
rect 1862 2682 1863 3127
rect 1977 2562 1978 2683
rect 1880 2684 1881 3127
rect 1893 2562 1894 2685
rect 1887 2562 1888 2687
rect 3155 2686 3156 3127
rect 1886 2688 1887 3127
rect 1929 2562 1930 2689
rect 1424 2690 1425 3127
rect 1928 2690 1929 3127
rect 1892 2692 1893 3127
rect 1905 2562 1906 2693
rect 1898 2694 1899 3127
rect 1935 2562 1936 2695
rect 1904 2696 1905 3127
rect 1941 2562 1942 2697
rect 1911 2562 1912 2699
rect 2964 2562 2965 2699
rect 1910 2700 1911 3127
rect 1953 2562 1954 2701
rect 1916 2702 1917 3127
rect 1959 2562 1960 2703
rect 1934 2704 1935 3127
rect 1965 2562 1966 2705
rect 1940 2706 1941 3127
rect 3027 2562 3028 2707
rect 1946 2708 1947 3127
rect 1995 2562 1996 2709
rect 1952 2710 1953 3127
rect 1983 2562 1984 2711
rect 1958 2712 1959 3127
rect 1989 2562 1990 2713
rect 1964 2714 1965 3127
rect 3024 2562 3025 2715
rect 1970 2716 1971 3127
rect 3015 2562 3016 2717
rect 1976 2718 1977 3127
rect 2007 2562 2008 2719
rect 1982 2720 1983 3127
rect 2001 2562 2002 2721
rect 1988 2722 1989 3127
rect 3107 2562 3108 2723
rect 1994 2724 1995 3127
rect 2031 2562 2032 2725
rect 2000 2726 2001 3127
rect 2025 2562 2026 2727
rect 2006 2728 2007 3127
rect 2037 2562 2038 2729
rect 2019 2562 2020 2731
rect 2792 2730 2793 3127
rect 2018 2732 2019 3127
rect 2043 2562 2044 2733
rect 2024 2734 2025 3127
rect 2055 2562 2056 2735
rect 2030 2736 2031 3127
rect 2085 2562 2086 2737
rect 2036 2738 2037 3127
rect 2067 2562 2068 2739
rect 2042 2740 2043 3127
rect 2079 2562 2080 2741
rect 1483 2562 1484 2743
rect 2078 2742 2079 3127
rect 1446 2562 1447 2745
rect 1482 2744 1483 3127
rect 2054 2744 2055 3127
rect 3226 2744 3227 3127
rect 2061 2562 2062 2747
rect 2930 2746 2931 3127
rect 2060 2748 2061 3127
rect 2073 2562 2074 2749
rect 1432 2562 1433 2751
rect 2072 2750 2073 3127
rect 1431 2752 1432 3127
rect 1599 2562 1600 2753
rect 1598 2754 1599 3127
rect 2943 2562 2944 2755
rect 2084 2756 2085 3127
rect 2103 2562 2104 2757
rect 2097 2562 2098 2759
rect 2102 2758 2103 3127
rect 2091 2562 2092 2761
rect 2096 2760 2097 3127
rect 2090 2762 2091 3127
rect 2109 2562 2110 2763
rect 1471 2562 1472 2765
rect 2108 2764 2109 3127
rect 1470 2766 1471 3127
rect 2066 2766 2067 3127
rect 2114 2766 2115 3127
rect 2121 2562 2122 2767
rect 2120 2768 2121 3127
rect 2127 2562 2128 2769
rect 1495 2770 1496 3127
rect 2126 2770 2127 3127
rect 2144 2770 2145 3127
rect 2145 2562 2146 2771
rect 2150 2770 2151 3127
rect 2157 2562 2158 2771
rect 2156 2772 2157 3127
rect 2163 2562 2164 2773
rect 2162 2774 2163 3127
rect 2205 2562 2206 2775
rect 2174 2776 2175 3127
rect 2175 2562 2176 2777
rect 2180 2776 2181 3127
rect 2199 2562 2200 2777
rect 2187 2562 2188 2779
rect 2222 2778 2223 3127
rect 2186 2780 2187 3127
rect 3152 2780 3153 3127
rect 2196 2562 2197 2783
rect 2231 2782 2232 3127
rect 2198 2784 2199 3127
rect 2217 2562 2218 2785
rect 2204 2786 2205 3127
rect 2253 2562 2254 2787
rect 2216 2788 2217 3127
rect 3185 2788 3186 3127
rect 2229 2562 2230 2791
rect 2258 2790 2259 3127
rect 2193 2562 2194 2793
rect 2228 2792 2229 3127
rect 2192 2794 2193 3127
rect 3107 2794 3108 3127
rect 2241 2562 2242 2797
rect 2967 2562 2968 2797
rect 2240 2798 2241 3127
rect 2553 2562 2554 2799
rect 2250 2562 2251 2801
rect 2285 2800 2286 3127
rect 2252 2802 2253 3127
rect 2547 2562 2548 2803
rect 2271 2562 2272 2805
rect 2306 2804 2307 3127
rect 2270 2806 2271 3127
rect 2577 2562 2578 2807
rect 2295 2562 2296 2809
rect 2318 2808 2319 3127
rect 2294 2810 2295 3127
rect 2325 2562 2326 2811
rect 2301 2562 2302 2813
rect 2324 2812 2325 3127
rect 2316 2562 2317 2815
rect 2351 2814 2352 3127
rect 2364 2562 2365 2815
rect 2876 2814 2877 3127
rect 2334 2562 2335 2817
rect 2363 2816 2364 3127
rect 2310 2562 2311 2819
rect 2333 2818 2334 3127
rect 2370 2562 2371 2819
rect 2405 2818 2406 3127
rect 2376 2562 2377 2821
rect 2387 2820 2388 3127
rect 2340 2562 2341 2823
rect 2375 2822 2376 3127
rect 2436 2562 2437 2823
rect 2495 2822 2496 3127
rect 2451 2562 2452 2825
rect 2919 2562 2920 2825
rect 2409 2562 2410 2827
rect 2450 2826 2451 3127
rect 2403 2562 2404 2829
rect 2408 2828 2409 3127
rect 2367 2562 2368 2831
rect 2402 2830 2403 3127
rect 2460 2562 2461 2831
rect 2501 2830 2502 3127
rect 2493 2562 2494 2833
rect 2552 2832 2553 3127
rect 2433 2562 2434 2835
rect 2492 2834 2493 3127
rect 1429 2562 1430 2837
rect 2432 2836 2433 3127
rect 2499 2562 2500 2837
rect 2546 2836 2547 3127
rect 2457 2562 2458 2839
rect 2498 2838 2499 3127
rect 2415 2562 2416 2841
rect 2456 2840 2457 3127
rect 2379 2562 2380 2843
rect 2414 2842 2415 3127
rect 2378 2844 2379 3127
rect 2385 2562 2386 2845
rect 2373 2562 2374 2847
rect 2384 2846 2385 3127
rect 2337 2562 2338 2849
rect 2372 2848 2373 3127
rect 2289 2562 2290 2851
rect 2336 2850 2337 3127
rect 2529 2562 2530 2851
rect 2576 2850 2577 3127
rect 2481 2562 2482 2853
rect 2528 2852 2529 3127
rect 2439 2562 2440 2855
rect 2480 2854 2481 3127
rect 2397 2562 2398 2857
rect 2438 2856 2439 3127
rect 2361 2562 2362 2859
rect 2396 2858 2397 3127
rect 2331 2562 2332 2861
rect 2360 2860 2361 3127
rect 2283 2562 2284 2863
rect 2330 2862 2331 3127
rect 2247 2562 2248 2865
rect 2282 2864 2283 3127
rect 2246 2866 2247 3127
rect 2517 2562 2518 2867
rect 2475 2562 2476 2869
rect 2516 2868 2517 3127
rect 2474 2870 2475 3127
rect 2916 2562 2917 2871
rect 2613 2562 2614 2873
rect 3061 2562 3062 2873
rect 2601 2562 2602 2875
rect 2612 2874 2613 3127
rect 2571 2562 2572 2877
rect 2600 2876 2601 3127
rect 2523 2562 2524 2879
rect 2570 2878 2571 3127
rect 1586 2880 1587 3127
rect 2522 2880 2523 3127
rect 2655 2562 2656 2881
rect 3229 2880 3230 3127
rect 2595 2562 2596 2883
rect 2654 2882 2655 3127
rect 2594 2884 2595 3127
rect 3189 2884 3190 3127
rect 2745 2562 2746 2887
rect 2816 2886 2817 3127
rect 2691 2562 2692 2889
rect 2744 2888 2745 3127
rect 2631 2562 2632 2891
rect 2690 2890 2691 3127
rect 2787 2562 2788 2891
rect 3240 2890 3241 3127
rect 2721 2562 2722 2893
rect 2786 2892 2787 3127
rect 2667 2562 2668 2895
rect 2720 2894 2721 3127
rect 2666 2896 2667 3127
rect 3064 2562 3065 2897
rect 2796 2562 2797 2899
rect 2888 2898 2889 3127
rect 2805 2562 2806 2901
rect 2936 2900 2937 3127
rect 2739 2562 2740 2903
rect 2804 2902 2805 3127
rect 2685 2562 2686 2905
rect 2738 2904 2739 3127
rect 2211 2562 2212 2907
rect 2684 2906 2685 3127
rect 2210 2908 2211 3127
rect 2349 2562 2350 2909
rect 2313 2562 2314 2911
rect 2348 2910 2349 3127
rect 2277 2562 2278 2913
rect 2312 2912 2313 3127
rect 2276 2914 2277 3127
rect 2511 2562 2512 2915
rect 2487 2562 2488 2917
rect 2510 2916 2511 3127
rect 2445 2562 2446 2919
rect 2486 2918 2487 3127
rect 1692 2562 1693 2921
rect 2444 2920 2445 3127
rect 2811 2562 2812 2921
rect 2942 2920 2943 3127
rect 1505 2922 1506 3127
rect 2810 2922 2811 3127
rect 2826 2562 2827 2923
rect 2906 2922 2907 3127
rect 2829 2562 2830 2925
rect 2918 2924 2919 3127
rect 2763 2562 2764 2927
rect 2828 2926 2829 3127
rect 2762 2928 2763 3127
rect 3247 2928 3248 3127
rect 2835 2562 2836 2931
rect 3026 2930 3027 3127
rect 2757 2562 2758 2933
rect 2834 2932 2835 3127
rect 2697 2562 2698 2935
rect 2756 2934 2757 3127
rect 2643 2562 2644 2937
rect 2696 2936 2697 3127
rect 2642 2938 2643 3127
rect 3233 2938 3234 3127
rect 2841 2562 2842 2941
rect 3097 2562 3098 2941
rect 2775 2562 2776 2943
rect 2840 2942 2841 3127
rect 2709 2562 2710 2945
rect 2774 2944 2775 3127
rect 2637 2562 2638 2947
rect 2708 2946 2709 3127
rect 2636 2948 2637 3127
rect 2894 2948 2895 3127
rect 2847 2562 2848 2951
rect 2954 2950 2955 3127
rect 2781 2562 2782 2953
rect 2846 2952 2847 3127
rect 2727 2562 2728 2955
rect 2780 2954 2781 3127
rect 2673 2562 2674 2957
rect 2726 2956 2727 3127
rect 2619 2562 2620 2959
rect 2672 2958 2673 3127
rect 2618 2960 2619 3127
rect 3219 2960 3220 3127
rect 2853 2562 2854 2963
rect 2948 2962 2949 3127
rect 2769 2562 2770 2965
rect 2852 2964 2853 3127
rect 2703 2562 2704 2967
rect 2768 2966 2769 3127
rect 2649 2562 2650 2969
rect 2702 2968 2703 3127
rect 2589 2562 2590 2971
rect 2648 2970 2649 3127
rect 2588 2972 2589 3127
rect 3192 2972 3193 3127
rect 2865 2562 2866 2975
rect 2960 2974 2961 3127
rect 2799 2562 2800 2977
rect 2864 2976 2865 3127
rect 2733 2562 2734 2979
rect 2798 2978 2799 3127
rect 2133 2562 2134 2981
rect 2732 2980 2733 3127
rect 2132 2982 2133 3127
rect 2139 2562 2140 2983
rect 2138 2984 2139 3127
rect 2169 2562 2170 2985
rect 1467 2562 1468 2987
rect 2168 2986 2169 3127
rect 1466 2988 1467 3127
rect 1640 2988 1641 3127
rect 2868 2562 2869 2989
rect 2966 2988 2967 3127
rect 2870 2990 2871 3127
rect 3222 2990 3223 3127
rect 2883 2562 2884 2993
rect 3059 2992 3060 3127
rect 2886 2562 2887 2995
rect 3032 2994 3033 3127
rect 2898 2562 2899 2997
rect 3014 2996 3015 3127
rect 2910 2562 2911 2999
rect 3057 2562 3058 2999
rect 2823 2562 2824 3001
rect 2909 3000 2910 3127
rect 2751 2562 2752 3003
rect 2822 3002 2823 3127
rect 2679 2562 2680 3005
rect 2750 3004 2751 3127
rect 2625 2562 2626 3007
rect 2678 3006 2679 3127
rect 2583 2562 2584 3009
rect 2624 3008 2625 3127
rect 2535 2562 2536 3011
rect 2582 3010 2583 3127
rect 2534 3012 2535 3127
rect 2897 3012 2898 3127
rect 2880 2562 2881 3015
rect 3056 3014 3057 3127
rect 1803 2562 1804 3017
rect 2879 3016 2880 3127
rect 1802 3018 1803 3127
rect 1815 2562 1816 3019
rect 1502 3020 1503 3127
rect 1814 3020 1815 3127
rect 2924 3020 2925 3127
rect 3125 2562 3126 3021
rect 2928 2562 2929 3023
rect 3071 3022 3072 3127
rect 2940 2562 2941 3025
rect 3068 3024 3069 3127
rect 2946 2562 2947 3027
rect 3086 3026 3087 3127
rect 2963 3028 2964 3127
rect 3118 2562 3119 3029
rect 2972 3030 2973 3127
rect 3100 2562 3101 3031
rect 2996 3032 2997 3127
rect 3243 3032 3244 3127
rect 3000 2562 3001 3035
rect 3140 3034 3141 3127
rect 3003 2562 3004 3037
rect 3143 3036 3144 3127
rect 2508 2562 2509 3039
rect 3002 3038 3003 3127
rect 3006 2562 3007 3039
rect 3146 3038 3147 3127
rect 1791 2562 1792 3041
rect 3005 3040 3006 3127
rect 1790 3042 1791 3127
rect 1809 2562 1810 3043
rect 1808 3044 1809 3127
rect 1821 2562 1822 3045
rect 1820 3046 1821 3127
rect 1827 2562 1828 3047
rect 1826 3048 1827 3127
rect 1869 2562 1870 3049
rect 1868 3050 1869 3127
rect 2013 2562 2014 3051
rect 2012 3052 2013 3127
rect 3012 2562 3013 3053
rect 3009 2562 3010 3055
rect 3149 3054 3150 3127
rect 2892 2562 2893 3057
rect 3008 3056 3009 3127
rect 2715 2562 2716 3059
rect 2891 3058 2892 3127
rect 2661 2562 2662 3061
rect 2714 3060 2715 3127
rect 2607 2562 2608 3063
rect 2660 3062 2661 3127
rect 2559 2562 2560 3065
rect 2606 3064 2607 3127
rect 2558 3066 2559 3127
rect 2565 2562 2566 3067
rect 2541 2562 2542 3069
rect 2564 3068 2565 3127
rect 2463 2562 2464 3071
rect 2540 3070 2541 3127
rect 2421 2562 2422 3073
rect 2462 3072 2463 3127
rect 1589 3074 1590 3127
rect 2420 3074 2421 3127
rect 3018 2562 3019 3075
rect 3158 3074 3159 3127
rect 3021 2562 3022 3077
rect 3161 3076 3162 3127
rect 2904 2562 2905 3079
rect 3020 3078 3021 3127
rect 3036 2562 3037 3079
rect 3179 3078 3180 3127
rect 3044 3080 3045 3127
rect 3167 3080 3168 3127
rect 3048 2562 3049 3083
rect 3054 2562 3055 3083
rect 3051 2562 3052 3085
rect 3176 3084 3177 3127
rect 2874 2562 2875 3087
rect 3050 3086 3051 3127
rect 3073 2562 3074 3087
rect 3213 3086 3214 3127
rect 2366 3088 2367 3127
rect 3074 3088 3075 3127
rect 3076 2562 3077 3089
rect 3216 3088 3217 3127
rect 2300 3090 2301 3127
rect 3077 3090 3078 3127
rect 3079 2562 3080 3091
rect 3111 2562 3112 3091
rect 2922 2562 2923 3093
rect 3080 3092 3081 3127
rect 2970 2562 2971 3095
rect 3110 3094 3111 3127
rect 3091 2562 3092 3097
rect 3201 3096 3202 3127
rect 2952 2562 2953 3099
rect 3092 3098 3093 3127
rect 3094 2562 3095 3099
rect 3204 3098 3205 3127
rect 3104 2562 3105 3101
rect 3182 3100 3183 3127
rect 2505 2562 2506 3103
rect 3104 3102 3105 3127
rect 2469 2562 2470 3105
rect 2504 3104 2505 3127
rect 2427 2562 2428 3107
rect 2468 3106 2469 3127
rect 2391 2562 2392 3109
rect 2426 3108 2427 3127
rect 2355 2562 2356 3111
rect 2390 3110 2391 3127
rect 2343 2562 2344 3113
rect 2354 3112 2355 3127
rect 2265 2562 2266 3115
rect 2342 3114 2343 3127
rect 2235 2562 2236 3117
rect 2264 3116 2265 3127
rect 1460 2562 1461 3119
rect 2234 3118 2235 3127
rect 1459 3120 1460 3127
rect 2288 3120 2289 3127
rect 3121 2562 3122 3121
rect 3236 3120 3237 3127
rect 2982 2562 2983 3123
rect 3122 3122 3123 3127
rect 3128 2562 3129 3123
rect 3250 3122 3251 3127
rect 2988 2562 2989 3125
rect 3128 3124 3129 3127
rect 1417 3131 1418 3134
rect 1922 3131 1923 3134
rect 1420 3131 1421 3136
rect 2048 3131 2049 3136
rect 1427 3131 1428 3138
rect 1916 3131 1917 3138
rect 1431 3131 1432 3140
rect 2387 3131 2388 3140
rect 1431 3141 1432 3700
rect 2156 3131 2157 3142
rect 1441 3131 1442 3144
rect 2302 3143 2303 3700
rect 1459 3131 1460 3146
rect 1946 3131 1947 3146
rect 1463 3131 1464 3148
rect 1688 3131 1689 3148
rect 1427 3149 1428 3700
rect 1687 3149 1688 3700
rect 1450 3131 1451 3152
rect 1462 3151 1463 3700
rect 1438 3131 1439 3154
rect 1450 3153 1451 3700
rect 1438 3155 1439 3700
rect 2612 3131 2613 3156
rect 1466 3131 1467 3158
rect 1904 3131 1905 3158
rect 1468 3159 1469 3700
rect 3037 3159 3038 3700
rect 1473 3131 1474 3162
rect 2060 3131 2061 3162
rect 1485 3163 1486 3700
rect 2282 3131 2283 3164
rect 1488 3131 1489 3166
rect 2222 3131 2223 3166
rect 1491 3131 1492 3168
rect 2114 3131 2115 3168
rect 1495 3131 1496 3170
rect 2042 3131 2043 3170
rect 1482 3131 1483 3172
rect 1494 3171 1495 3700
rect 1498 3131 1499 3172
rect 2036 3131 2037 3172
rect 1502 3131 1503 3174
rect 2072 3131 2073 3174
rect 1505 3131 1506 3176
rect 2012 3131 2013 3176
rect 1507 3177 1508 3700
rect 1568 3131 1569 3178
rect 1514 3131 1515 3180
rect 1519 3179 1520 3700
rect 1526 3131 1527 3180
rect 1531 3179 1532 3700
rect 1525 3181 1526 3700
rect 1616 3131 1617 3182
rect 1528 3183 1529 3700
rect 2501 3131 2502 3184
rect 1538 3131 1539 3186
rect 1543 3185 1544 3700
rect 1562 3131 1563 3186
rect 1567 3185 1568 3700
rect 1556 3131 1557 3188
rect 1561 3187 1562 3700
rect 1478 3189 1479 3700
rect 1555 3189 1556 3700
rect 1586 3131 1587 3190
rect 2024 3131 2025 3190
rect 1580 3131 1581 3192
rect 1585 3191 1586 3700
rect 1574 3131 1575 3194
rect 1579 3193 1580 3700
rect 1475 3195 1476 3700
rect 1573 3195 1574 3700
rect 1592 3131 1593 3196
rect 1615 3195 1616 3700
rect 1601 3131 1602 3198
rect 1604 3131 1605 3198
rect 1434 3131 1435 3200
rect 1603 3199 1604 3700
rect 1434 3201 1435 3700
rect 1612 3201 1613 3700
rect 1609 3203 1610 3700
rect 3044 3131 3045 3204
rect 1633 3205 1634 3700
rect 1634 3131 1635 3206
rect 1639 3205 1640 3700
rect 1640 3131 1641 3206
rect 1658 3131 1659 3206
rect 3074 3131 3075 3206
rect 1652 3131 1653 3208
rect 1657 3207 1658 3700
rect 1663 3207 1664 3700
rect 1664 3131 1665 3208
rect 1669 3207 1670 3700
rect 1670 3131 1671 3208
rect 1675 3207 1676 3700
rect 1676 3131 1677 3208
rect 1681 3207 1682 3700
rect 1682 3131 1683 3208
rect 1694 3131 1695 3208
rect 1699 3207 1700 3700
rect 1712 3131 1713 3208
rect 3243 3131 3244 3208
rect 1706 3131 1707 3210
rect 1711 3209 1712 3700
rect 1717 3209 1718 3700
rect 1718 3131 1719 3210
rect 1724 3131 1725 3210
rect 2422 3209 2423 3700
rect 1723 3211 1724 3700
rect 3247 3131 3248 3212
rect 1748 3131 1749 3214
rect 1777 3213 1778 3700
rect 1736 3131 1737 3216
rect 1747 3215 1748 3700
rect 1753 3215 1754 3700
rect 1754 3131 1755 3216
rect 1759 3215 1760 3700
rect 1760 3131 1761 3216
rect 1765 3215 1766 3700
rect 1766 3131 1767 3216
rect 1844 3131 1845 3216
rect 1921 3215 1922 3700
rect 1802 3131 1803 3218
rect 1843 3217 1844 3700
rect 1772 3131 1773 3220
rect 1801 3219 1802 3700
rect 1742 3131 1743 3222
rect 1771 3221 1772 3700
rect 1730 3131 1731 3224
rect 1741 3223 1742 3700
rect 1424 3131 1425 3226
rect 1729 3225 1730 3700
rect 1424 3227 1425 3700
rect 1693 3227 1694 3700
rect 1862 3131 1863 3228
rect 3152 3131 3153 3228
rect 1820 3131 1821 3230
rect 1861 3229 1862 3700
rect 1819 3231 1820 3700
rect 1826 3131 1827 3232
rect 1825 3233 1826 3700
rect 1832 3131 1833 3234
rect 1796 3131 1797 3236
rect 1831 3235 1832 3700
rect 1795 3237 1796 3700
rect 1850 3131 1851 3238
rect 1790 3131 1791 3240
rect 1849 3239 1850 3700
rect 1789 3241 1790 3700
rect 1808 3131 1809 3242
rect 1807 3243 1808 3700
rect 1838 3131 1839 3244
rect 1837 3245 1838 3700
rect 1856 3131 1857 3246
rect 1873 3245 1874 3700
rect 1880 3131 1881 3246
rect 1879 3247 1880 3700
rect 1892 3131 1893 3248
rect 1868 3131 1869 3250
rect 1891 3249 1892 3700
rect 1814 3131 1815 3252
rect 1867 3251 1868 3700
rect 1784 3131 1785 3254
rect 1813 3253 1814 3700
rect 1903 3253 1904 3700
rect 1928 3131 1929 3254
rect 1915 3255 1916 3700
rect 2792 3131 2793 3256
rect 1927 3257 1928 3700
rect 1952 3131 1953 3258
rect 1621 3259 1622 3700
rect 1951 3259 1952 3700
rect 1945 3261 1946 3700
rect 1976 3131 1977 3262
rect 1975 3263 1976 3700
rect 2000 3131 2001 3264
rect 1999 3265 2000 3700
rect 2030 3131 2031 3266
rect 1482 3267 1483 3700
rect 2029 3267 2030 3700
rect 2011 3269 2012 3700
rect 2066 3131 2067 3270
rect 2023 3271 2024 3700
rect 2090 3131 2091 3272
rect 2035 3273 2036 3700
rect 2096 3131 2097 3274
rect 2041 3275 2042 3700
rect 2102 3131 2103 3276
rect 2047 3277 2048 3700
rect 2078 3131 2079 3278
rect 2054 3131 2055 3280
rect 2065 3279 2066 3700
rect 2053 3281 2054 3700
rect 2108 3131 2109 3282
rect 2059 3283 2060 3700
rect 2120 3131 2121 3284
rect 2071 3285 2072 3700
rect 2138 3131 2139 3286
rect 2080 3287 2081 3700
rect 2879 3131 2880 3288
rect 2089 3289 2090 3700
rect 2150 3131 2151 3290
rect 2095 3291 2096 3700
rect 2180 3131 2181 3292
rect 2101 3293 2102 3700
rect 2186 3131 2187 3294
rect 2107 3295 2108 3700
rect 2174 3131 2175 3296
rect 2113 3297 2114 3700
rect 2162 3131 2163 3298
rect 1598 3131 1599 3300
rect 2161 3299 2162 3700
rect 1510 3301 1511 3700
rect 1597 3301 1598 3700
rect 2119 3301 2120 3700
rect 2666 3131 2667 3302
rect 2132 3131 2133 3304
rect 3155 3131 3156 3304
rect 2131 3305 2132 3700
rect 2210 3131 2211 3306
rect 2137 3307 2138 3700
rect 2270 3131 2271 3308
rect 2149 3309 2150 3700
rect 2216 3131 2217 3310
rect 2155 3311 2156 3700
rect 2252 3131 2253 3312
rect 2173 3313 2174 3700
rect 2228 3131 2229 3314
rect 1456 3131 1457 3316
rect 2227 3315 2228 3700
rect 1456 3317 1457 3700
rect 2177 3131 2178 3318
rect 2176 3319 2177 3700
rect 2231 3131 2232 3320
rect 2179 3321 2180 3700
rect 2234 3131 2235 3322
rect 2185 3323 2186 3700
rect 2588 3131 2589 3324
rect 2194 3325 2195 3700
rect 2285 3131 2286 3326
rect 2204 3131 2205 3328
rect 3136 3327 3137 3700
rect 2203 3329 2204 3700
rect 2264 3131 2265 3330
rect 2206 3331 2207 3700
rect 2351 3131 2352 3332
rect 2209 3333 2210 3700
rect 2258 3131 2259 3334
rect 2215 3335 2216 3700
rect 2600 3131 2601 3336
rect 2221 3337 2222 3700
rect 2564 3131 2565 3338
rect 2233 3339 2234 3700
rect 2288 3131 2289 3340
rect 2240 3131 2241 3342
rect 3189 3131 3190 3342
rect 2239 3343 2240 3700
rect 2660 3131 2661 3344
rect 2198 3131 2199 3346
rect 2659 3345 2660 3700
rect 2197 3347 2198 3700
rect 2594 3131 2595 3348
rect 2251 3349 2252 3700
rect 2342 3131 2343 3350
rect 2257 3351 2258 3700
rect 2300 3131 2301 3352
rect 1441 3353 1442 3700
rect 2299 3353 2300 3700
rect 2263 3355 2264 3700
rect 2366 3131 2367 3356
rect 2269 3357 2270 3700
rect 2306 3131 2307 3358
rect 2276 3131 2277 3360
rect 3077 3131 3078 3360
rect 1886 3131 1887 3362
rect 3076 3361 3077 3700
rect 1885 3363 1886 3700
rect 1898 3131 1899 3364
rect 1897 3365 1898 3700
rect 1910 3131 1911 3366
rect 1909 3367 1910 3700
rect 1934 3131 1935 3368
rect 1933 3369 1934 3700
rect 1958 3131 1959 3370
rect 1957 3371 1958 3700
rect 1982 3131 1983 3372
rect 1589 3131 1590 3374
rect 1981 3373 1982 3700
rect 2275 3373 2276 3700
rect 2312 3131 2313 3374
rect 2281 3375 2282 3700
rect 2330 3131 2331 3376
rect 2284 3377 2285 3700
rect 2333 3131 2334 3378
rect 2287 3379 2288 3700
rect 2336 3131 2337 3380
rect 2305 3381 2306 3700
rect 2534 3131 2535 3382
rect 2311 3383 2312 3700
rect 2897 3131 2898 3384
rect 2324 3131 2325 3386
rect 2329 3385 2330 3700
rect 2192 3131 2193 3388
rect 2323 3387 2324 3700
rect 1417 3389 1418 3700
rect 2191 3389 2192 3700
rect 2335 3389 2336 3700
rect 2546 3131 2547 3390
rect 2341 3391 2342 3700
rect 2384 3131 2385 3392
rect 2354 3131 2355 3394
rect 2662 3393 2663 3700
rect 2353 3395 2354 3700
rect 2474 3131 2475 3396
rect 2365 3397 2366 3700
rect 2498 3131 2499 3398
rect 2375 3131 2376 3400
rect 2410 3399 2411 3700
rect 2363 3131 2364 3402
rect 2374 3401 2375 3700
rect 2383 3401 2384 3700
rect 2690 3131 2691 3402
rect 2396 3131 2397 3404
rect 2894 3131 2895 3404
rect 2395 3405 2396 3700
rect 2480 3131 2481 3406
rect 2434 3407 2435 3700
rect 2495 3131 2496 3408
rect 2441 3131 2442 3410
rect 2446 3409 2447 3700
rect 2405 3131 2406 3412
rect 2440 3411 2441 3700
rect 1550 3131 1551 3414
rect 2404 3413 2405 3700
rect 2468 3131 2469 3414
rect 2497 3413 2498 3700
rect 2432 3131 2433 3416
rect 2467 3415 2468 3700
rect 2420 3131 2421 3418
rect 2431 3417 2432 3700
rect 2414 3131 2415 3420
rect 2419 3419 2420 3700
rect 2413 3421 2414 3700
rect 2510 3131 2511 3422
rect 2470 3423 2471 3700
rect 2876 3131 2877 3424
rect 2473 3425 2474 3700
rect 2570 3131 2571 3426
rect 2479 3427 2480 3700
rect 2696 3131 2697 3428
rect 2126 3131 2127 3430
rect 2695 3429 2696 3700
rect 2125 3431 2126 3700
rect 2672 3131 2673 3432
rect 2504 3131 2505 3434
rect 3185 3131 3186 3434
rect 2486 3131 2487 3436
rect 2503 3435 2504 3700
rect 2450 3131 2451 3438
rect 2485 3437 2486 3700
rect 2444 3131 2445 3440
rect 2449 3439 2450 3700
rect 2438 3131 2439 3442
rect 2443 3441 2444 3700
rect 2402 3131 2403 3444
rect 2437 3443 2438 3700
rect 1500 3445 1501 3700
rect 2401 3445 2402 3700
rect 2509 3445 2510 3700
rect 3182 3131 3183 3446
rect 2528 3131 2529 3448
rect 2545 3447 2546 3700
rect 2527 3449 2528 3700
rect 2654 3131 2655 3450
rect 2533 3451 2534 3700
rect 2576 3131 2577 3452
rect 2552 3131 2553 3454
rect 3104 3131 3105 3454
rect 2551 3455 2552 3700
rect 2582 3131 2583 3456
rect 2558 3131 2559 3458
rect 3192 3131 3193 3458
rect 2557 3459 2558 3700
rect 3107 3131 3108 3460
rect 2563 3461 2564 3700
rect 2606 3131 2607 3462
rect 2569 3463 2570 3700
rect 3198 3463 3199 3700
rect 2575 3465 2576 3700
rect 3195 3465 3196 3700
rect 2581 3467 2582 3700
rect 2648 3131 2649 3468
rect 2587 3469 2588 3700
rect 2624 3131 2625 3470
rect 2599 3471 2600 3700
rect 2963 3131 2964 3472
rect 2605 3473 2606 3700
rect 2636 3131 2637 3474
rect 2611 3475 2612 3700
rect 2642 3131 2643 3476
rect 2623 3477 2624 3700
rect 3236 3131 3237 3478
rect 2629 3479 2630 3700
rect 3240 3131 3241 3480
rect 2635 3481 2636 3700
rect 2714 3131 2715 3482
rect 2647 3483 2648 3700
rect 2720 3131 2721 3484
rect 2653 3485 2654 3700
rect 2726 3131 2727 3486
rect 2665 3487 2666 3700
rect 3118 3487 3119 3700
rect 2671 3489 2672 3700
rect 2738 3131 2739 3490
rect 1970 3131 1971 3492
rect 2737 3491 2738 3700
rect 1420 3493 1421 3700
rect 1969 3493 1970 3700
rect 2684 3131 2685 3494
rect 3115 3493 3116 3700
rect 1503 3495 1504 3700
rect 2683 3495 2684 3700
rect 2689 3495 2690 3700
rect 2744 3131 2745 3496
rect 2708 3131 2709 3498
rect 3226 3131 3227 3498
rect 2707 3499 2708 3700
rect 3250 3131 3251 3500
rect 2713 3501 2714 3700
rect 2756 3131 2757 3502
rect 2719 3503 2720 3700
rect 2750 3131 2751 3504
rect 2725 3505 2726 3700
rect 2768 3131 2769 3506
rect 2731 3507 2732 3700
rect 2732 3131 2733 3508
rect 2743 3507 2744 3700
rect 2798 3131 2799 3508
rect 2749 3509 2750 3700
rect 2804 3131 2805 3510
rect 2755 3511 2756 3700
rect 3188 3511 3189 3700
rect 2767 3513 2768 3700
rect 3229 3131 3230 3514
rect 2774 3131 2775 3516
rect 3170 3515 3171 3700
rect 2773 3517 2774 3700
rect 2828 3131 2829 3518
rect 1940 3131 1941 3520
rect 2827 3519 2828 3700
rect 1624 3521 1625 3700
rect 1939 3521 1940 3700
rect 2791 3521 2792 3700
rect 2822 3131 2823 3522
rect 2797 3523 2798 3700
rect 2834 3131 2835 3524
rect 2803 3525 2804 3700
rect 3219 3131 3220 3526
rect 2641 3527 2642 3700
rect 3219 3527 3220 3700
rect 2821 3529 2822 3700
rect 2846 3131 2847 3530
rect 2833 3531 2834 3700
rect 2912 3131 2913 3532
rect 2845 3533 2846 3700
rect 2864 3131 2865 3534
rect 2852 3131 2853 3536
rect 2863 3535 2864 3700
rect 2870 3131 2871 3536
rect 2884 3535 2885 3700
rect 2869 3537 2870 3700
rect 3152 3537 3153 3700
rect 2875 3539 2876 3700
rect 2924 3131 2925 3540
rect 2881 3541 2882 3700
rect 2891 3131 2892 3542
rect 2888 3131 2889 3544
rect 3073 3543 3074 3700
rect 2887 3545 2888 3700
rect 2930 3131 2931 3546
rect 2893 3547 2894 3700
rect 2936 3131 2937 3548
rect 2905 3549 2906 3700
rect 2906 3131 2907 3550
rect 2908 3549 2909 3700
rect 2909 3131 2910 3550
rect 2911 3549 2912 3700
rect 2942 3131 2943 3550
rect 2918 3131 2919 3552
rect 3155 3551 3156 3700
rect 2917 3553 2918 3700
rect 2972 3131 2973 3554
rect 2923 3555 2924 3700
rect 3005 3131 3006 3556
rect 2935 3557 2936 3700
rect 2966 3131 2967 3558
rect 1470 3131 1471 3560
rect 2965 3559 2966 3700
rect 1471 3561 1472 3700
rect 2348 3131 2349 3562
rect 2347 3563 2348 3700
rect 2408 3131 2409 3564
rect 2372 3131 2373 3566
rect 2407 3565 2408 3700
rect 2360 3131 2361 3568
rect 2371 3567 2372 3700
rect 2359 3569 2360 3700
rect 2492 3131 2493 3570
rect 2491 3571 2492 3700
rect 2618 3131 2619 3572
rect 2617 3573 2618 3700
rect 2702 3131 2703 3574
rect 2701 3575 2702 3700
rect 2762 3131 2763 3576
rect 2761 3577 2762 3700
rect 3191 3577 3192 3700
rect 2944 3579 2945 3700
rect 2960 3131 2961 3580
rect 2948 3131 2949 3582
rect 3052 3581 3053 3700
rect 2947 3583 2948 3700
rect 2984 3131 2985 3584
rect 2971 3585 2972 3700
rect 3008 3131 3009 3586
rect 2977 3587 2978 3700
rect 3014 3131 3015 3588
rect 2983 3589 2984 3700
rect 3020 3131 3021 3590
rect 3002 3131 3003 3592
rect 3040 3591 3041 3700
rect 3001 3593 3002 3700
rect 3026 3131 3027 3594
rect 3013 3595 3014 3700
rect 3164 3131 3165 3596
rect 3019 3597 3020 3700
rect 3056 3131 3057 3598
rect 3022 3599 3023 3700
rect 3059 3131 3060 3600
rect 3034 3601 3035 3700
rect 3071 3131 3072 3602
rect 3043 3603 3044 3700
rect 3080 3131 3081 3604
rect 3050 3131 3051 3606
rect 3167 3131 3168 3606
rect 2144 3131 2145 3608
rect 3049 3607 3050 3700
rect 2143 3609 2144 3700
rect 2246 3131 2247 3610
rect 2245 3611 2246 3700
rect 2294 3131 2295 3612
rect 2293 3613 2294 3700
rect 2378 3131 2379 3614
rect 2377 3615 2378 3700
rect 2426 3131 2427 3616
rect 2390 3131 2391 3618
rect 2425 3617 2426 3700
rect 2389 3619 2390 3700
rect 3133 3619 3134 3700
rect 3055 3621 3056 3700
rect 3086 3131 3087 3622
rect 3061 3623 3062 3700
rect 3092 3131 3093 3624
rect 3079 3625 3080 3700
rect 3110 3131 3111 3626
rect 3091 3627 3092 3700
rect 3122 3131 3123 3628
rect 3097 3629 3098 3700
rect 3143 3131 3144 3630
rect 2996 3131 2997 3632
rect 3142 3631 3143 3700
rect 2995 3633 2996 3700
rect 3032 3131 3033 3634
rect 3031 3635 3032 3700
rect 3068 3131 3069 3636
rect 3109 3635 3110 3700
rect 3146 3131 3147 3636
rect 2786 3131 2787 3638
rect 3145 3637 3146 3700
rect 2785 3639 2786 3700
rect 2816 3131 2817 3640
rect 1964 3131 1965 3642
rect 2815 3641 2816 3700
rect 1963 3643 1964 3700
rect 1988 3131 1989 3644
rect 1987 3645 1988 3700
rect 1994 3131 1995 3646
rect 1993 3647 1994 3700
rect 2006 3131 2007 3648
rect 2005 3649 2006 3700
rect 2018 3131 2019 3650
rect 2017 3651 2018 3700
rect 2084 3131 2085 3652
rect 2083 3653 2084 3700
rect 2168 3131 2169 3654
rect 2167 3655 2168 3700
rect 2678 3131 2679 3656
rect 2677 3657 2678 3700
rect 3209 3657 3210 3700
rect 3112 3659 3113 3700
rect 3149 3131 3150 3660
rect 3121 3661 3122 3700
rect 3158 3131 3159 3662
rect 3124 3663 3125 3700
rect 3161 3131 3162 3664
rect 3128 3131 3129 3666
rect 3222 3131 3223 3666
rect 3127 3667 3128 3700
rect 3173 3667 3174 3700
rect 3130 3669 3131 3700
rect 3140 3131 3141 3670
rect 3139 3671 3140 3700
rect 3179 3131 3180 3672
rect 3164 3673 3165 3700
rect 3201 3131 3202 3674
rect 2318 3131 2319 3676
rect 3202 3675 3203 3700
rect 2317 3677 2318 3700
rect 2540 3131 2541 3678
rect 2522 3131 2523 3680
rect 2539 3679 2540 3700
rect 2516 3131 2517 3682
rect 2521 3681 2522 3700
rect 2515 3683 2516 3700
rect 3148 3683 3149 3700
rect 3167 3683 3168 3700
rect 3204 3131 3205 3684
rect 2593 3685 2594 3700
rect 3205 3685 3206 3700
rect 3176 3131 3177 3688
rect 3233 3131 3234 3688
rect 3182 3689 3183 3700
rect 3213 3131 3214 3690
rect 2941 3691 2942 3700
rect 3212 3691 3213 3700
rect 3185 3693 3186 3700
rect 3216 3131 3217 3694
rect 2954 3131 2955 3696
rect 3216 3695 3217 3700
rect 2953 3697 2954 3700
rect 2990 3131 2991 3698
rect 1417 3704 1418 3707
rect 1927 3704 1928 3707
rect 1434 3704 1435 3709
rect 2089 3704 2090 3709
rect 1434 3710 1435 4295
rect 1585 3704 1586 3711
rect 1438 3704 1439 3713
rect 1519 3704 1520 3713
rect 1438 3714 1439 4295
rect 1573 3704 1574 3715
rect 1450 3714 1451 4295
rect 1450 3704 1451 3715
rect 1456 3714 1457 4295
rect 1456 3704 1457 3715
rect 1462 3714 1463 4295
rect 1462 3704 1463 3715
rect 1468 3704 1469 3717
rect 2209 3704 2210 3717
rect 1475 3704 1476 3719
rect 2194 3704 2195 3719
rect 1478 3704 1479 3721
rect 1531 3704 1532 3721
rect 1485 3704 1486 3723
rect 1813 3704 1814 3723
rect 1468 3724 1469 4295
rect 1814 3724 1815 4295
rect 1485 3726 1486 4295
rect 2737 3704 2738 3727
rect 1494 3726 1495 4295
rect 1494 3704 1495 3727
rect 1503 3704 1504 3729
rect 1909 3704 1910 3729
rect 1503 3730 1504 4295
rect 1843 3704 1844 3731
rect 1507 3704 1508 3733
rect 1574 3732 1575 4295
rect 1507 3734 1508 4295
rect 1615 3704 1616 3735
rect 1510 3704 1511 3737
rect 3227 3736 3228 4295
rect 1514 3738 1515 4295
rect 3221 3738 3222 4295
rect 1517 3740 1518 4295
rect 2173 3704 2174 3741
rect 1528 3704 1529 3743
rect 3112 3704 3113 3743
rect 1543 3704 1544 3745
rect 1544 3744 1545 4295
rect 1555 3704 1556 3745
rect 1556 3744 1557 4295
rect 1561 3704 1562 3745
rect 1562 3744 1563 4295
rect 1567 3704 1568 3745
rect 1568 3744 1569 4295
rect 1579 3704 1580 3745
rect 1580 3744 1581 4295
rect 1592 3744 1593 4295
rect 1597 3704 1598 3745
rect 1598 3746 1599 4295
rect 1765 3704 1766 3747
rect 1603 3704 1604 3749
rect 1604 3748 1605 4295
rect 1612 3704 1613 3749
rect 2149 3704 2150 3749
rect 1624 3704 1625 3751
rect 2665 3704 2666 3751
rect 1628 3752 1629 4295
rect 1663 3704 1664 3753
rect 1424 3704 1425 3755
rect 1664 3754 1665 4295
rect 1417 3756 1418 4295
rect 1424 3756 1425 4295
rect 1633 3704 1634 3757
rect 2003 3756 2004 4295
rect 1639 3704 1640 3759
rect 1640 3758 1641 4295
rect 1652 3758 1653 4295
rect 2434 3704 2435 3759
rect 1675 3704 1676 3761
rect 3198 3704 3199 3761
rect 1706 3762 1707 4295
rect 1879 3704 1880 3763
rect 1717 3704 1718 3765
rect 1784 3764 1785 4295
rect 1669 3704 1670 3767
rect 1718 3766 1719 4295
rect 1670 3768 1671 4295
rect 1687 3704 1688 3769
rect 1688 3770 1689 4295
rect 1693 3704 1694 3771
rect 1529 3772 1530 4295
rect 1694 3772 1695 4295
rect 1736 3772 1737 4295
rect 1771 3704 1772 3773
rect 1482 3704 1483 3775
rect 1772 3774 1773 4295
rect 1482 3776 1483 4295
rect 2143 3704 2144 3777
rect 1844 3778 1845 4295
rect 1969 3704 1970 3779
rect 1856 3780 1857 4295
rect 1939 3704 1940 3781
rect 1871 3782 1872 4295
rect 2176 3704 2177 3783
rect 1880 3784 1881 4295
rect 1981 3704 1982 3785
rect 1910 3786 1911 4295
rect 2041 3704 2042 3787
rect 1928 3788 1929 4295
rect 2107 3704 2108 3789
rect 1940 3790 1941 4295
rect 2083 3704 2084 3791
rect 1961 3792 1962 4295
rect 2206 3704 2207 3793
rect 1970 3794 1971 4295
rect 2047 3704 2048 3795
rect 1982 3796 1983 4295
rect 2227 3704 2228 3797
rect 1609 3704 1610 3799
rect 2228 3798 2229 4295
rect 1510 3800 1511 4295
rect 1610 3800 1611 4295
rect 2027 3800 2028 4295
rect 2302 3704 2303 3801
rect 2042 3802 2043 4295
rect 2269 3704 2270 3803
rect 2051 3804 2052 4295
rect 2284 3704 2285 3805
rect 2063 3806 2064 4295
rect 2410 3704 2411 3807
rect 2078 3808 2079 4295
rect 2287 3704 2288 3809
rect 2084 3810 2085 4295
rect 2341 3704 2342 3811
rect 2090 3812 2091 4295
rect 2437 3704 2438 3813
rect 2099 3814 2100 4295
rect 2440 3704 2441 3815
rect 2105 3816 2106 4295
rect 2404 3704 2405 3817
rect 2108 3818 2109 4295
rect 2251 3704 2252 3819
rect 2059 3704 2060 3821
rect 2252 3820 2253 4295
rect 2060 3822 2061 4295
rect 2407 3704 2408 3823
rect 2137 3704 2138 3825
rect 3216 3704 3217 3825
rect 2138 3826 2139 4295
rect 2353 3704 2354 3827
rect 2144 3828 2145 4295
rect 2461 3704 2462 3829
rect 2150 3830 2151 4295
rect 2443 3704 2444 3831
rect 2174 3832 2175 4295
rect 2503 3704 2504 3833
rect 2197 3704 2198 3835
rect 2408 3834 2409 4295
rect 1500 3704 1501 3837
rect 2198 3836 2199 4295
rect 2210 3836 2211 4295
rect 2365 3704 2366 3837
rect 2131 3704 2132 3839
rect 2366 3838 2367 4295
rect 2132 3840 2133 4295
rect 2347 3704 2348 3841
rect 2215 3704 2216 3843
rect 3252 3842 3253 4295
rect 2216 3844 2217 4295
rect 2521 3704 2522 3845
rect 2101 3704 2102 3847
rect 2522 3846 2523 4295
rect 2102 3848 2103 4295
rect 2401 3704 2402 3849
rect 2185 3704 2186 3851
rect 2402 3850 2403 4295
rect 2186 3852 2187 4295
rect 2359 3704 2360 3853
rect 2257 3704 2258 3855
rect 2342 3854 2343 4295
rect 2258 3856 2259 4295
rect 2515 3704 2516 3857
rect 2167 3704 2168 3859
rect 2516 3858 2517 4295
rect 2168 3860 2169 4295
rect 2455 3704 2456 3861
rect 2263 3704 2264 3863
rect 3291 3862 3292 4295
rect 2161 3704 2162 3865
rect 2264 3864 2265 4295
rect 2162 3866 2163 4295
rect 2497 3704 2498 3867
rect 2239 3704 2240 3869
rect 2498 3868 2499 4295
rect 2240 3870 2241 4295
rect 2539 3704 2540 3871
rect 2270 3872 2271 4295
rect 2662 3704 2663 3873
rect 2288 3874 2289 4295
rect 2293 3704 2294 3875
rect 2294 3876 2295 4295
rect 2533 3704 2534 3877
rect 2317 3704 2318 3879
rect 2360 3878 2361 4295
rect 2318 3880 2319 4295
rect 2389 3704 2390 3881
rect 2348 3882 2349 4295
rect 2569 3704 2570 3883
rect 2354 3884 2355 4295
rect 2575 3704 2576 3885
rect 2390 3886 2391 4295
rect 2605 3704 2606 3887
rect 2323 3704 2324 3889
rect 2606 3888 2607 4295
rect 2324 3890 2325 4295
rect 2473 3704 2474 3891
rect 1999 3704 2000 3893
rect 2474 3892 2475 4295
rect 2000 3894 2001 4295
rect 2191 3704 2192 3895
rect 2192 3896 2193 4295
rect 2395 3704 2396 3897
rect 2396 3898 2397 4295
rect 2611 3704 2612 3899
rect 2422 3704 2423 3901
rect 2612 3900 2613 4295
rect 2438 3902 2439 4295
rect 2623 3704 2624 3903
rect 2444 3904 2445 4295
rect 2557 3704 2558 3905
rect 1993 3704 1994 3907
rect 2558 3906 2559 4295
rect 2446 3704 2447 3909
rect 2927 3908 2928 4295
rect 2456 3910 2457 4295
rect 3288 3910 3289 4295
rect 2462 3912 2463 4295
rect 3202 3704 3203 3913
rect 2479 3704 2480 3915
rect 2534 3914 2535 4295
rect 2119 3704 2120 3917
rect 2480 3916 2481 4295
rect 2120 3918 2121 4295
rect 2431 3704 2432 3919
rect 2432 3920 2433 4295
rect 2581 3704 2582 3921
rect 2485 3704 2486 3923
rect 3231 3922 3232 4295
rect 2125 3704 2126 3925
rect 2486 3924 2487 4295
rect 2126 3926 2127 4295
rect 2467 3704 2468 3927
rect 2468 3928 2469 4295
rect 2527 3704 2528 3929
rect 2504 3930 2505 4295
rect 2641 3704 2642 3931
rect 2509 3704 2510 3933
rect 3205 3704 3206 3933
rect 2510 3934 2511 4295
rect 3267 3934 3268 4295
rect 2528 3936 2529 4295
rect 3073 3704 3074 3937
rect 2540 3938 2541 4295
rect 2617 3704 2618 3939
rect 1849 3704 1850 3941
rect 2618 3940 2619 4295
rect 1621 3704 1622 3943
rect 1850 3942 1851 4295
rect 2563 3704 2564 3943
rect 3195 3704 3196 3943
rect 2383 3704 2384 3945
rect 2564 3944 2565 4295
rect 2155 3704 2156 3947
rect 2384 3946 2385 4295
rect 2156 3948 2157 4295
rect 2377 3704 2378 3949
rect 2005 3704 2006 3951
rect 2378 3950 2379 4295
rect 2006 3952 2007 4295
rect 2281 3704 2282 3953
rect 2282 3954 2283 4295
rect 2335 3704 2336 3955
rect 2336 3956 2337 4295
rect 2593 3704 2594 3957
rect 2570 3958 2571 4295
rect 2635 3704 2636 3959
rect 1753 3704 1754 3961
rect 2636 3960 2637 4295
rect 1478 3962 1479 4295
rect 1754 3962 1755 4295
rect 2576 3962 2577 4295
rect 2647 3704 2648 3963
rect 2582 3964 2583 4295
rect 2671 3704 2672 3965
rect 2594 3966 2595 4295
rect 3305 3966 3306 4295
rect 2624 3968 2625 4295
rect 2701 3704 2702 3969
rect 2642 3970 2643 4295
rect 2713 3704 2714 3971
rect 2659 3704 2660 3973
rect 2897 3972 2898 4295
rect 2660 3974 2661 4295
rect 3170 3704 3171 3975
rect 2666 3976 2667 4295
rect 3118 3704 3119 3977
rect 2672 3978 2673 4295
rect 2731 3704 2732 3979
rect 2683 3704 2684 3981
rect 3302 3980 3303 4295
rect 2684 3982 2685 4295
rect 2749 3704 2750 3983
rect 2689 3704 2690 3985
rect 3212 3704 3213 3985
rect 2690 3986 2691 4295
rect 2755 3704 2756 3987
rect 2695 3704 2696 3989
rect 3115 3704 3116 3989
rect 2696 3990 2697 4295
rect 2761 3704 2762 3991
rect 2702 3992 2703 4295
rect 2767 3704 2768 3993
rect 2714 3994 2715 4295
rect 3188 3704 3189 3995
rect 2725 3704 2726 3997
rect 3173 3704 3174 3997
rect 1861 3704 1862 3999
rect 2726 3998 2727 4295
rect 1862 4000 1863 4295
rect 2017 3704 2018 4001
rect 2018 4002 2019 4295
rect 2329 3704 2330 4003
rect 1987 3704 1988 4005
rect 2330 4004 2331 4295
rect 1988 4006 1989 4295
rect 2233 3704 2234 4007
rect 2234 4008 2235 4295
rect 3234 4008 3235 4295
rect 2732 4010 2733 4295
rect 2803 3704 2804 4011
rect 2743 3704 2744 4013
rect 3284 4012 3285 4295
rect 2744 4014 2745 4295
rect 2791 3704 2792 4015
rect 2750 4016 2751 4295
rect 2797 3704 2798 4017
rect 2756 4018 2757 4295
rect 2809 3704 2810 4019
rect 2762 4020 2763 4295
rect 2815 3704 2816 4021
rect 1807 3704 1808 4023
rect 2816 4022 2817 4295
rect 1808 4024 1809 4295
rect 1867 3704 1868 4025
rect 1868 4026 1869 4295
rect 2023 3704 2024 4027
rect 2024 4028 2025 4295
rect 2299 3704 2300 4029
rect 2300 4030 2301 4295
rect 2551 3704 2552 4031
rect 2065 3704 2066 4033
rect 2552 4032 2553 4295
rect 1475 4034 1476 4295
rect 2066 4034 2067 4295
rect 2768 4034 2769 4295
rect 2821 3704 2822 4035
rect 1795 3704 1796 4037
rect 2822 4036 2823 4295
rect 1796 4038 1797 4295
rect 1903 3704 1904 4039
rect 1500 4040 1501 4295
rect 1904 4040 1905 4295
rect 2779 3704 2780 4041
rect 3191 3704 3192 4041
rect 1825 3704 1826 4043
rect 2780 4042 2781 4295
rect 1826 4044 1827 4295
rect 1945 3704 1946 4045
rect 1946 4046 1947 4295
rect 2095 3704 2096 4047
rect 2096 4048 2097 4295
rect 2425 3704 2426 4049
rect 2426 4050 2427 4295
rect 2599 3704 2600 4051
rect 2600 4052 2601 4295
rect 2677 3704 2678 4053
rect 2678 4054 2679 4295
rect 3281 4054 3282 4295
rect 2792 4056 2793 4295
rect 2845 3704 2846 4057
rect 1709 4058 1710 4295
rect 2846 4058 2847 4295
rect 2798 4060 2799 4295
rect 3249 4060 3250 4295
rect 2804 4062 2805 4295
rect 2857 3704 2858 4063
rect 2080 3704 2081 4065
rect 2858 4064 2859 4295
rect 2081 4066 2082 4295
rect 2374 3704 2375 4067
rect 2810 4066 2811 4295
rect 2863 3704 2864 4067
rect 1747 3704 1748 4069
rect 2864 4068 2865 4295
rect 1748 4070 1749 4295
rect 1837 3704 1838 4071
rect 1838 4072 1839 4295
rect 1957 3704 1958 4073
rect 1958 4074 1959 4295
rect 2203 3704 2204 4075
rect 2204 4076 2205 4295
rect 2413 3704 2414 4077
rect 2113 3704 2114 4079
rect 2414 4078 2415 4295
rect 2114 4080 2115 4295
rect 2419 3704 2420 4081
rect 2420 4082 2421 4295
rect 2587 3704 2588 4083
rect 2588 4084 2589 4295
rect 2653 3704 2654 4085
rect 2654 4086 2655 4295
rect 2719 3704 2720 4087
rect 2720 4088 2721 4295
rect 2785 3704 2786 4089
rect 1921 3704 1922 4091
rect 2786 4090 2787 4295
rect 1922 4092 1923 4295
rect 2071 3704 2072 4093
rect 2053 3704 2054 4095
rect 2072 4094 2073 4295
rect 2054 4096 2055 4295
rect 2371 3704 2372 4097
rect 2221 3704 2222 4099
rect 2372 4098 2373 4295
rect 2222 4100 2223 4295
rect 3298 4100 3299 4295
rect 2839 3704 2840 4103
rect 3274 4102 3275 4295
rect 1741 3704 1742 4105
rect 2840 4104 2841 4295
rect 1742 4106 1743 4295
rect 1777 3704 1778 4107
rect 1723 3704 1724 4109
rect 1778 4108 1779 4295
rect 1724 4110 1725 4295
rect 1801 3704 1802 4111
rect 1802 4112 1803 4295
rect 1897 3704 1898 4113
rect 1891 3704 1892 4115
rect 1898 4114 1899 4295
rect 1892 4116 1893 4295
rect 2011 3704 2012 4117
rect 2012 4118 2013 4295
rect 2275 3704 2276 4119
rect 2276 4120 2277 4295
rect 2311 3704 2312 4121
rect 2245 3704 2246 4123
rect 2312 4122 2313 4295
rect 2246 4124 2247 4295
rect 2545 3704 2546 4125
rect 2029 3704 2030 4127
rect 2546 4126 2547 4295
rect 2852 4126 2853 4295
rect 2881 3704 2882 4127
rect 2855 4128 2856 4295
rect 3133 3704 3134 4129
rect 2869 3704 2870 4131
rect 2882 4130 2883 4295
rect 2875 3704 2876 4133
rect 3155 3704 3156 4133
rect 2876 4134 2877 4295
rect 2905 3704 2906 4135
rect 2879 4136 2880 4295
rect 2908 3704 2909 4137
rect 2884 3704 2885 4139
rect 3277 4138 3278 4295
rect 2900 4140 2901 4295
rect 3270 4140 3271 4295
rect 2906 4142 2907 4295
rect 3215 4142 3216 4295
rect 2917 3704 2918 4145
rect 2990 4144 2991 4295
rect 2918 4146 2919 4295
rect 3052 3704 3053 4147
rect 2923 3704 2924 4149
rect 3076 3704 3077 4149
rect 1601 4150 1602 4295
rect 2924 4150 2925 4295
rect 2941 3704 2942 4151
rect 2969 4150 2970 4295
rect 1525 3704 1526 4153
rect 2942 4152 2943 4295
rect 1526 4154 1527 4295
rect 1657 3704 1658 4155
rect 1427 3704 1428 4157
rect 1658 4156 1659 4295
rect 1427 4158 1428 4295
rect 2843 4158 2844 4295
rect 2971 3704 2972 4159
rect 3026 4158 3027 4295
rect 2893 3704 2894 4161
rect 2972 4160 2973 4295
rect 1759 3704 1760 4163
rect 2894 4162 2895 4295
rect 1760 4164 1761 4295
rect 1831 3704 1832 4165
rect 1681 3704 1682 4167
rect 1832 4166 1833 4295
rect 1682 4168 1683 4295
rect 1711 3704 1712 4169
rect 1699 3704 1700 4171
rect 1712 4170 1713 4295
rect 1700 4172 1701 4295
rect 1729 3704 1730 4173
rect 1730 4174 1731 4295
rect 1819 3704 1820 4175
rect 1820 4176 1821 4295
rect 1933 3704 1934 4177
rect 1934 4178 1935 4295
rect 3158 4178 3159 4295
rect 3001 3704 3002 4181
rect 3068 4180 3069 4295
rect 2947 3704 2948 4183
rect 3002 4182 3003 4295
rect 2944 3704 2945 4185
rect 2948 4184 2949 4295
rect 2470 3704 2471 4187
rect 2945 4186 2946 4295
rect 3008 4186 3009 4295
rect 3219 3704 3220 4187
rect 3019 3704 3020 4189
rect 3104 4188 3105 4295
rect 3020 4190 3021 4295
rect 3295 4190 3296 4295
rect 3022 3704 3023 4193
rect 3107 4192 3108 4295
rect 3031 3704 3032 4195
rect 3101 4194 3102 4295
rect 2977 3704 2978 4197
rect 3032 4196 3033 4295
rect 2911 3704 2912 4199
rect 2978 4198 2979 4295
rect 2912 4200 2913 4295
rect 3136 3704 3137 4201
rect 3034 3704 3035 4203
rect 3086 4202 3087 4295
rect 3040 3704 3041 4205
rect 3113 4204 3114 4295
rect 3043 3704 3044 4207
rect 3134 4206 3135 4295
rect 3044 4208 3045 4295
rect 3142 3704 3143 4209
rect 2648 4210 2649 4295
rect 3143 4210 3144 4295
rect 3049 3704 3050 4213
rect 3145 3704 3146 4213
rect 2965 3704 2966 4215
rect 3050 4214 3051 4295
rect 2966 4216 2967 4295
rect 3209 3704 3210 4217
rect 3055 3704 3056 4219
rect 3146 4218 3147 4295
rect 3061 3704 3062 4221
rect 3203 4220 3204 4295
rect 2995 3704 2996 4223
rect 3062 4222 3063 4295
rect 2887 3704 2888 4225
rect 2996 4224 2997 4295
rect 1915 3704 1916 4227
rect 2888 4226 2889 4295
rect 1431 3704 1432 4229
rect 1916 4228 1917 4295
rect 1431 4230 1432 4295
rect 1586 4230 1587 4295
rect 3091 3704 3092 4231
rect 3176 4230 3177 4295
rect 3109 3704 3110 4233
rect 3197 4232 3198 4295
rect 3037 3704 3038 4235
rect 3110 4234 3111 4295
rect 2983 3704 2984 4237
rect 3038 4236 3039 4295
rect 2935 3704 2936 4239
rect 2984 4238 2985 4295
rect 2936 4240 2937 4295
rect 3148 3704 3149 4241
rect 3121 3704 3122 4243
rect 3200 4242 3201 4295
rect 3122 4244 3123 4295
rect 3224 4244 3225 4295
rect 3124 3704 3125 4247
rect 3161 4246 3162 4295
rect 3127 3704 3128 4249
rect 3206 4248 3207 4295
rect 1420 3704 1421 4251
rect 3128 4250 3129 4295
rect 1420 4252 1421 4295
rect 1994 4252 1995 4295
rect 3130 3704 3131 4253
rect 3209 4252 3210 4295
rect 3139 3704 3140 4255
rect 3218 4254 3219 4295
rect 2305 3704 2306 4257
rect 3140 4256 3141 4295
rect 1963 3704 1964 4259
rect 2306 4258 2307 4295
rect 1964 4260 1965 4295
rect 2035 3704 2036 4261
rect 1471 3704 1472 4263
rect 2036 4262 2037 4295
rect 1471 4264 1472 4295
rect 2030 4264 2031 4295
rect 3152 3704 3153 4265
rect 3194 4264 3195 4295
rect 3164 3704 3165 4267
rect 3243 4266 3244 4295
rect 3079 3704 3080 4269
rect 3164 4268 3165 4295
rect 3013 3704 3014 4271
rect 3080 4270 3081 4295
rect 2953 3704 2954 4273
rect 3014 4272 3015 4295
rect 2833 3704 2834 4275
rect 2954 4274 2955 4295
rect 1789 3704 1790 4277
rect 2834 4276 2835 4295
rect 1790 4278 1791 4295
rect 1885 3704 1886 4279
rect 1886 4280 1887 4295
rect 1951 3704 1952 4281
rect 1441 3704 1442 4283
rect 1952 4282 1953 4295
rect 1441 4284 1442 4295
rect 2048 4284 2049 4295
rect 3167 3704 3168 4285
rect 3246 4284 3247 4295
rect 3182 3704 3183 4287
rect 3261 4286 3262 4295
rect 3097 3704 3098 4289
rect 3182 4288 3183 4295
rect 3098 4290 3099 4295
rect 3212 4290 3213 4295
rect 3185 3704 3186 4293
rect 3264 4292 3265 4295
rect 1431 4299 1432 4302
rect 1580 4299 1581 4302
rect 1441 4299 1442 4304
rect 1550 4303 1551 4918
rect 1441 4305 1442 4918
rect 2024 4299 2025 4306
rect 1450 4305 1451 4918
rect 1450 4299 1451 4306
rect 1456 4305 1457 4918
rect 1456 4299 1457 4306
rect 1462 4305 1463 4918
rect 1462 4299 1463 4306
rect 1468 4299 1469 4308
rect 2042 4299 2043 4308
rect 1468 4309 1469 4918
rect 2006 4299 2007 4310
rect 1494 4309 1495 4918
rect 1494 4299 1495 4310
rect 1503 4299 1504 4312
rect 1910 4299 1911 4312
rect 1510 4299 1511 4314
rect 1622 4313 1623 4918
rect 1510 4315 1511 4918
rect 1922 4299 1923 4316
rect 1517 4299 1518 4318
rect 3311 4317 3312 4918
rect 1517 4319 1518 4918
rect 1940 4299 1941 4320
rect 1526 4299 1527 4322
rect 1652 4299 1653 4322
rect 1485 4299 1486 4324
rect 1526 4323 1527 4918
rect 1485 4325 1486 4918
rect 2000 4299 2001 4326
rect 1541 4327 1542 4918
rect 2828 4299 2829 4328
rect 1586 4299 1587 4330
rect 1616 4329 1617 4918
rect 1601 4299 1602 4332
rect 3243 4299 3244 4332
rect 1610 4299 1611 4334
rect 1634 4333 1635 4918
rect 1434 4299 1435 4336
rect 1610 4335 1611 4918
rect 1628 4299 1629 4336
rect 1652 4335 1653 4918
rect 1507 4299 1508 4338
rect 1628 4337 1629 4918
rect 1507 4339 1508 4918
rect 1838 4299 1839 4340
rect 1500 4299 1501 4342
rect 1838 4341 1839 4918
rect 1500 4343 1501 4918
rect 1778 4299 1779 4344
rect 1640 4299 1641 4346
rect 1676 4345 1677 4918
rect 1604 4299 1605 4348
rect 1640 4347 1641 4918
rect 1661 4347 1662 4918
rect 3032 4299 3033 4348
rect 1709 4299 1710 4350
rect 2858 4299 2859 4350
rect 1514 4299 1515 4352
rect 2858 4351 2859 4918
rect 1478 4299 1479 4354
rect 1514 4353 1515 4918
rect 1778 4353 1779 4918
rect 2864 4299 2865 4354
rect 1856 4299 1857 4356
rect 2000 4355 2001 4918
rect 1434 4357 1435 4918
rect 1856 4357 1857 4918
rect 1868 4299 1869 4358
rect 2042 4357 2043 4918
rect 1754 4299 1755 4360
rect 1868 4359 1869 4918
rect 1424 4299 1425 4362
rect 1754 4361 1755 4918
rect 1424 4363 1425 4918
rect 1742 4299 1743 4364
rect 1712 4299 1713 4366
rect 1742 4365 1743 4918
rect 1712 4367 1713 4918
rect 1832 4299 1833 4368
rect 1832 4369 1833 4918
rect 2846 4299 2847 4370
rect 1871 4299 1872 4372
rect 2045 4371 2046 4918
rect 1880 4299 1881 4374
rect 2024 4373 2025 4918
rect 1772 4299 1773 4376
rect 1880 4375 1881 4918
rect 1682 4299 1683 4378
rect 1772 4377 1773 4918
rect 1886 4299 1887 4378
rect 2006 4377 2007 4918
rect 1886 4379 1887 4918
rect 2834 4299 2835 4380
rect 1898 4299 1899 4382
rect 1922 4381 1923 4918
rect 1898 4383 1899 4918
rect 2822 4299 2823 4384
rect 1940 4385 1941 4918
rect 3300 4385 3301 4918
rect 1961 4299 1962 4388
rect 2147 4387 2148 4918
rect 2003 4299 2004 4390
rect 2159 4389 2160 4918
rect 2027 4299 2028 4392
rect 2231 4391 2232 4918
rect 2051 4299 2052 4394
rect 2273 4393 2274 4918
rect 2063 4299 2064 4396
rect 2291 4395 2292 4918
rect 2081 4299 2082 4398
rect 2279 4397 2280 4918
rect 2099 4299 2100 4400
rect 2321 4399 2322 4918
rect 2105 4299 2106 4402
rect 2327 4401 2328 4918
rect 2216 4299 2217 4404
rect 3234 4299 3235 4404
rect 2216 4405 2217 4918
rect 2474 4299 2475 4406
rect 2246 4299 2247 4408
rect 2474 4407 2475 4918
rect 2288 4299 2289 4410
rect 3143 4299 3144 4410
rect 2060 4299 2061 4412
rect 2288 4411 2289 4918
rect 1892 4299 1893 4414
rect 2060 4413 2061 4918
rect 1748 4299 1749 4416
rect 1892 4415 1893 4918
rect 1748 4417 1749 4918
rect 1784 4299 1785 4418
rect 1784 4419 1785 4918
rect 2612 4299 2613 4420
rect 2357 4421 2358 4918
rect 2897 4299 2898 4422
rect 2402 4299 2403 4424
rect 3370 4423 3371 4918
rect 2192 4299 2193 4426
rect 2402 4425 2403 4918
rect 2108 4299 2109 4428
rect 2192 4427 2193 4918
rect 2429 4427 2430 4918
rect 2843 4299 2844 4428
rect 2438 4299 2439 4430
rect 2612 4429 2613 4918
rect 2438 4431 2439 4918
rect 2546 4299 2547 4432
rect 2354 4299 2355 4434
rect 2546 4433 2547 4918
rect 2186 4299 2187 4436
rect 2354 4435 2355 4918
rect 2186 4437 2187 4918
rect 2558 4299 2559 4438
rect 2384 4299 2385 4440
rect 2558 4439 2559 4918
rect 2162 4299 2163 4442
rect 2384 4441 2385 4918
rect 2162 4443 2163 4918
rect 2252 4299 2253 4444
rect 2252 4445 2253 4918
rect 2270 4299 2271 4446
rect 2048 4299 2049 4448
rect 2270 4447 2271 4918
rect 2048 4449 2049 4918
rect 2306 4299 2307 4450
rect 2138 4299 2139 4452
rect 2306 4451 2307 4918
rect 1976 4299 1977 4454
rect 2138 4453 2139 4918
rect 1478 4455 1479 4918
rect 1976 4455 1977 4918
rect 2450 4299 2451 4456
rect 3395 4455 3396 4918
rect 2222 4299 2223 4458
rect 2450 4457 2451 4918
rect 2018 4299 2019 4460
rect 2222 4459 2223 4918
rect 1874 4299 1875 4462
rect 2018 4461 2019 4918
rect 1760 4299 1761 4464
rect 1874 4463 1875 4918
rect 1503 4465 1504 4918
rect 1760 4465 1761 4918
rect 2504 4299 2505 4466
rect 3367 4465 3368 4918
rect 2294 4299 2295 4468
rect 2504 4467 2505 4918
rect 1427 4299 1428 4470
rect 2294 4469 2295 4918
rect 1427 4471 1428 4918
rect 2108 4471 2109 4918
rect 2594 4299 2595 4472
rect 2738 4471 2739 4918
rect 2426 4299 2427 4474
rect 2594 4473 2595 4918
rect 2210 4299 2211 4476
rect 2426 4475 2427 4918
rect 2078 4299 2079 4478
rect 2210 4477 2211 4918
rect 1904 4299 1905 4480
rect 2078 4479 2079 4918
rect 1808 4299 1809 4482
rect 1904 4481 1905 4918
rect 1420 4299 1421 4484
rect 1808 4483 1809 4918
rect 1420 4485 1421 4918
rect 2246 4485 2247 4918
rect 2684 4299 2685 4486
rect 3281 4299 3282 4486
rect 2534 4299 2535 4488
rect 2684 4487 2685 4918
rect 2414 4299 2415 4490
rect 2534 4489 2535 4918
rect 2414 4491 2415 4918
rect 3326 4491 3327 4918
rect 2690 4299 2691 4494
rect 2828 4493 2829 4918
rect 2540 4299 2541 4496
rect 2690 4495 2691 4918
rect 2348 4299 2349 4498
rect 2540 4497 2541 4918
rect 2126 4299 2127 4500
rect 2348 4499 2349 4918
rect 1970 4299 1971 4502
rect 2126 4501 2127 4918
rect 1820 4299 1821 4504
rect 1970 4503 1971 4918
rect 1820 4505 1821 4918
rect 2924 4299 2925 4506
rect 2696 4299 2697 4508
rect 2834 4507 2835 4918
rect 2696 4509 2697 4918
rect 2726 4299 2727 4510
rect 2582 4299 2583 4512
rect 2726 4511 2727 4918
rect 2390 4299 2391 4514
rect 2582 4513 2583 4918
rect 1417 4299 1418 4516
rect 2390 4515 2391 4918
rect 1417 4517 1418 4918
rect 1482 4299 1483 4518
rect 1482 4519 1483 4918
rect 1994 4299 1995 4520
rect 1850 4299 1851 4522
rect 1994 4521 1995 4918
rect 1475 4299 1476 4524
rect 1850 4523 1851 4918
rect 2708 4299 2709 4524
rect 3023 4523 3024 4918
rect 2570 4299 2571 4526
rect 2708 4525 2709 4918
rect 2408 4299 2409 4528
rect 2570 4527 2571 4918
rect 2198 4299 2199 4530
rect 2408 4529 2409 4918
rect 2030 4299 2031 4532
rect 2198 4531 2199 4918
rect 2030 4533 2031 4918
rect 2456 4299 2457 4534
rect 2456 4535 2457 4918
rect 3398 4535 3399 4918
rect 2714 4299 2715 4538
rect 3333 4537 3334 4918
rect 2576 4299 2577 4540
rect 2714 4539 2715 4918
rect 2480 4299 2481 4542
rect 2576 4541 2577 4918
rect 2282 4299 2283 4544
rect 2480 4543 2481 4918
rect 1438 4299 1439 4546
rect 2282 4545 2283 4918
rect 2786 4299 2787 4546
rect 2924 4545 2925 4918
rect 2648 4299 2649 4548
rect 2786 4547 2787 4918
rect 2516 4299 2517 4550
rect 2648 4549 2649 4918
rect 2324 4299 2325 4552
rect 2516 4551 2517 4918
rect 2102 4299 2103 4554
rect 2324 4553 2325 4918
rect 1964 4299 1965 4556
rect 2102 4555 2103 4918
rect 1538 4557 1539 4918
rect 1964 4557 1965 4918
rect 2792 4299 2793 4558
rect 2930 4557 2931 4918
rect 2654 4299 2655 4560
rect 2792 4559 2793 4918
rect 2492 4299 2493 4562
rect 2654 4561 2655 4918
rect 2342 4299 2343 4564
rect 2492 4563 2493 4918
rect 2120 4299 2121 4566
rect 2342 4565 2343 4918
rect 1946 4299 1947 4568
rect 2120 4567 2121 4918
rect 1946 4569 1947 4918
rect 3252 4299 3253 4570
rect 2822 4571 2823 4918
rect 3284 4299 3285 4572
rect 2840 4299 2841 4574
rect 3374 4573 3375 4918
rect 2702 4299 2703 4576
rect 2840 4575 2841 4918
rect 2564 4299 2565 4578
rect 2702 4577 2703 4918
rect 2522 4299 2523 4580
rect 2564 4579 2565 4918
rect 2372 4299 2373 4582
rect 2522 4581 2523 4918
rect 2180 4299 2181 4584
rect 2372 4583 2373 4918
rect 2180 4585 2181 4918
rect 2264 4299 2265 4586
rect 2084 4299 2085 4588
rect 2264 4587 2265 4918
rect 1928 4299 1929 4590
rect 2084 4589 2085 4918
rect 1814 4299 1815 4592
rect 1928 4591 1929 4918
rect 1814 4593 1815 4918
rect 2636 4299 2637 4594
rect 2486 4299 2487 4596
rect 2636 4595 2637 4918
rect 2360 4299 2361 4598
rect 2486 4597 2487 4918
rect 2150 4299 2151 4600
rect 2360 4599 2361 4918
rect 2150 4601 2151 4918
rect 2228 4299 2229 4602
rect 1438 4603 1439 4918
rect 2228 4603 2229 4918
rect 2855 4299 2856 4604
rect 2870 4603 2871 4918
rect 2864 4605 2865 4918
rect 3323 4605 3324 4918
rect 2876 4299 2877 4608
rect 3270 4299 3271 4608
rect 2744 4299 2745 4610
rect 2876 4609 2877 4918
rect 2600 4299 2601 4612
rect 2744 4611 2745 4918
rect 2420 4299 2421 4614
rect 2600 4613 2601 4918
rect 2204 4299 2205 4616
rect 2420 4615 2421 4918
rect 1471 4299 1472 4618
rect 2204 4617 2205 4918
rect 1471 4619 1472 4918
rect 2012 4299 2013 4620
rect 1844 4299 1845 4622
rect 2012 4621 2013 4918
rect 1724 4299 1725 4624
rect 1844 4623 1845 4918
rect 1664 4299 1665 4626
rect 1724 4625 1725 4918
rect 1529 4299 1530 4628
rect 1664 4627 1665 4918
rect 1529 4629 1530 4918
rect 1604 4629 1605 4918
rect 2906 4299 2907 4630
rect 3158 4299 3159 4630
rect 2906 4631 2907 4918
rect 3291 4299 3292 4632
rect 2918 4299 2919 4634
rect 3215 4299 3216 4634
rect 2816 4299 2817 4636
rect 2918 4635 2919 4918
rect 2678 4299 2679 4638
rect 2816 4637 2817 4918
rect 2552 4299 2553 4640
rect 2678 4639 2679 4918
rect 2336 4299 2337 4642
rect 2552 4641 2553 4918
rect 2114 4299 2115 4644
rect 2336 4643 2337 4918
rect 1952 4299 1953 4646
rect 2114 4645 2115 4918
rect 1796 4299 1797 4648
rect 1952 4647 1953 4918
rect 1796 4649 1797 4918
rect 2894 4299 2895 4650
rect 2762 4299 2763 4652
rect 2894 4651 2895 4918
rect 2624 4299 2625 4654
rect 2762 4653 2763 4918
rect 2462 4299 2463 4656
rect 2624 4655 2625 4918
rect 2240 4299 2241 4658
rect 2462 4657 2463 4918
rect 2036 4299 2037 4660
rect 2240 4659 2241 4918
rect 1862 4299 1863 4662
rect 2036 4661 2037 4918
rect 1730 4299 1731 4664
rect 1862 4663 1863 4918
rect 1670 4299 1671 4666
rect 1730 4665 1731 4918
rect 2921 4665 2922 4918
rect 2927 4299 2928 4666
rect 2945 4299 2946 4666
rect 2999 4665 3000 4918
rect 2966 4299 2967 4668
rect 3092 4667 3093 4918
rect 2966 4669 2967 4918
rect 3237 4669 3238 4918
rect 2969 4299 2970 4672
rect 3095 4671 3096 4918
rect 3002 4299 3003 4674
rect 3116 4673 3117 4918
rect 2852 4299 2853 4676
rect 3002 4675 3003 4918
rect 2720 4299 2721 4678
rect 2852 4677 2853 4918
rect 2588 4299 2589 4680
rect 2720 4679 2721 4918
rect 2396 4299 2397 4682
rect 2588 4681 2589 4918
rect 2174 4299 2175 4684
rect 2396 4683 2397 4918
rect 1988 4299 1989 4686
rect 2174 4685 2175 4918
rect 1431 4687 1432 4918
rect 1988 4687 1989 4918
rect 3005 4687 3006 4918
rect 3288 4299 3289 4688
rect 3014 4299 3015 4690
rect 3032 4689 3033 4918
rect 3014 4691 3015 4918
rect 3212 4299 3213 4692
rect 3038 4299 3039 4694
rect 3295 4299 3296 4694
rect 2972 4299 2973 4696
rect 3038 4695 3039 4918
rect 1706 4299 1707 4698
rect 2972 4697 2973 4918
rect 1706 4699 1707 4918
rect 1718 4299 1719 4700
rect 1658 4299 1659 4702
rect 1718 4701 1719 4918
rect 1658 4703 1659 4918
rect 3305 4299 3306 4704
rect 2996 4299 2997 4706
rect 3304 4705 3305 4918
rect 2942 4299 2943 4708
rect 2996 4707 2997 4918
rect 2942 4709 2943 4918
rect 3274 4299 3275 4710
rect 3056 4711 3057 4918
rect 3377 4711 3378 4918
rect 3062 4299 3063 4714
rect 3158 4713 3159 4918
rect 2936 4299 2937 4716
rect 3062 4715 3063 4918
rect 2798 4299 2799 4718
rect 2936 4717 2937 4918
rect 2660 4299 2661 4720
rect 2798 4719 2799 4918
rect 2498 4299 2499 4722
rect 2660 4721 2661 4918
rect 2318 4299 2319 4724
rect 2498 4723 2499 4918
rect 2090 4299 2091 4726
rect 2318 4725 2319 4918
rect 2090 4727 2091 4918
rect 3298 4299 3299 4728
rect 3068 4299 3069 4730
rect 3152 4729 3153 4918
rect 2948 4299 2949 4732
rect 3068 4731 3069 4918
rect 2804 4299 2805 4734
rect 2948 4733 2949 4918
rect 2672 4299 2673 4736
rect 2804 4735 2805 4918
rect 2528 4299 2529 4738
rect 2672 4737 2673 4918
rect 2366 4299 2367 4740
rect 2528 4739 2529 4918
rect 2144 4299 2145 4742
rect 2366 4741 2367 4918
rect 1958 4299 1959 4744
rect 2144 4743 2145 4918
rect 1802 4299 1803 4746
rect 1958 4745 1959 4918
rect 1802 4747 1803 4918
rect 2900 4299 2901 4748
rect 2768 4299 2769 4750
rect 2900 4749 2901 4918
rect 2630 4299 2631 4752
rect 2768 4751 2769 4918
rect 2468 4299 2469 4754
rect 2630 4753 2631 4918
rect 2234 4299 2235 4756
rect 2468 4755 2469 4918
rect 2234 4757 2235 4918
rect 2312 4299 2313 4758
rect 2096 4299 2097 4760
rect 2312 4759 2313 4918
rect 1934 4299 1935 4762
rect 2096 4761 2097 4918
rect 1790 4299 1791 4764
rect 1934 4763 1935 4918
rect 1700 4299 1701 4766
rect 1790 4765 1791 4918
rect 1598 4299 1599 4768
rect 1700 4767 1701 4918
rect 1568 4299 1569 4770
rect 1598 4769 1599 4918
rect 3074 4769 3075 4918
rect 3277 4299 3278 4770
rect 3080 4299 3081 4772
rect 3249 4299 3250 4772
rect 2990 4299 2991 4774
rect 3080 4773 3081 4918
rect 2990 4775 2991 4918
rect 3384 4775 3385 4918
rect 3098 4299 3099 4778
rect 3188 4777 3189 4918
rect 2978 4299 2979 4780
rect 3098 4779 3099 4918
rect 2888 4299 2889 4782
rect 2978 4781 2979 4918
rect 2756 4299 2757 4784
rect 2888 4783 2889 4918
rect 2666 4299 2667 4786
rect 2756 4785 2757 4918
rect 2510 4299 2511 4788
rect 2666 4787 2667 4918
rect 2300 4299 2301 4790
rect 2510 4789 2511 4918
rect 2132 4299 2133 4792
rect 2300 4791 2301 4918
rect 2072 4299 2073 4794
rect 2132 4793 2133 4918
rect 1916 4299 1917 4796
rect 2072 4795 2073 4918
rect 1916 4797 1917 4918
rect 2618 4299 2619 4798
rect 2444 4299 2445 4800
rect 2618 4799 2619 4918
rect 2258 4299 2259 4802
rect 2444 4801 2445 4918
rect 2066 4299 2067 4804
rect 2258 4803 2259 4918
rect 2066 4805 2067 4918
rect 2378 4299 2379 4806
rect 2168 4299 2169 4808
rect 2378 4807 2379 4918
rect 1982 4299 1983 4810
rect 2168 4809 2169 4918
rect 1826 4299 1827 4812
rect 1982 4811 1983 4918
rect 1736 4299 1737 4814
rect 1826 4813 1827 4918
rect 1688 4299 1689 4816
rect 1736 4815 1737 4918
rect 1688 4817 1689 4918
rect 1694 4299 1695 4818
rect 3101 4299 3102 4818
rect 3191 4817 3192 4918
rect 3104 4299 3105 4820
rect 3215 4819 3216 4918
rect 2984 4299 2985 4822
rect 3104 4821 3105 4918
rect 3128 4299 3129 4822
rect 3224 4299 3225 4822
rect 3050 4299 3051 4824
rect 3128 4823 3129 4918
rect 2912 4299 2913 4826
rect 3050 4825 3051 4918
rect 2774 4299 2775 4828
rect 2912 4827 2913 4918
rect 2774 4829 2775 4918
rect 3302 4299 3303 4830
rect 3134 4299 3135 4832
rect 3227 4299 3228 4832
rect 3026 4299 3027 4834
rect 3134 4833 3135 4918
rect 2882 4299 2883 4836
rect 3026 4835 3027 4918
rect 2750 4299 2751 4838
rect 2882 4837 2883 4918
rect 2750 4839 2751 4918
rect 2780 4299 2781 4840
rect 2642 4299 2643 4842
rect 2780 4841 2781 4918
rect 2642 4843 2643 4918
rect 3360 4843 3361 4918
rect 3140 4299 3141 4846
rect 3161 4299 3162 4846
rect 3164 4299 3165 4846
rect 3243 4845 3244 4918
rect 3107 4299 3108 4848
rect 3164 4847 3165 4918
rect 3176 4299 3177 4848
rect 3320 4847 3321 4918
rect 3086 4299 3087 4850
rect 3176 4849 3177 4918
rect 3194 4299 3195 4850
rect 3273 4849 3274 4918
rect 3110 4299 3111 4852
rect 3194 4851 3195 4918
rect 3008 4299 3009 4854
rect 3110 4853 3111 4918
rect 2954 4299 2955 4856
rect 3008 4855 3009 4918
rect 2810 4299 2811 4858
rect 2954 4857 2955 4918
rect 2732 4299 2733 4860
rect 2810 4859 2811 4918
rect 2606 4299 2607 4862
rect 2732 4861 2733 4918
rect 2432 4299 2433 4864
rect 2606 4863 2607 4918
rect 2276 4299 2277 4866
rect 2432 4865 2433 4918
rect 2054 4299 2055 4868
rect 2276 4867 2277 4918
rect 2054 4869 2055 4918
rect 2330 4299 2331 4870
rect 2156 4299 2157 4872
rect 2330 4871 2331 4918
rect 2156 4873 2157 4918
rect 3231 4299 3232 4874
rect 3170 4875 3171 4918
rect 3230 4875 3231 4918
rect 3197 4299 3198 4878
rect 3276 4877 3277 4918
rect 3113 4299 3114 4880
rect 3197 4879 3198 4918
rect 3200 4299 3201 4880
rect 3294 4879 3295 4918
rect 3200 4881 3201 4918
rect 3221 4299 3222 4882
rect 3203 4299 3204 4884
rect 3224 4883 3225 4918
rect 3044 4299 3045 4886
rect 3203 4885 3204 4918
rect 1475 4887 1476 4918
rect 3044 4887 3045 4918
rect 3206 4299 3207 4888
rect 3285 4887 3286 4918
rect 3122 4299 3123 4890
rect 3206 4889 3207 4918
rect 3020 4299 3021 4892
rect 3122 4891 3123 4918
rect 2879 4299 2880 4894
rect 3020 4893 3021 4918
rect 3209 4299 3210 4894
rect 3288 4893 3289 4918
rect 3212 4895 3213 4918
rect 3307 4895 3308 4918
rect 3218 4299 3219 4898
rect 3233 4897 3234 4918
rect 3146 4299 3147 4900
rect 3218 4899 3219 4918
rect 3240 4899 3241 4918
rect 3314 4899 3315 4918
rect 3246 4299 3247 4902
rect 3317 4901 3318 4918
rect 3261 4299 3262 4904
rect 3354 4903 3355 4918
rect 3182 4299 3183 4906
rect 3261 4905 3262 4918
rect 3264 4299 3265 4906
rect 3357 4905 3358 4918
rect 3267 4299 3268 4908
rect 3297 4907 3298 4918
rect 3291 4909 3292 4918
rect 3363 4909 3364 4918
rect 3330 4911 3331 4918
rect 3381 4911 3382 4918
rect 3336 4913 3337 4918
rect 3388 4913 3389 4918
rect 3342 4915 3343 4918
rect 3391 4915 3392 4918
rect 1434 4922 1435 4925
rect 1952 4922 1953 4925
rect 1438 4922 1439 4927
rect 2138 4922 2139 4927
rect 1447 4928 1448 5573
rect 2060 4922 2061 4929
rect 1471 4922 1472 4931
rect 2006 4922 2007 4931
rect 1478 4922 1479 4933
rect 1970 4922 1971 4933
rect 1477 4934 1478 5573
rect 1988 4922 1989 4935
rect 1482 4922 1483 4937
rect 2156 4922 2157 4937
rect 1488 4938 1489 5573
rect 2327 4922 2328 4939
rect 1491 4940 1492 5573
rect 2282 4922 2283 4941
rect 1503 4922 1504 4943
rect 1748 4922 1749 4943
rect 1514 4922 1515 4945
rect 2312 4922 2313 4945
rect 1510 4922 1511 4947
rect 2312 4946 2313 5573
rect 1517 4922 1518 4949
rect 2879 4948 2880 5573
rect 1519 4950 1520 5573
rect 2192 4922 2193 4951
rect 1526 4922 1527 4953
rect 1904 4922 1905 4953
rect 1526 4954 1527 5573
rect 2504 4922 2505 4955
rect 1529 4922 1530 4957
rect 3014 4922 3015 4957
rect 1538 4922 1539 4959
rect 1886 4922 1887 4959
rect 1541 4922 1542 4961
rect 1838 4922 1839 4961
rect 1468 4922 1469 4963
rect 1838 4962 1839 5573
rect 1462 4922 1463 4965
rect 1468 4964 1469 5573
rect 1456 4922 1457 4967
rect 1462 4966 1463 5573
rect 1450 4922 1451 4969
rect 1456 4968 1457 5573
rect 1544 4968 1545 5573
rect 1544 4922 1545 4969
rect 1556 4922 1557 4969
rect 2825 4968 2826 5573
rect 1574 4922 1575 4971
rect 1586 4970 1587 5573
rect 1580 4972 1581 5573
rect 2147 4922 2148 4973
rect 1634 4922 1635 4975
rect 1646 4974 1647 5573
rect 1622 4922 1623 4977
rect 1634 4976 1635 5573
rect 1610 4922 1611 4979
rect 1622 4978 1623 5573
rect 1598 4922 1599 4981
rect 1610 4980 1611 5573
rect 1562 4922 1563 4983
rect 1598 4982 1599 5573
rect 1550 4922 1551 4985
rect 1562 4984 1563 5573
rect 1652 4922 1653 4985
rect 1670 4984 1671 5573
rect 1640 4922 1641 4987
rect 1652 4986 1653 5573
rect 1628 4922 1629 4989
rect 1640 4988 1641 5573
rect 1616 4922 1617 4991
rect 1628 4990 1629 5573
rect 1694 4990 1695 5573
rect 1718 4922 1719 4991
rect 1742 4922 1743 4991
rect 1766 4990 1767 5573
rect 1742 4992 1743 5573
rect 1790 4922 1791 4993
rect 1748 4994 1749 5573
rect 1754 4922 1755 4995
rect 1688 4922 1689 4997
rect 1754 4996 1755 5573
rect 1481 4998 1482 5573
rect 1688 4998 1689 5573
rect 1790 4998 1791 5573
rect 1844 4922 1845 4999
rect 1829 5000 1830 5573
rect 2045 4922 2046 5001
rect 1844 5002 1845 5573
rect 2072 4922 2073 5003
rect 1904 5004 1905 5573
rect 2288 4922 2289 5005
rect 1661 4922 1662 5007
rect 2288 5006 2289 5573
rect 1907 5008 1908 5573
rect 2291 4922 2292 5009
rect 1910 5010 1911 5573
rect 2228 4922 2229 5011
rect 1937 5012 1938 5573
rect 2231 4922 2232 5013
rect 1952 5014 1953 5573
rect 2240 4922 2241 5015
rect 1970 5016 1971 5573
rect 2348 4922 2349 5017
rect 1976 4922 1977 5019
rect 2192 5018 2193 5573
rect 1976 5020 1977 5573
rect 2342 4922 2343 5021
rect 1982 4922 1983 5023
rect 2156 5022 2157 5573
rect 1982 5024 1983 5573
rect 2204 4922 2205 5025
rect 1988 5026 1989 5573
rect 2366 4922 2367 5027
rect 2006 5028 2007 5573
rect 2360 4922 2361 5029
rect 2060 5030 2061 5573
rect 2264 4922 2265 5031
rect 2069 5032 2070 5573
rect 2273 4922 2274 5033
rect 2072 5034 2073 5573
rect 2300 4922 2301 5035
rect 2102 4922 2103 5037
rect 2348 5036 2349 5573
rect 2102 5038 2103 5573
rect 2402 4922 2403 5039
rect 2132 4922 2133 5041
rect 2360 5040 2361 5573
rect 2132 5042 2133 5573
rect 2408 4922 2409 5043
rect 2126 4922 2127 5045
rect 2408 5044 2409 5573
rect 2126 5046 2127 5573
rect 2462 4922 2463 5047
rect 2138 5048 2139 5573
rect 2420 4922 2421 5049
rect 2150 4922 2151 5051
rect 2228 5050 2229 5573
rect 2150 5052 2151 5573
rect 2426 4922 2427 5053
rect 2159 4922 2160 5055
rect 2573 5054 2574 5573
rect 2180 4922 2181 5057
rect 2300 5056 2301 5573
rect 2090 4922 2091 5059
rect 2180 5058 2181 5573
rect 2090 5060 2091 5573
rect 2450 4922 2451 5061
rect 2204 5062 2205 5573
rect 2510 4922 2511 5063
rect 2234 4922 2235 5065
rect 2240 5064 2241 5573
rect 2234 5066 2235 5573
rect 3326 4922 3327 5067
rect 2264 5068 2265 5573
rect 2540 4922 2541 5069
rect 2282 5070 2283 5573
rect 2294 4922 2295 5071
rect 2294 5072 2295 5573
rect 2492 4922 2493 5073
rect 1868 4922 1869 5075
rect 2492 5074 2493 5573
rect 2342 5076 2343 5573
rect 2594 4922 2595 5077
rect 1760 4922 1761 5079
rect 2594 5078 2595 5573
rect 1760 5080 1761 5573
rect 1862 4922 1863 5081
rect 1862 5082 1863 5573
rect 2144 4922 2145 5083
rect 2144 5084 2145 5573
rect 2474 4922 2475 5085
rect 1874 4922 1875 5087
rect 2474 5086 2475 5573
rect 1658 4922 1659 5089
rect 1874 5088 1875 5573
rect 1604 4922 1605 5091
rect 1658 5090 1659 5573
rect 1592 4922 1593 5093
rect 1604 5092 1605 5573
rect 1433 5094 1434 5573
rect 1592 5094 1593 5573
rect 2357 4922 2358 5095
rect 3035 5094 3036 5573
rect 2279 4922 2280 5097
rect 2357 5096 2358 5573
rect 2366 5096 2367 5573
rect 2600 4922 2601 5097
rect 2216 4922 2217 5099
rect 2600 5098 2601 5573
rect 2216 5100 2217 5573
rect 2480 4922 2481 5101
rect 1856 4922 1857 5103
rect 2480 5102 2481 5573
rect 1856 5104 1857 5573
rect 2108 4922 2109 5105
rect 2108 5106 2109 5573
rect 2354 4922 2355 5107
rect 1475 4922 1476 5109
rect 2354 5108 2355 5573
rect 1474 5110 1475 5573
rect 2114 4922 2115 5111
rect 2114 5112 2115 5573
rect 3451 5112 3452 5573
rect 2402 5114 2403 5573
rect 3468 5114 3469 5573
rect 2420 5116 2421 5573
rect 2630 4922 2631 5117
rect 2426 5118 2427 5573
rect 2624 4922 2625 5119
rect 2444 4922 2445 5121
rect 3304 4922 3305 5121
rect 2444 5122 2445 5573
rect 2528 4922 2529 5123
rect 1994 4922 1995 5125
rect 2528 5124 2529 5573
rect 1994 5126 1995 5573
rect 2174 4922 2175 5127
rect 1889 5128 1890 5573
rect 2174 5128 2175 5573
rect 2450 5128 2451 5573
rect 2654 4922 2655 5129
rect 2462 5130 2463 5573
rect 2642 4922 2643 5131
rect 2468 4922 2469 5133
rect 3454 5132 3455 5573
rect 2024 4922 2025 5135
rect 2468 5134 2469 5573
rect 2024 5136 2025 5573
rect 2210 4922 2211 5137
rect 2210 5138 2211 5573
rect 2432 4922 2433 5139
rect 2432 5140 2433 5573
rect 2570 4922 2571 5141
rect 1880 4922 1881 5143
rect 2570 5142 2571 5573
rect 1880 5144 1881 5573
rect 2084 4922 2085 5145
rect 2084 5146 2085 5573
rect 2306 4922 2307 5147
rect 1507 4922 1508 5149
rect 2306 5148 2307 5573
rect 2504 5148 2505 5573
rect 2660 4922 2661 5149
rect 2186 4922 2187 5151
rect 2660 5150 2661 5573
rect 2120 4922 2121 5153
rect 2186 5152 2187 5573
rect 2120 5154 2121 5573
rect 3323 4922 3324 5155
rect 2510 5156 2511 5573
rect 2666 4922 2667 5157
rect 1541 5158 1542 5573
rect 2666 5158 2667 5573
rect 2540 5160 2541 5573
rect 3333 4922 3334 5161
rect 2552 4922 2553 5163
rect 3381 4922 3382 5163
rect 2552 5164 2553 5573
rect 2684 4922 2685 5165
rect 2564 5164 2565 5573
rect 2564 4922 2565 5165
rect 2576 4922 2577 5167
rect 3458 5166 3459 5573
rect 2576 5168 2577 5573
rect 2672 4922 2673 5169
rect 1940 4922 1941 5171
rect 2672 5170 2673 5573
rect 1940 5172 1941 5573
rect 2318 4922 2319 5173
rect 2318 5174 2319 5573
rect 2582 4922 2583 5175
rect 2048 4922 2049 5177
rect 2582 5176 2583 5573
rect 2048 5178 2049 5573
rect 2414 4922 2415 5179
rect 2414 5180 2415 5573
rect 3367 4922 3368 5181
rect 2618 4922 2619 5183
rect 3370 4922 3371 5183
rect 2030 4922 2031 5185
rect 2618 5184 2619 5573
rect 2030 5186 2031 5573
rect 2378 4922 2379 5187
rect 2378 5188 2379 5573
rect 2606 4922 2607 5189
rect 2606 5190 2607 5573
rect 2708 4922 2709 5191
rect 2624 5192 2625 5573
rect 2738 4922 2739 5193
rect 2630 5194 2631 5573
rect 2714 4922 2715 5195
rect 2642 5196 2643 5573
rect 2678 4922 2679 5197
rect 2654 5198 2655 5573
rect 2732 4922 2733 5199
rect 1850 4922 1851 5201
rect 2732 5200 2733 5573
rect 1424 4922 1425 5203
rect 1850 5202 1851 5573
rect 1423 5204 1424 5573
rect 1556 5204 1557 5573
rect 2678 5204 2679 5573
rect 2780 4922 2781 5205
rect 1512 5206 1513 5573
rect 2780 5206 2781 5573
rect 2684 5208 2685 5573
rect 3307 4922 3308 5209
rect 2708 5210 2709 5573
rect 2798 4922 2799 5211
rect 2714 5212 2715 5573
rect 2792 4922 2793 5213
rect 2738 5214 2739 5573
rect 2828 4922 2829 5215
rect 2744 4922 2745 5217
rect 3407 5216 3408 5573
rect 2744 5218 2745 5573
rect 2834 4922 2835 5219
rect 2762 4922 2763 5221
rect 3429 5220 3430 5573
rect 2762 5222 2763 5573
rect 2852 4922 2853 5223
rect 2768 4922 2769 5225
rect 3363 4922 3364 5225
rect 2756 4922 2757 5227
rect 2768 5226 2769 5573
rect 2792 5226 2793 5573
rect 2864 4922 2865 5227
rect 2798 5228 2799 5573
rect 2876 4922 2877 5229
rect 1500 4922 1501 5231
rect 2876 5230 2877 5573
rect 1494 4922 1495 5233
rect 1500 5232 1501 5573
rect 2810 5232 2811 5573
rect 2810 4922 2811 5233
rect 2816 4922 2817 5233
rect 3461 5232 3462 5573
rect 1946 4922 1947 5235
rect 2816 5234 2817 5573
rect 1946 5236 1947 5573
rect 2324 4922 2325 5237
rect 2324 5238 2325 5573
rect 2588 4922 2589 5239
rect 2054 4922 2055 5241
rect 2588 5240 2589 5573
rect 2054 5242 2055 5573
rect 3465 5242 3466 5573
rect 2828 5244 2829 5573
rect 2900 4922 2901 5245
rect 2834 5246 2835 5573
rect 2906 4922 2907 5247
rect 2846 5248 2847 5573
rect 2888 4922 2889 5249
rect 2750 4922 2751 5251
rect 2888 5250 2889 5573
rect 2750 5252 2751 5573
rect 2840 4922 2841 5253
rect 1916 4922 1917 5255
rect 2840 5254 2841 5573
rect 1916 5256 1917 5573
rect 2270 4922 2271 5257
rect 2270 5258 2271 5573
rect 2516 4922 2517 5259
rect 2000 4922 2001 5261
rect 2516 5260 2517 5573
rect 2000 5262 2001 5573
rect 2384 4922 2385 5263
rect 1427 4922 1428 5265
rect 2384 5264 2385 5573
rect 1426 5266 1427 5573
rect 1877 5266 1878 5573
rect 2852 5266 2853 5573
rect 2894 4922 2895 5267
rect 2858 4922 2859 5269
rect 3400 5268 3401 5573
rect 2858 5270 2859 5573
rect 2930 4922 2931 5271
rect 1898 4922 1899 5273
rect 2930 5272 2931 5573
rect 1898 5274 1899 5573
rect 2222 4922 2223 5275
rect 2222 5276 2223 5573
rect 2252 4922 2253 5277
rect 2252 5278 2253 5573
rect 3327 5278 3328 5573
rect 2864 5280 2865 5573
rect 2936 4922 2937 5281
rect 2870 4922 2871 5283
rect 3444 5282 3445 5573
rect 2870 5284 2871 5573
rect 2912 4922 2913 5285
rect 2894 5286 2895 5573
rect 2948 4922 2949 5287
rect 1706 4922 1707 5289
rect 2948 5288 2949 5573
rect 1706 5290 1707 5573
rect 1730 4922 1731 5291
rect 1730 5292 1731 5573
rect 2321 4922 2322 5293
rect 2900 5292 2901 5573
rect 2954 4922 2955 5293
rect 1832 4922 1833 5295
rect 2954 5294 2955 5573
rect 1431 4922 1432 5297
rect 1832 5296 1833 5573
rect 1430 5298 1431 5573
rect 1538 5298 1539 5573
rect 2912 5298 2913 5573
rect 2966 4922 2967 5299
rect 2921 4922 2922 5301
rect 3107 5300 3108 5573
rect 2924 4922 2925 5303
rect 3240 4922 3241 5303
rect 2918 4922 2919 5305
rect 2924 5304 2925 5573
rect 2918 5306 2919 5573
rect 3237 4922 3238 5307
rect 2942 4922 2943 5309
rect 3384 4922 3385 5309
rect 1964 4922 1965 5311
rect 2942 5310 2943 5573
rect 1964 5312 1965 5573
rect 2198 4922 2199 5313
rect 2078 4922 2079 5315
rect 2198 5314 2199 5573
rect 2078 5316 2079 5573
rect 2330 4922 2331 5317
rect 2096 4922 2097 5319
rect 2330 5318 2331 5573
rect 2096 5320 2097 5573
rect 2456 4922 2457 5321
rect 2456 5322 2457 5573
rect 2558 4922 2559 5323
rect 2558 5324 2559 5573
rect 2636 4922 2637 5325
rect 2636 5326 2637 5573
rect 2702 4922 2703 5327
rect 2702 5328 2703 5573
rect 2774 4922 2775 5329
rect 2774 5330 2775 5573
rect 2804 4922 2805 5331
rect 2804 5332 2805 5573
rect 2882 4922 2883 5333
rect 2696 4922 2697 5335
rect 2882 5334 2883 5573
rect 2696 5336 2697 5573
rect 3323 5336 3324 5573
rect 2960 5338 2961 5573
rect 3002 4922 3003 5339
rect 1712 4922 1713 5341
rect 3002 5340 3003 5573
rect 1712 5342 1713 5573
rect 1736 4922 1737 5343
rect 1664 4922 1665 5345
rect 1736 5344 1737 5573
rect 2963 5344 2964 5573
rect 3005 4922 3006 5345
rect 2966 5346 2967 5573
rect 2972 4922 2973 5347
rect 1808 4922 1809 5349
rect 2972 5348 2973 5573
rect 1808 5350 1809 5573
rect 1958 4922 1959 5351
rect 1958 5352 1959 5573
rect 2336 4922 2337 5353
rect 2336 5354 2337 5573
rect 2522 4922 2523 5355
rect 2066 4922 2067 5357
rect 2522 5356 2523 5573
rect 2066 5358 2067 5573
rect 2168 4922 2169 5359
rect 2168 5360 2169 5573
rect 2246 4922 2247 5361
rect 2246 5362 2247 5573
rect 2498 4922 2499 5363
rect 1928 4922 1929 5365
rect 2498 5364 2499 5573
rect 1928 5366 1929 5573
rect 2258 4922 2259 5367
rect 2258 5368 2259 5573
rect 2546 4922 2547 5369
rect 2546 5370 2547 5573
rect 2690 4922 2691 5371
rect 2690 5372 2691 5573
rect 2786 4922 2787 5373
rect 2786 5374 2787 5573
rect 3447 5374 3448 5573
rect 2981 5376 2982 5573
rect 3023 4922 3024 5377
rect 2429 4922 2430 5379
rect 3023 5378 3024 5573
rect 2984 5380 2985 5573
rect 3026 4922 3027 5381
rect 1778 4922 1779 5383
rect 3026 5382 3027 5573
rect 1444 5384 1445 5573
rect 1778 5384 1779 5573
rect 2999 4922 3000 5385
rect 3221 5384 3222 5573
rect 3014 5386 3015 5573
rect 3056 4922 3057 5387
rect 3032 4922 3033 5389
rect 3146 5388 3147 5573
rect 1796 4922 1797 5391
rect 3032 5390 3033 5573
rect 1796 5392 1797 5573
rect 1826 4922 1827 5393
rect 1826 5394 1827 5573
rect 2042 4922 2043 5395
rect 2042 5396 2043 5573
rect 2372 4922 2373 5397
rect 2372 5398 2373 5573
rect 2612 4922 2613 5399
rect 2612 5400 2613 5573
rect 2726 4922 2727 5401
rect 2726 5402 2727 5573
rect 2822 4922 2823 5403
rect 1515 5404 1516 5573
rect 2822 5404 2823 5573
rect 3050 4922 3051 5405
rect 3374 4922 3375 5405
rect 1820 4922 1821 5407
rect 3050 5406 3051 5573
rect 1820 5408 1821 5573
rect 2036 4922 2037 5409
rect 2036 5410 2037 5573
rect 2390 4922 2391 5411
rect 2162 4922 2163 5413
rect 2390 5412 2391 5573
rect 1485 4922 1486 5415
rect 2162 5414 2163 5573
rect 1484 5416 1485 5573
rect 1676 4922 1677 5417
rect 1676 5418 1677 5573
rect 3422 5418 3423 5573
rect 3056 5420 3057 5573
rect 3068 4922 3069 5421
rect 3068 5422 3069 5573
rect 3297 4922 3298 5423
rect 3092 5422 3093 5573
rect 3092 4922 3093 5423
rect 3095 5422 3096 5573
rect 3095 4922 3096 5423
rect 3098 4922 3099 5425
rect 3140 5424 3141 5573
rect 3116 4922 3117 5427
rect 3419 5426 3420 5573
rect 3104 4922 3105 5429
rect 3116 5428 3117 5573
rect 1700 4922 1701 5431
rect 3104 5430 3105 5573
rect 1700 5432 1701 5573
rect 1724 4922 1725 5433
rect 1724 5434 1725 5573
rect 1772 4922 1773 5435
rect 1417 4922 1418 5437
rect 1772 5436 1773 5573
rect 3170 4922 3171 5437
rect 3278 5436 3279 5573
rect 3170 5438 3171 5573
rect 3311 4922 3312 5439
rect 3182 5440 3183 5573
rect 3314 4922 3315 5441
rect 3188 4922 3189 5443
rect 3248 5442 3249 5573
rect 3128 4922 3129 5445
rect 3188 5444 3189 5573
rect 3038 4922 3039 5447
rect 3128 5446 3129 5573
rect 1437 5448 1438 5573
rect 3038 5448 3039 5573
rect 3203 4922 3204 5449
rect 3263 5448 3264 5573
rect 3206 4922 3207 5451
rect 3266 5450 3267 5573
rect 3158 4922 3159 5453
rect 3206 5452 3207 5573
rect 3134 4922 3135 5455
rect 3158 5454 3159 5573
rect 3044 4922 3045 5457
rect 3134 5456 3135 5573
rect 1802 4922 1803 5459
rect 3044 5458 3045 5573
rect 1802 5460 1803 5573
rect 1934 4922 1935 5461
rect 1441 4922 1442 5463
rect 1934 5462 1935 5573
rect 1440 5464 1441 5573
rect 2012 4922 2013 5465
rect 2012 5466 2013 5573
rect 2396 4922 2397 5467
rect 2396 5468 2397 5573
rect 3426 5468 3427 5573
rect 3212 4922 3213 5471
rect 3308 5470 3309 5573
rect 3164 4922 3165 5473
rect 3212 5472 3213 5573
rect 3122 4922 3123 5475
rect 3164 5474 3165 5573
rect 3080 4922 3081 5477
rect 3122 5476 3123 5573
rect 3074 4922 3075 5479
rect 3080 5478 3081 5573
rect 3062 4922 3063 5481
rect 3074 5480 3075 5573
rect 1522 5482 1523 5573
rect 3062 5482 3063 5573
rect 3215 4922 3216 5483
rect 3311 5482 3312 5573
rect 3218 4922 3219 5485
rect 3314 5484 3315 5573
rect 2996 4922 2997 5487
rect 3218 5486 3219 5573
rect 1814 4922 1815 5489
rect 2996 5488 2997 5573
rect 1529 5490 1530 5573
rect 1814 5490 1815 5573
rect 3224 4922 3225 5491
rect 3296 5490 3297 5573
rect 3176 4922 3177 5493
rect 3224 5492 3225 5573
rect 3236 5492 3237 5573
rect 3377 4922 3378 5493
rect 3243 4922 3244 5495
rect 3333 5494 3334 5573
rect 3251 5496 3252 5573
rect 3395 4922 3396 5497
rect 2990 4922 2991 5499
rect 3396 5498 3397 5573
rect 2990 5500 2991 5573
rect 3393 5500 3394 5573
rect 3273 4922 3274 5503
rect 3369 5502 3370 5573
rect 3272 5504 3273 5573
rect 3300 4922 3301 5505
rect 3276 4922 3277 5507
rect 3372 5506 3373 5573
rect 3194 4922 3195 5509
rect 3275 5508 3276 5573
rect 3194 5510 3195 5573
rect 3197 4922 3198 5511
rect 3285 4922 3286 5511
rect 3381 5510 3382 5573
rect 3230 4922 3231 5513
rect 3284 5512 3285 5573
rect 3191 4922 3192 5515
rect 3230 5514 3231 5573
rect 3288 4922 3289 5515
rect 3384 5514 3385 5573
rect 3317 4922 3318 5517
rect 3413 5516 3414 5573
rect 3320 4922 3321 5519
rect 3339 5518 3340 5573
rect 2720 4922 2721 5521
rect 3320 5520 3321 5573
rect 1922 4922 1923 5523
rect 2720 5522 2721 5573
rect 1922 5524 1923 5573
rect 2276 4922 2277 5525
rect 2276 5526 2277 5573
rect 2486 4922 2487 5527
rect 2486 5528 2487 5573
rect 2534 4922 2535 5529
rect 2534 5530 2535 5573
rect 2648 4922 2649 5531
rect 2438 4922 2439 5533
rect 2648 5532 2649 5573
rect 2018 4922 2019 5535
rect 2438 5534 2439 5573
rect 1886 5536 1887 5573
rect 2018 5536 2019 5573
rect 3330 4922 3331 5537
rect 3398 4922 3399 5537
rect 2936 5538 2937 5573
rect 3330 5538 3331 5573
rect 3336 4922 3337 5539
rect 3441 5538 3442 5573
rect 3342 4922 3343 5541
rect 3438 5540 3439 5573
rect 3354 4922 3355 5543
rect 3391 4922 3392 5543
rect 3294 4922 3295 5545
rect 3390 5544 3391 5573
rect 3357 4922 3358 5547
rect 3388 4922 3389 5547
rect 3261 4922 3262 5549
rect 3357 5548 3358 5573
rect 3200 4922 3201 5551
rect 3260 5550 3261 5573
rect 3152 4922 3153 5553
rect 3200 5552 3201 5573
rect 3110 4922 3111 5555
rect 3152 5554 3153 5573
rect 3008 4922 3009 5557
rect 3110 5556 3111 5573
rect 2978 4922 2979 5559
rect 3008 5558 3009 5573
rect 2978 5560 2979 5573
rect 3020 4922 3021 5561
rect 1784 4922 1785 5563
rect 3020 5562 3021 5573
rect 1784 5564 1785 5573
rect 1892 4922 1893 5565
rect 1420 4922 1421 5567
rect 1892 5566 1893 5573
rect 3291 4922 3292 5567
rect 3387 5566 3388 5573
rect 3233 4922 3234 5569
rect 3290 5568 3291 5573
rect 3360 4922 3361 5569
rect 3416 5568 3417 5573
rect 3403 5570 3404 5573
rect 3410 5570 3411 5573
rect 1420 5579 1421 6172
rect 1832 5577 1833 5580
rect 1423 5577 1424 5582
rect 1919 5581 1920 6172
rect 1433 5577 1434 5584
rect 1907 5577 1908 5584
rect 1434 5585 1435 6172
rect 1694 5577 1695 5586
rect 1437 5577 1438 5588
rect 1967 5587 1968 6172
rect 1438 5589 1439 6172
rect 2780 5577 2781 5590
rect 1440 5577 1441 5592
rect 2594 5577 2595 5592
rect 1441 5593 1442 6172
rect 1592 5577 1593 5594
rect 1444 5577 1445 5596
rect 1652 5577 1653 5596
rect 1445 5597 1446 6172
rect 1580 5577 1581 5598
rect 1456 5577 1457 5600
rect 1457 5599 1458 6172
rect 1462 5577 1463 5600
rect 1463 5599 1464 6172
rect 1468 5577 1469 5600
rect 1469 5599 1470 6172
rect 1481 5577 1482 5600
rect 2573 5577 2574 5600
rect 1482 5601 1483 6172
rect 2180 5577 2181 5602
rect 1477 5577 1478 5604
rect 2180 5603 2181 6172
rect 1484 5577 1485 5606
rect 2567 5605 2568 6172
rect 1488 5577 1489 5608
rect 2246 5577 2247 5608
rect 1500 5577 1501 5610
rect 1501 5609 1502 6172
rect 1515 5577 1516 5610
rect 2996 5577 2997 5610
rect 1519 5577 1520 5612
rect 1556 5577 1557 5612
rect 1522 5577 1523 5614
rect 3020 5577 3021 5614
rect 1532 5615 1533 6172
rect 1658 5577 1659 5616
rect 1535 5617 1536 6172
rect 1652 5617 1653 6172
rect 1541 5577 1542 5620
rect 2672 5577 2673 5620
rect 1544 5577 1545 5622
rect 1550 5621 1551 6172
rect 1544 5623 1545 6172
rect 2768 5577 2769 5624
rect 1547 5625 1548 6172
rect 2234 5577 2235 5626
rect 1556 5627 1557 6172
rect 1562 5577 1563 5628
rect 1568 5627 1569 6172
rect 1877 5577 1878 5628
rect 1580 5629 1581 6172
rect 1586 5577 1587 5630
rect 1592 5629 1593 6172
rect 1604 5577 1605 5630
rect 1604 5631 1605 6172
rect 1889 5577 1890 5632
rect 1426 5577 1427 5634
rect 1889 5633 1890 6172
rect 1427 5635 1428 6172
rect 1874 5577 1875 5636
rect 1616 5637 1617 6172
rect 1622 5577 1623 5638
rect 1622 5639 1623 6172
rect 1628 5577 1629 5640
rect 1598 5577 1599 5642
rect 1628 5641 1629 6172
rect 1598 5643 1599 6172
rect 1610 5577 1611 5644
rect 1430 5577 1431 5646
rect 1610 5645 1611 6172
rect 1646 5645 1647 6172
rect 1646 5577 1647 5646
rect 1664 5645 1665 6172
rect 1676 5577 1677 5646
rect 1676 5647 1677 6172
rect 1688 5577 1689 5648
rect 1682 5649 1683 6172
rect 1700 5577 1701 5650
rect 1688 5651 1689 6172
rect 1706 5577 1707 5652
rect 1694 5653 1695 6172
rect 1712 5577 1713 5654
rect 1700 5655 1701 6172
rect 1730 5577 1731 5656
rect 1712 5657 1713 6172
rect 1724 5577 1725 5658
rect 1526 5577 1527 5660
rect 1724 5659 1725 6172
rect 1525 5661 1526 6172
rect 2072 5577 2073 5662
rect 1718 5663 1719 6172
rect 1766 5577 1767 5664
rect 1730 5665 1731 6172
rect 1742 5577 1743 5666
rect 1742 5667 1743 6172
rect 1748 5577 1749 5668
rect 1670 5577 1671 5670
rect 1748 5669 1749 6172
rect 1754 5577 1755 5670
rect 3396 5577 3397 5670
rect 1754 5671 1755 6172
rect 2876 5577 2877 5672
rect 1760 5671 1761 6172
rect 1760 5577 1761 5672
rect 1766 5673 1767 6172
rect 1796 5577 1797 5674
rect 1736 5577 1737 5676
rect 1796 5675 1797 6172
rect 1431 5677 1432 6172
rect 1736 5677 1737 6172
rect 1772 5677 1773 6172
rect 1772 5577 1773 5678
rect 1778 5677 1779 6172
rect 1778 5577 1779 5678
rect 1784 5677 1785 6172
rect 1784 5577 1785 5678
rect 1790 5677 1791 6172
rect 1790 5577 1791 5678
rect 1802 5677 1803 6172
rect 1802 5577 1803 5678
rect 1808 5577 1809 5678
rect 1832 5677 1833 6172
rect 1485 5679 1486 6172
rect 1808 5679 1809 6172
rect 1814 5679 1815 6172
rect 1814 5577 1815 5680
rect 1820 5679 1821 6172
rect 1820 5577 1821 5680
rect 1826 5679 1827 6172
rect 1826 5577 1827 5680
rect 1829 5679 1830 6172
rect 1829 5577 1830 5680
rect 1838 5679 1839 6172
rect 1838 5577 1839 5680
rect 1844 5679 1845 6172
rect 1844 5577 1845 5680
rect 1850 5679 1851 6172
rect 1850 5577 1851 5680
rect 1868 5679 1869 6172
rect 2069 5577 2070 5680
rect 1874 5681 1875 6172
rect 1880 5577 1881 5682
rect 1880 5683 1881 6172
rect 2066 5577 2067 5684
rect 1886 5577 1887 5686
rect 2957 5685 2958 6172
rect 1424 5687 1425 6172
rect 1886 5687 1887 6172
rect 1925 5687 1926 6172
rect 1937 5577 1938 5688
rect 1952 5687 1953 6172
rect 1952 5577 1953 5688
rect 1988 5577 1989 5688
rect 3461 5577 3462 5688
rect 1940 5577 1941 5690
rect 1988 5689 1989 6172
rect 1928 5577 1929 5692
rect 1940 5691 1941 6172
rect 1928 5693 1929 6172
rect 1994 5577 1995 5694
rect 1946 5577 1947 5696
rect 1994 5695 1995 6172
rect 1922 5577 1923 5698
rect 1946 5697 1947 6172
rect 1910 5577 1911 5700
rect 1922 5699 1923 6172
rect 1898 5577 1899 5702
rect 1910 5701 1911 6172
rect 1417 5703 1418 6172
rect 1898 5703 1899 6172
rect 2033 5703 2034 6172
rect 2240 5577 2241 5704
rect 2042 5577 2043 5706
rect 2072 5705 2073 6172
rect 2030 5577 2031 5708
rect 2042 5707 2043 6172
rect 2120 5577 2121 5708
rect 3454 5577 3455 5708
rect 2090 5577 2091 5710
rect 2120 5709 2121 6172
rect 2054 5577 2055 5712
rect 2090 5711 2091 6172
rect 2036 5577 2037 5714
rect 2054 5713 2055 6172
rect 2036 5715 2037 6172
rect 2060 5577 2061 5716
rect 2012 5577 2013 5718
rect 2060 5717 2061 6172
rect 2012 5719 2013 6172
rect 2018 5577 2019 5720
rect 1970 5577 1971 5722
rect 2018 5721 2019 6172
rect 1489 5723 1490 6172
rect 1970 5723 1971 6172
rect 2204 5723 2205 6172
rect 2204 5577 2205 5724
rect 2234 5723 2235 6172
rect 2282 5577 2283 5724
rect 2228 5577 2229 5726
rect 2282 5725 2283 6172
rect 2186 5577 2187 5728
rect 2228 5727 2229 6172
rect 2240 5727 2241 6172
rect 2252 5577 2253 5728
rect 2246 5729 2247 6172
rect 2270 5577 2271 5730
rect 2252 5731 2253 6172
rect 2258 5577 2259 5732
rect 2258 5733 2259 6172
rect 2264 5577 2265 5734
rect 2264 5735 2265 6172
rect 3361 5735 3362 6172
rect 2270 5737 2271 6172
rect 2294 5577 2295 5738
rect 2276 5577 2277 5740
rect 3327 5577 3328 5740
rect 2276 5741 2277 6172
rect 2288 5577 2289 5742
rect 2198 5577 2199 5744
rect 2288 5743 2289 6172
rect 2198 5745 2199 6172
rect 2210 5577 2211 5746
rect 2210 5747 2211 6172
rect 2216 5577 2217 5748
rect 2156 5577 2157 5750
rect 2216 5749 2217 6172
rect 2144 5577 2145 5752
rect 2156 5751 2157 6172
rect 2114 5577 2115 5754
rect 2144 5753 2145 6172
rect 2084 5577 2085 5756
rect 2114 5755 2115 6172
rect 1474 5577 1475 5758
rect 2084 5757 2085 6172
rect 1475 5759 1476 6172
rect 2186 5759 2187 6172
rect 2294 5759 2295 6172
rect 2306 5577 2307 5760
rect 2300 5577 2301 5762
rect 3465 5577 3466 5762
rect 2300 5763 2301 6172
rect 2312 5577 2313 5764
rect 2306 5765 2307 6172
rect 2318 5577 2319 5766
rect 2312 5767 2313 6172
rect 2324 5577 2325 5768
rect 2318 5769 2319 6172
rect 2330 5577 2331 5770
rect 2324 5771 2325 6172
rect 2348 5577 2349 5772
rect 2330 5773 2331 6172
rect 2354 5577 2355 5774
rect 2333 5775 2334 6172
rect 2357 5577 2358 5776
rect 2336 5577 2337 5778
rect 3354 5777 3355 6172
rect 2336 5779 2337 6172
rect 2366 5577 2367 5780
rect 2348 5781 2349 6172
rect 2378 5577 2379 5782
rect 2354 5783 2355 6172
rect 2360 5577 2361 5784
rect 2360 5785 2361 6172
rect 2384 5577 2385 5786
rect 2366 5787 2367 6172
rect 2396 5577 2397 5788
rect 2378 5789 2379 6172
rect 2402 5577 2403 5790
rect 2384 5791 2385 6172
rect 3330 5577 3331 5792
rect 2390 5791 2391 6172
rect 2390 5577 2391 5792
rect 2396 5793 2397 6172
rect 2414 5577 2415 5794
rect 2402 5795 2403 6172
rect 2426 5577 2427 5796
rect 2408 5577 2409 5798
rect 2414 5797 2415 6172
rect 2408 5799 2409 6172
rect 3405 5799 3406 6172
rect 2420 5577 2421 5802
rect 3451 5577 3452 5802
rect 2222 5577 2223 5804
rect 3451 5803 3452 6172
rect 2192 5577 2193 5806
rect 2222 5805 2223 6172
rect 1478 5807 1479 6172
rect 2192 5807 2193 6172
rect 2420 5807 2421 6172
rect 2438 5577 2439 5808
rect 2426 5809 2427 6172
rect 2450 5577 2451 5810
rect 2438 5811 2439 6172
rect 2456 5577 2457 5812
rect 2450 5813 2451 6172
rect 2468 5577 2469 5814
rect 2456 5815 2457 6172
rect 2474 5577 2475 5816
rect 2468 5817 2469 6172
rect 3323 5577 3324 5818
rect 2474 5819 2475 6172
rect 2492 5577 2493 5820
rect 2486 5577 2487 5822
rect 3320 5577 3321 5822
rect 2486 5823 2487 6172
rect 3395 5823 3396 6172
rect 2492 5825 2493 6172
rect 2504 5577 2505 5826
rect 2504 5827 2505 6172
rect 2516 5577 2517 5828
rect 2516 5829 2517 6172
rect 2528 5577 2529 5830
rect 2528 5831 2529 6172
rect 2540 5577 2541 5832
rect 2540 5833 2541 6172
rect 2552 5577 2553 5834
rect 2582 5833 2583 6172
rect 2582 5577 2583 5834
rect 2591 5833 2592 6172
rect 2879 5577 2880 5834
rect 2594 5835 2595 6172
rect 2618 5577 2619 5836
rect 2606 5577 2607 5838
rect 2618 5837 2619 6172
rect 2606 5839 2607 6172
rect 2648 5577 2649 5840
rect 2630 5839 2631 6172
rect 2630 5577 2631 5840
rect 2636 5839 2637 6172
rect 2636 5577 2637 5840
rect 2642 5839 2643 6172
rect 2642 5577 2643 5840
rect 2648 5841 2649 6172
rect 2666 5577 2667 5842
rect 2654 5841 2655 6172
rect 2654 5577 2655 5842
rect 2672 5841 2673 6172
rect 2678 5577 2679 5842
rect 2678 5843 2679 6172
rect 2684 5577 2685 5844
rect 2684 5845 2685 6172
rect 2690 5577 2691 5846
rect 2690 5847 2691 6172
rect 2702 5577 2703 5848
rect 2696 5577 2697 5850
rect 3365 5849 3366 6172
rect 2696 5851 2697 6172
rect 2708 5577 2709 5852
rect 2702 5853 2703 6172
rect 2714 5577 2715 5854
rect 2708 5855 2709 6172
rect 2720 5577 2721 5856
rect 2714 5857 2715 6172
rect 3468 5577 3469 5858
rect 2720 5859 2721 6172
rect 2726 5577 2727 5860
rect 2726 5861 2727 6172
rect 3407 5577 3408 5862
rect 2756 5863 2757 6172
rect 2762 5577 2763 5864
rect 2762 5865 2763 6172
rect 2774 5577 2775 5866
rect 2768 5867 2769 6172
rect 2822 5577 2823 5868
rect 2774 5869 2775 6172
rect 3403 5577 3404 5870
rect 2780 5871 2781 6172
rect 3447 5577 3448 5872
rect 2432 5577 2433 5874
rect 3448 5873 3449 6172
rect 2432 5875 2433 6172
rect 2444 5577 2445 5876
rect 2444 5877 2445 6172
rect 2462 5577 2463 5878
rect 2462 5879 2463 6172
rect 2480 5577 2481 5880
rect 2480 5881 2481 6172
rect 2498 5577 2499 5882
rect 2498 5883 2499 6172
rect 2510 5577 2511 5884
rect 2510 5885 2511 6172
rect 2522 5577 2523 5886
rect 2522 5887 2523 6172
rect 2534 5577 2535 5888
rect 2534 5889 2535 6172
rect 2546 5577 2547 5890
rect 2546 5891 2547 6172
rect 2558 5577 2559 5892
rect 2558 5893 2559 6172
rect 2564 5577 2565 5894
rect 2564 5895 2565 6172
rect 2570 5577 2571 5896
rect 2570 5897 2571 6172
rect 2576 5577 2577 5898
rect 1516 5899 1517 6172
rect 2576 5899 2577 6172
rect 2786 5577 2787 5900
rect 3429 5577 3430 5900
rect 2786 5901 2787 6172
rect 2798 5577 2799 5902
rect 2792 5577 2793 5904
rect 3444 5577 3445 5904
rect 2792 5905 2793 6172
rect 2804 5577 2805 5906
rect 1512 5577 1513 5908
rect 2804 5907 2805 6172
rect 1513 5909 1514 6172
rect 1904 5577 1905 5910
rect 1904 5911 1905 6172
rect 1934 5577 1935 5912
rect 1916 5577 1917 5914
rect 1934 5913 1935 6172
rect 1892 5577 1893 5916
rect 1916 5915 1917 6172
rect 1491 5577 1492 5918
rect 1892 5917 1893 6172
rect 1492 5919 1493 6172
rect 2600 5577 2601 5920
rect 2600 5921 2601 6172
rect 2612 5577 2613 5922
rect 2612 5923 2613 6172
rect 2624 5577 2625 5924
rect 2624 5925 2625 6172
rect 2660 5577 2661 5926
rect 1538 5577 1539 5928
rect 2660 5927 2661 6172
rect 2798 5927 2799 6172
rect 2816 5577 2817 5928
rect 2801 5929 2802 6172
rect 3023 5577 3024 5930
rect 2807 5931 2808 6172
rect 2825 5577 2826 5932
rect 2810 5577 2811 5934
rect 3400 5577 3401 5934
rect 2810 5935 2811 6172
rect 2828 5577 2829 5936
rect 2816 5937 2817 6172
rect 2834 5577 2835 5938
rect 2822 5939 2823 6172
rect 2840 5577 2841 5940
rect 2828 5941 2829 6172
rect 2846 5577 2847 5942
rect 2834 5943 2835 6172
rect 2852 5577 2853 5944
rect 2840 5945 2841 6172
rect 2858 5577 2859 5946
rect 2846 5947 2847 6172
rect 2864 5577 2865 5948
rect 2852 5949 2853 6172
rect 2870 5577 2871 5950
rect 2858 5951 2859 6172
rect 3026 5577 3027 5952
rect 2864 5953 2865 6172
rect 2882 5577 2883 5954
rect 2870 5955 2871 6172
rect 2888 5577 2889 5956
rect 2876 5957 2877 6172
rect 2894 5577 2895 5958
rect 2882 5959 2883 6172
rect 2900 5577 2901 5960
rect 2888 5961 2889 6172
rect 2963 5577 2964 5962
rect 2900 5963 2901 6172
rect 2912 5577 2913 5964
rect 2906 5965 2907 6172
rect 3351 5965 3352 6172
rect 2912 5967 2913 6172
rect 2918 5577 2919 5968
rect 2918 5969 2919 6172
rect 2924 5577 2925 5970
rect 2924 5971 2925 6172
rect 2930 5577 2931 5972
rect 2930 5973 2931 6172
rect 2936 5577 2937 5974
rect 2936 5975 2937 6172
rect 2942 5577 2943 5976
rect 2942 5977 2943 6172
rect 2972 5577 2973 5978
rect 2948 5577 2949 5980
rect 3444 5979 3445 6172
rect 2948 5981 2949 6172
rect 2954 5577 2955 5982
rect 2954 5983 2955 6172
rect 2960 5577 2961 5984
rect 2960 5985 2961 6172
rect 2966 5577 2967 5986
rect 2966 5987 2967 6172
rect 3032 5577 3033 5988
rect 2972 5989 2973 6172
rect 2978 5577 2979 5990
rect 2975 5991 2976 6172
rect 2981 5577 2982 5992
rect 2978 5993 2979 6172
rect 2984 5577 2985 5994
rect 2984 5995 2985 6172
rect 2990 5577 2991 5996
rect 2990 5997 2991 6172
rect 3393 5577 3394 5998
rect 2996 5999 2997 6172
rect 3044 5577 3045 6000
rect 3011 6001 3012 6172
rect 3035 5577 3036 6002
rect 3020 6003 3021 6172
rect 3062 5577 3063 6004
rect 3026 6005 3027 6172
rect 3068 5577 3069 6006
rect 3044 6007 3045 6172
rect 3074 5577 3075 6008
rect 3062 6009 3063 6172
rect 3110 5577 3111 6010
rect 3068 6011 3069 6172
rect 3095 5577 3096 6012
rect 3074 6013 3075 6172
rect 3092 5577 3093 6014
rect 3086 6015 3087 6172
rect 3128 5577 3129 6016
rect 3092 6017 3093 6172
rect 3116 5577 3117 6018
rect 3098 6019 3099 6172
rect 3134 5577 3135 6020
rect 3104 5577 3105 6022
rect 3110 6021 3111 6172
rect 3104 6023 3105 6172
rect 3140 5577 3141 6024
rect 3107 5577 3108 6026
rect 3113 6025 3114 6172
rect 3134 6025 3135 6172
rect 3182 5577 3183 6026
rect 3140 6027 3141 6172
rect 3188 5577 3189 6028
rect 3152 5577 3153 6030
rect 3422 5577 3423 6030
rect 2126 5577 2127 6032
rect 3423 6031 3424 6172
rect 2096 5577 2097 6034
rect 2126 6033 2127 6172
rect 2096 6035 2097 6172
rect 2150 5577 2151 6036
rect 2138 5577 2139 6038
rect 2150 6037 2151 6172
rect 2138 6039 2139 6172
rect 2162 5577 2163 6040
rect 2162 6041 2163 6172
rect 2168 5577 2169 6042
rect 2168 6043 2169 6172
rect 2174 5577 2175 6044
rect 1447 5577 1448 6046
rect 2174 6045 2175 6172
rect 1448 6047 1449 6172
rect 2552 6047 2553 6172
rect 3146 5577 3147 6048
rect 3152 6047 3153 6172
rect 3146 6049 3147 6172
rect 3194 5577 3195 6050
rect 3158 5577 3159 6052
rect 3402 6051 3403 6172
rect 3158 6053 3159 6172
rect 3206 5577 3207 6054
rect 3164 5577 3165 6056
rect 3282 6055 3283 6172
rect 3164 6057 3165 6172
rect 3200 5577 3201 6058
rect 3176 6059 3177 6172
rect 3224 5577 3225 6060
rect 3182 6061 3183 6172
rect 3230 5577 3231 6062
rect 3188 6063 3189 6172
rect 3430 6063 3431 6172
rect 3200 6065 3201 6172
rect 3248 5577 3249 6066
rect 3203 6067 3204 6172
rect 3251 5577 3252 6068
rect 3206 6069 3207 6172
rect 3218 5577 3219 6070
rect 3209 6071 3210 6172
rect 3221 5577 3222 6072
rect 3218 6073 3219 6172
rect 3260 5577 3261 6074
rect 3221 6075 3222 6172
rect 3263 5577 3264 6076
rect 3224 6077 3225 6172
rect 3266 5577 3267 6078
rect 3230 6079 3231 6172
rect 3272 5577 3273 6080
rect 2588 5577 2589 6082
rect 3272 6081 3273 6172
rect 2588 6083 2589 6172
rect 2732 5577 2733 6084
rect 2732 6085 2733 6172
rect 2738 5577 2739 6086
rect 2738 6087 2739 6172
rect 2744 5577 2745 6088
rect 2744 6089 2745 6172
rect 2750 5577 2751 6090
rect 3233 6089 3234 6172
rect 3275 5577 3276 6090
rect 1640 5577 1641 6092
rect 3275 6091 3276 6172
rect 1634 5577 1635 6094
rect 1640 6093 1641 6172
rect 3242 6093 3243 6172
rect 3284 5577 3285 6094
rect 3248 6095 3249 6172
rect 3290 5577 3291 6096
rect 3260 6097 3261 6172
rect 3308 5577 3309 6098
rect 3263 6099 3264 6172
rect 3311 5577 3312 6100
rect 3266 6101 3267 6172
rect 3314 5577 3315 6102
rect 3285 6103 3286 6172
rect 3333 5577 3334 6104
rect 3291 6105 3292 6172
rect 3339 5577 3340 6106
rect 2030 6107 2031 6172
rect 3339 6107 3340 6172
rect 3296 5577 3297 6110
rect 3398 6109 3399 6172
rect 3309 6111 3310 6172
rect 3357 5577 3358 6112
rect 2066 6113 2067 6172
rect 3358 6113 3359 6172
rect 3315 6115 3316 6172
rect 3384 5577 3385 6116
rect 3321 6117 3322 6172
rect 3369 5577 3370 6118
rect 2666 6119 2667 6172
rect 3368 6119 3369 6172
rect 3324 6121 3325 6172
rect 3372 5577 3373 6122
rect 3342 6123 3343 6172
rect 3381 5577 3382 6124
rect 3345 6125 3346 6172
rect 3387 5577 3388 6126
rect 3348 6127 3349 6172
rect 3390 5577 3391 6128
rect 3371 6129 3372 6172
rect 3413 5577 3414 6130
rect 3374 6131 3375 6172
rect 3416 5577 3417 6132
rect 3377 6133 3378 6172
rect 3434 6133 3435 6172
rect 3389 6135 3390 6172
rect 3419 5577 3420 6136
rect 2342 5577 2343 6138
rect 3420 6137 3421 6172
rect 2342 6139 2343 6172
rect 2372 5577 2373 6140
rect 2372 6141 2373 6172
rect 3426 5577 3427 6142
rect 3236 5577 3237 6144
rect 3427 6143 3428 6172
rect 3236 6145 3237 6172
rect 3278 5577 3279 6146
rect 3116 6147 3117 6172
rect 3279 6147 3280 6172
rect 3410 5577 3411 6148
rect 3458 5577 3459 6148
rect 3414 6149 3415 6172
rect 3438 5577 3439 6150
rect 3392 6151 3393 6172
rect 3437 6151 3438 6172
rect 3417 6153 3418 6172
rect 3441 5577 3442 6154
rect 3014 5577 3015 6156
rect 3441 6155 3442 6172
rect 3014 6157 3015 6172
rect 3038 5577 3039 6158
rect 3038 6159 3039 6172
rect 3050 5577 3051 6160
rect 3050 6161 3051 6172
rect 3056 5577 3057 6162
rect 3056 6163 3057 6172
rect 3080 5577 3081 6164
rect 3080 6165 3081 6172
rect 3122 5577 3123 6166
rect 3122 6167 3123 6172
rect 3170 5577 3171 6168
rect 3170 6169 3171 6172
rect 3212 5577 3213 6170
rect 1417 6176 1418 6179
rect 1850 6176 1851 6179
rect 1417 6180 1418 6809
rect 1513 6176 1514 6181
rect 1420 6176 1421 6183
rect 2186 6176 2187 6183
rect 1420 6184 1421 6809
rect 1668 6184 1669 6809
rect 1424 6176 1425 6187
rect 1812 6186 1813 6809
rect 1424 6188 1425 6809
rect 1604 6176 1605 6189
rect 1427 6176 1428 6191
rect 1482 6176 1483 6191
rect 1427 6192 1428 6809
rect 1598 6176 1599 6193
rect 1431 6176 1432 6195
rect 1674 6194 1675 6809
rect 1431 6196 1432 6809
rect 1692 6196 1693 6809
rect 1434 6176 1435 6199
rect 1730 6176 1731 6199
rect 1434 6200 1435 6809
rect 1441 6176 1442 6201
rect 1438 6176 1439 6203
rect 2166 6202 2167 6809
rect 1438 6204 1439 6809
rect 1686 6204 1687 6809
rect 1441 6206 1442 6809
rect 1742 6176 1743 6207
rect 1448 6176 1449 6209
rect 2288 6176 2289 6209
rect 1448 6210 1449 6809
rect 2844 6210 2845 6809
rect 1457 6176 1458 6213
rect 1475 6176 1476 6213
rect 1457 6214 1458 6809
rect 1463 6176 1464 6215
rect 1463 6216 1464 6809
rect 1469 6176 1470 6217
rect 1469 6218 1470 6809
rect 2807 6176 2808 6219
rect 1472 6220 1473 6809
rect 2636 6176 2637 6221
rect 1476 6222 1477 6809
rect 1746 6222 1747 6809
rect 1478 6176 1479 6225
rect 2438 6176 2439 6225
rect 1479 6226 1480 6809
rect 1628 6176 1629 6227
rect 1485 6176 1486 6229
rect 2522 6176 2523 6229
rect 1489 6176 1490 6231
rect 2546 6176 2547 6231
rect 1492 6176 1493 6233
rect 1766 6176 1767 6233
rect 1494 6234 1495 6809
rect 1501 6176 1502 6235
rect 1500 6236 1501 6809
rect 1644 6236 1645 6809
rect 1503 6238 1504 6809
rect 1700 6176 1701 6239
rect 1512 6240 1513 6809
rect 1547 6176 1548 6241
rect 1516 6176 1517 6243
rect 1889 6176 1890 6243
rect 1515 6244 1516 6809
rect 2180 6176 2181 6245
rect 1518 6246 1519 6809
rect 1550 6176 1551 6247
rect 1525 6176 1526 6249
rect 1676 6176 1677 6249
rect 1524 6250 1525 6809
rect 1556 6176 1557 6251
rect 1528 6176 1529 6253
rect 2096 6176 2097 6253
rect 1532 6176 1533 6255
rect 3011 6176 3012 6255
rect 1539 6256 1540 6809
rect 1770 6256 1771 6809
rect 1542 6258 1543 6809
rect 1580 6176 1581 6259
rect 1554 6260 1555 6809
rect 1592 6176 1593 6261
rect 1560 6262 1561 6809
rect 1610 6176 1611 6263
rect 1566 6264 1567 6809
rect 1616 6176 1617 6265
rect 1572 6266 1573 6809
rect 1622 6176 1623 6267
rect 1584 6268 1585 6809
rect 2726 6176 2727 6269
rect 1587 6270 1588 6809
rect 2804 6176 2805 6271
rect 1596 6272 1597 6809
rect 1646 6176 1647 6273
rect 1608 6274 1609 6809
rect 2648 6176 2649 6275
rect 1611 6276 1612 6809
rect 2340 6276 2341 6809
rect 1614 6278 1615 6809
rect 1664 6176 1665 6279
rect 1620 6280 1621 6809
rect 1682 6176 1683 6281
rect 1626 6282 1627 6809
rect 1688 6176 1689 6283
rect 1632 6284 1633 6809
rect 1694 6176 1695 6285
rect 1652 6176 1653 6287
rect 2033 6176 2034 6287
rect 1656 6288 1657 6809
rect 1712 6176 1713 6289
rect 1662 6290 1663 6809
rect 1724 6176 1725 6291
rect 1680 6292 1681 6809
rect 1736 6176 1737 6293
rect 1698 6294 1699 6809
rect 1718 6176 1719 6295
rect 1710 6296 1711 6809
rect 1754 6176 1755 6297
rect 1716 6298 1717 6809
rect 1796 6176 1797 6299
rect 1722 6300 1723 6809
rect 1790 6176 1791 6301
rect 1728 6302 1729 6809
rect 2564 6176 2565 6303
rect 1734 6304 1735 6809
rect 1760 6176 1761 6305
rect 1740 6306 1741 6809
rect 2474 6176 2475 6307
rect 1752 6308 1753 6809
rect 2456 6176 2457 6309
rect 1758 6310 1759 6809
rect 1772 6176 1773 6311
rect 1764 6312 1765 6809
rect 1778 6176 1779 6313
rect 1776 6314 1777 6809
rect 2360 6176 2361 6315
rect 1782 6316 1783 6809
rect 1784 6176 1785 6317
rect 1788 6316 1789 6809
rect 2462 6176 2463 6317
rect 1794 6318 1795 6809
rect 2588 6176 2589 6319
rect 1800 6320 1801 6809
rect 1868 6176 1869 6321
rect 1802 6176 1803 6323
rect 1836 6322 1837 6809
rect 1806 6324 1807 6809
rect 1808 6176 1809 6325
rect 1814 6176 1815 6325
rect 1818 6324 1819 6809
rect 1820 6176 1821 6325
rect 1842 6324 1843 6809
rect 1824 6326 1825 6809
rect 2292 6326 2293 6809
rect 1826 6176 1827 6329
rect 1848 6328 1849 6809
rect 1827 6330 1828 6809
rect 2540 6176 2541 6331
rect 1829 6176 1830 6333
rect 1851 6332 1852 6809
rect 1830 6334 1831 6809
rect 1832 6176 1833 6335
rect 1838 6176 1839 6335
rect 1854 6334 1855 6809
rect 1844 6176 1845 6337
rect 1890 6336 1891 6809
rect 1856 6176 1857 6339
rect 1878 6338 1879 6809
rect 1860 6340 1861 6809
rect 2798 6176 2799 6341
rect 1862 6176 1863 6343
rect 1884 6342 1885 6809
rect 1866 6344 1867 6809
rect 2216 6176 2217 6345
rect 1872 6346 1873 6809
rect 2222 6176 2223 6347
rect 1874 6176 1875 6349
rect 2016 6348 2017 6809
rect 1880 6176 1881 6351
rect 2088 6350 2089 6809
rect 1886 6176 1887 6353
rect 3451 6176 3452 6353
rect 1568 6176 1569 6355
rect 1887 6354 1888 6809
rect 1892 6176 1893 6355
rect 1950 6354 1951 6809
rect 1896 6356 1897 6809
rect 1916 6176 1917 6357
rect 1898 6176 1899 6359
rect 1908 6358 1909 6809
rect 1902 6360 1903 6809
rect 1910 6176 1911 6361
rect 1904 6176 1905 6363
rect 1938 6362 1939 6809
rect 1905 6364 1906 6809
rect 1919 6176 1920 6365
rect 1914 6366 1915 6809
rect 1940 6176 1941 6367
rect 1920 6368 1921 6809
rect 1922 6176 1923 6369
rect 1928 6176 1929 6369
rect 2082 6368 2083 6809
rect 1932 6370 1933 6809
rect 1934 6176 1935 6371
rect 1944 6370 1945 6809
rect 1946 6176 1947 6371
rect 1956 6370 1957 6809
rect 1958 6176 1959 6371
rect 1962 6370 1963 6809
rect 1970 6176 1971 6371
rect 1964 6176 1965 6373
rect 1980 6372 1981 6809
rect 1974 6374 1975 6809
rect 1994 6176 1995 6375
rect 1976 6176 1977 6377
rect 2064 6376 2065 6809
rect 1982 6176 1983 6379
rect 1992 6378 1993 6809
rect 1986 6380 1987 6809
rect 2000 6176 2001 6381
rect 1998 6382 1999 6809
rect 2018 6176 2019 6383
rect 1925 6176 1926 6385
rect 2019 6384 2020 6809
rect 1445 6176 1446 6387
rect 1926 6386 1927 6809
rect 1445 6388 1446 6809
rect 1952 6176 1953 6389
rect 2004 6388 2005 6809
rect 2006 6176 2007 6389
rect 2010 6388 2011 6809
rect 2012 6176 2013 6389
rect 2022 6388 2023 6809
rect 2024 6176 2025 6389
rect 2028 6388 2029 6809
rect 2048 6176 2049 6389
rect 2030 6176 2031 6391
rect 2234 6176 2235 6391
rect 2034 6392 2035 6809
rect 2072 6176 2073 6393
rect 2036 6176 2037 6395
rect 2070 6394 2071 6809
rect 2040 6396 2041 6809
rect 2060 6176 2061 6397
rect 2042 6176 2043 6399
rect 2052 6398 2053 6809
rect 2046 6400 2047 6809
rect 2054 6176 2055 6401
rect 2058 6400 2059 6809
rect 3361 6176 3362 6401
rect 2066 6176 2067 6403
rect 3402 6176 3403 6403
rect 2076 6404 2077 6809
rect 2090 6176 2091 6405
rect 1967 6176 1968 6407
rect 2091 6406 2092 6809
rect 1968 6408 1969 6809
rect 1988 6176 1989 6409
rect 2078 6176 2079 6409
rect 3227 6408 3228 6809
rect 2084 6176 2085 6411
rect 2160 6410 2161 6809
rect 2094 6412 2095 6809
rect 2102 6176 2103 6413
rect 2100 6414 2101 6809
rect 2108 6176 2109 6415
rect 2106 6416 2107 6809
rect 2114 6176 2115 6417
rect 2112 6418 2113 6809
rect 2126 6176 2127 6419
rect 2118 6420 2119 6809
rect 2144 6176 2145 6421
rect 2120 6176 2121 6423
rect 3289 6422 3290 6809
rect 2124 6424 2125 6809
rect 3423 6176 3424 6425
rect 2130 6426 2131 6809
rect 2132 6176 2133 6427
rect 2136 6426 2137 6809
rect 2192 6176 2193 6427
rect 2138 6176 2139 6429
rect 2172 6428 2173 6809
rect 2142 6430 2143 6809
rect 2156 6176 2157 6431
rect 2148 6432 2149 6809
rect 2150 6176 2151 6433
rect 2154 6432 2155 6809
rect 2162 6176 2163 6433
rect 2168 6176 2169 6433
rect 2178 6432 2179 6809
rect 2174 6176 2175 6435
rect 2184 6434 2185 6809
rect 2181 6436 2182 6809
rect 2567 6176 2568 6437
rect 2190 6438 2191 6809
rect 2204 6176 2205 6439
rect 2196 6440 2197 6809
rect 2324 6176 2325 6441
rect 2198 6176 2199 6443
rect 2214 6442 2215 6809
rect 2202 6444 2203 6809
rect 2318 6176 2319 6445
rect 2208 6446 2209 6809
rect 2210 6176 2211 6447
rect 2220 6446 2221 6809
rect 2228 6176 2229 6447
rect 2223 6448 2224 6809
rect 2591 6176 2592 6449
rect 2226 6450 2227 6809
rect 2294 6176 2295 6451
rect 2232 6452 2233 6809
rect 2300 6176 2301 6453
rect 2238 6454 2239 6809
rect 2354 6176 2355 6455
rect 2240 6176 2241 6457
rect 2268 6456 2269 6809
rect 2244 6458 2245 6809
rect 2264 6176 2265 6459
rect 2246 6176 2247 6461
rect 2262 6460 2263 6809
rect 2250 6462 2251 6809
rect 2252 6176 2253 6463
rect 2256 6462 2257 6809
rect 2258 6176 2259 6463
rect 2270 6176 2271 6463
rect 2274 6462 2275 6809
rect 2276 6176 2277 6463
rect 2286 6462 2287 6809
rect 2282 6176 2283 6465
rect 2298 6464 2299 6809
rect 2304 6464 2305 6809
rect 2330 6176 2331 6465
rect 2306 6176 2307 6467
rect 2310 6466 2311 6809
rect 2307 6468 2308 6809
rect 2333 6176 2334 6469
rect 2312 6176 2313 6471
rect 2316 6470 2317 6809
rect 2322 6470 2323 6809
rect 2390 6176 2391 6471
rect 2328 6472 2329 6809
rect 3405 6176 3406 6473
rect 2334 6474 2335 6809
rect 2414 6176 2415 6475
rect 2336 6176 2337 6477
rect 2346 6476 2347 6809
rect 2337 6478 2338 6809
rect 2801 6176 2802 6479
rect 2342 6176 2343 6481
rect 3444 6176 3445 6481
rect 2348 6176 2349 6483
rect 2352 6482 2353 6809
rect 2358 6482 2359 6809
rect 2660 6176 2661 6483
rect 2364 6484 2365 6809
rect 2408 6176 2409 6485
rect 2366 6176 2367 6487
rect 2376 6486 2377 6809
rect 2370 6488 2371 6809
rect 2420 6176 2421 6489
rect 2372 6176 2373 6491
rect 2394 6490 2395 6809
rect 2378 6176 2379 6493
rect 2382 6492 2383 6809
rect 2384 6176 2385 6493
rect 3268 6492 3269 6809
rect 2396 6176 2397 6495
rect 2406 6494 2407 6809
rect 2400 6496 2401 6809
rect 2402 6176 2403 6497
rect 2412 6496 2413 6809
rect 3420 6176 3421 6497
rect 2418 6498 2419 6809
rect 3300 6498 3301 6809
rect 2424 6500 2425 6809
rect 2450 6176 2451 6501
rect 2426 6176 2427 6503
rect 2430 6502 2431 6809
rect 1640 6176 1641 6505
rect 2427 6504 2428 6809
rect 2432 6176 2433 6505
rect 2436 6504 2437 6809
rect 2442 6504 2443 6809
rect 2480 6176 2481 6505
rect 2444 6176 2445 6507
rect 2448 6506 2449 6809
rect 2454 6506 2455 6809
rect 2468 6176 2469 6507
rect 2460 6508 2461 6809
rect 2708 6176 2709 6509
rect 2466 6510 2467 6809
rect 2858 6176 2859 6511
rect 2472 6512 2473 6809
rect 2486 6176 2487 6513
rect 2478 6514 2479 6809
rect 2624 6176 2625 6515
rect 2484 6516 2485 6809
rect 2582 6176 2583 6517
rect 2490 6518 2491 6809
rect 2504 6176 2505 6519
rect 2492 6176 2493 6521
rect 3395 6176 3396 6521
rect 2496 6522 2497 6809
rect 2510 6176 2511 6523
rect 2498 6176 2499 6525
rect 3398 6176 3399 6525
rect 2502 6526 2503 6809
rect 2552 6176 2553 6527
rect 2508 6528 2509 6809
rect 2528 6176 2529 6529
rect 2514 6530 2515 6809
rect 2558 6176 2559 6531
rect 2516 6176 2517 6533
rect 2520 6532 2521 6809
rect 2526 6532 2527 6809
rect 2570 6176 2571 6533
rect 2532 6534 2533 6809
rect 2576 6176 2577 6535
rect 2534 6176 2535 6537
rect 3351 6176 3352 6537
rect 2538 6538 2539 6809
rect 3275 6176 3276 6539
rect 2544 6540 2545 6809
rect 2822 6176 2823 6541
rect 2550 6542 2551 6809
rect 2762 6176 2763 6543
rect 2556 6544 2557 6809
rect 2600 6176 2601 6545
rect 2562 6546 2563 6809
rect 3166 6546 3167 6809
rect 2568 6548 2569 6809
rect 2606 6176 2607 6549
rect 2574 6550 2575 6809
rect 2618 6176 2619 6551
rect 2580 6552 2581 6809
rect 2942 6176 2943 6553
rect 2586 6554 2587 6809
rect 2630 6176 2631 6555
rect 2592 6556 2593 6809
rect 2642 6176 2643 6557
rect 2594 6176 2595 6559
rect 3156 6558 3157 6809
rect 2598 6560 2599 6809
rect 2654 6176 2655 6561
rect 2604 6562 2605 6809
rect 2666 6176 2667 6563
rect 2610 6564 2611 6809
rect 2702 6176 2703 6565
rect 2616 6566 2617 6809
rect 2672 6176 2673 6567
rect 2622 6568 2623 6809
rect 2678 6176 2679 6569
rect 2628 6570 2629 6809
rect 2684 6176 2685 6571
rect 2634 6572 2635 6809
rect 2690 6176 2691 6573
rect 2640 6574 2641 6809
rect 3358 6176 3359 6575
rect 2646 6576 2647 6809
rect 2696 6176 2697 6577
rect 2652 6578 2653 6809
rect 3365 6176 3366 6579
rect 2658 6580 2659 6809
rect 3368 6176 3369 6581
rect 2664 6582 2665 6809
rect 2714 6176 2715 6583
rect 2670 6584 2671 6809
rect 2720 6176 2721 6585
rect 2676 6586 2677 6809
rect 2732 6176 2733 6587
rect 2682 6588 2683 6809
rect 2738 6176 2739 6589
rect 2688 6590 2689 6809
rect 2744 6176 2745 6591
rect 2706 6592 2707 6809
rect 2774 6176 2775 6593
rect 2712 6594 2713 6809
rect 2864 6176 2865 6595
rect 2718 6596 2719 6809
rect 2870 6176 2871 6597
rect 2724 6598 2725 6809
rect 2786 6176 2787 6599
rect 2730 6600 2731 6809
rect 2792 6176 2793 6601
rect 2736 6602 2737 6809
rect 2810 6176 2811 6603
rect 2742 6604 2743 6809
rect 2816 6176 2817 6605
rect 2748 6606 2749 6809
rect 2828 6176 2829 6607
rect 2754 6608 2755 6809
rect 2834 6176 2835 6609
rect 2766 6610 2767 6809
rect 2840 6176 2841 6611
rect 2772 6612 2773 6809
rect 2846 6176 2847 6613
rect 2778 6614 2779 6809
rect 2900 6176 2901 6615
rect 2784 6616 2785 6809
rect 2906 6176 2907 6617
rect 2790 6618 2791 6809
rect 2912 6176 2913 6619
rect 1535 6176 1536 6621
rect 2913 6620 2914 6809
rect 1536 6622 1537 6809
rect 2768 6176 2769 6623
rect 2796 6622 2797 6809
rect 2876 6176 2877 6623
rect 2802 6624 2803 6809
rect 2882 6176 2883 6625
rect 2808 6626 2809 6809
rect 2888 6176 2889 6627
rect 2820 6628 2821 6809
rect 2918 6176 2919 6629
rect 2826 6630 2827 6809
rect 2924 6176 2925 6631
rect 2832 6632 2833 6809
rect 2930 6176 2931 6633
rect 2838 6634 2839 6809
rect 2936 6176 2937 6635
rect 2850 6636 2851 6809
rect 2948 6176 2949 6637
rect 2856 6638 2857 6809
rect 2954 6176 2955 6639
rect 2859 6640 2860 6809
rect 2957 6176 2958 6641
rect 2862 6642 2863 6809
rect 2960 6176 2961 6643
rect 2868 6644 2869 6809
rect 2966 6176 2967 6645
rect 2874 6646 2875 6809
rect 2972 6176 2973 6647
rect 2877 6648 2878 6809
rect 3296 6648 3297 6809
rect 2880 6650 2881 6809
rect 2978 6176 2979 6651
rect 2886 6652 2887 6809
rect 2990 6176 2991 6653
rect 2892 6654 2893 6809
rect 3002 6176 3003 6655
rect 2898 6656 2899 6809
rect 2996 6176 2997 6657
rect 2904 6658 2905 6809
rect 3014 6176 3015 6659
rect 1748 6176 1749 6661
rect 3015 6660 3016 6809
rect 2910 6662 2911 6809
rect 3008 6176 3009 6663
rect 2916 6664 2917 6809
rect 3020 6176 3021 6665
rect 2922 6666 2923 6809
rect 3026 6176 3027 6667
rect 2928 6668 2929 6809
rect 3441 6176 3442 6669
rect 2940 6670 2941 6809
rect 3044 6176 3045 6671
rect 2946 6672 2947 6809
rect 3056 6176 3057 6673
rect 2952 6674 2953 6809
rect 3050 6176 3051 6675
rect 2958 6676 2959 6809
rect 3038 6176 3039 6677
rect 2964 6678 2965 6809
rect 3068 6176 3069 6679
rect 2970 6680 2971 6809
rect 3074 6176 3075 6681
rect 2975 6176 2976 6683
rect 3293 6682 3294 6809
rect 2976 6684 2977 6809
rect 3062 6176 3063 6685
rect 2982 6686 2983 6809
rect 3080 6176 3081 6687
rect 2988 6688 2989 6809
rect 3086 6176 3087 6689
rect 2994 6690 2995 6809
rect 3092 6176 3093 6691
rect 3000 6692 3001 6809
rect 3098 6176 3099 6693
rect 3006 6694 3007 6809
rect 3104 6176 3105 6695
rect 3012 6696 3013 6809
rect 3110 6176 3111 6697
rect 3018 6698 3019 6809
rect 3116 6176 3117 6699
rect 2852 6176 2853 6701
rect 3117 6700 3118 6809
rect 3024 6702 3025 6809
rect 3122 6176 3123 6703
rect 3036 6704 3037 6809
rect 3239 6704 3240 6809
rect 3048 6706 3049 6809
rect 3134 6176 3135 6707
rect 3054 6708 3055 6809
rect 3152 6176 3153 6709
rect 3060 6710 3061 6809
rect 3164 6176 3165 6711
rect 3066 6712 3067 6809
rect 3170 6176 3171 6713
rect 3078 6714 3079 6809
rect 3206 6176 3207 6715
rect 3081 6716 3082 6809
rect 3209 6176 3210 6717
rect 3090 6718 3091 6809
rect 3176 6176 3177 6719
rect 3102 6720 3103 6809
rect 3188 6176 3189 6721
rect 3105 6722 3106 6809
rect 3182 6176 3183 6723
rect 3108 6724 3109 6809
rect 3218 6176 3219 6725
rect 3111 6726 3112 6809
rect 3221 6176 3222 6727
rect 3113 6176 3114 6729
rect 3354 6176 3355 6729
rect 3114 6730 3115 6809
rect 3224 6176 3225 6731
rect 2780 6176 2781 6733
rect 3224 6732 3225 6809
rect 3120 6734 3121 6809
rect 3230 6176 3231 6735
rect 3123 6736 3124 6809
rect 3233 6176 3234 6737
rect 3126 6738 3127 6809
rect 3236 6176 3237 6739
rect 3030 6740 3031 6809
rect 3236 6740 3237 6809
rect 3132 6742 3133 6809
rect 3248 6176 3249 6743
rect 3140 6176 3141 6745
rect 3279 6176 3280 6745
rect 3144 6746 3145 6809
rect 3260 6176 3261 6747
rect 2756 6176 2757 6749
rect 3261 6748 3262 6809
rect 3146 6176 3147 6751
rect 3282 6176 3283 6751
rect 3147 6752 3148 6809
rect 3263 6176 3264 6753
rect 2700 6754 2701 6809
rect 3264 6754 3265 6809
rect 3150 6756 3151 6809
rect 3266 6176 3267 6757
rect 3158 6176 3159 6759
rect 3233 6758 3234 6809
rect 2984 6176 2985 6761
rect 3159 6760 3160 6809
rect 3163 6760 3164 6809
rect 3303 6760 3304 6809
rect 3169 6762 3170 6809
rect 3285 6176 3286 6763
rect 2280 6764 2281 6809
rect 3286 6764 3287 6809
rect 3181 6766 3182 6809
rect 3309 6176 3310 6767
rect 3187 6768 3188 6809
rect 3315 6176 3316 6769
rect 3193 6770 3194 6809
rect 3321 6176 3322 6771
rect 3196 6772 3197 6809
rect 3324 6176 3325 6773
rect 3200 6176 3201 6775
rect 3430 6176 3431 6775
rect 1544 6176 1545 6777
rect 3199 6776 3200 6809
rect 3203 6176 3204 6777
rect 3427 6176 3428 6777
rect 2612 6176 2613 6779
rect 3202 6778 3203 6809
rect 3211 6778 3212 6809
rect 3339 6176 3340 6779
rect 3214 6780 3215 6809
rect 3342 6176 3343 6781
rect 3217 6782 3218 6809
rect 3348 6176 3349 6783
rect 3220 6784 3221 6809
rect 3345 6176 3346 6785
rect 3230 6786 3231 6809
rect 3371 6176 3372 6787
rect 3242 6176 3243 6789
rect 3272 6176 3273 6789
rect 2388 6790 2389 6809
rect 3271 6790 3272 6809
rect 3243 6792 3244 6809
rect 3291 6176 3292 6793
rect 3246 6794 3247 6809
rect 3374 6176 3375 6795
rect 3255 6796 3256 6809
rect 3392 6176 3393 6797
rect 3258 6798 3259 6809
rect 3377 6176 3378 6799
rect 3280 6800 3281 6809
rect 3414 6176 3415 6801
rect 3283 6802 3284 6809
rect 3417 6176 3418 6803
rect 3389 6176 3390 6805
rect 3437 6176 3438 6805
rect 3434 6176 3435 6807
rect 3448 6176 3449 6807
rect 1427 6813 1428 6816
rect 1554 6813 1555 6816
rect 1434 6813 1435 6818
rect 1530 6817 1531 7370
rect 1438 6813 1439 6820
rect 1668 6813 1669 6820
rect 1441 6813 1442 6822
rect 1662 6813 1663 6822
rect 1445 6813 1446 6824
rect 2064 6813 2065 6824
rect 1448 6813 1449 6826
rect 1851 6813 1852 6826
rect 1454 6827 1455 7370
rect 1914 6813 1915 6828
rect 1472 6813 1473 6830
rect 1920 6813 1921 6830
rect 1476 6813 1477 6832
rect 2166 6813 2167 6832
rect 1417 6813 1418 6834
rect 1475 6833 1476 7370
rect 1479 6813 1480 6834
rect 2226 6813 2227 6834
rect 1478 6835 1479 7370
rect 2160 6813 2161 6836
rect 1482 6837 1483 7370
rect 2490 6813 2491 6838
rect 1503 6813 1504 6840
rect 1614 6813 1615 6840
rect 1512 6813 1513 6842
rect 2154 6813 2155 6842
rect 1512 6843 1513 7370
rect 2223 6813 2224 6844
rect 1536 6813 1537 6846
rect 2010 6813 2011 6846
rect 1524 6813 1525 6848
rect 1536 6847 1537 7370
rect 1518 6813 1519 6850
rect 1524 6849 1525 7370
rect 1542 6813 1543 6850
rect 1554 6849 1555 7370
rect 1548 6851 1549 7370
rect 2496 6813 2497 6852
rect 1551 6853 1552 7370
rect 1992 6813 1993 6854
rect 1566 6813 1567 6856
rect 1578 6855 1579 7370
rect 1424 6813 1425 6858
rect 1566 6857 1567 7370
rect 1599 6857 1600 7370
rect 2106 6813 2107 6858
rect 1608 6813 1609 6860
rect 1611 6813 1612 6860
rect 1596 6813 1597 6862
rect 1608 6861 1609 7370
rect 1596 6863 1597 7370
rect 1956 6813 1957 6864
rect 1469 6813 1470 6866
rect 1956 6865 1957 7370
rect 1463 6813 1464 6868
rect 1469 6867 1470 7370
rect 1457 6813 1458 6870
rect 1463 6869 1464 7370
rect 1620 6813 1621 6870
rect 1638 6869 1639 7370
rect 1620 6871 1621 7370
rect 2790 6813 2791 6872
rect 1623 6873 1624 7370
rect 2094 6813 2095 6874
rect 1632 6813 1633 6876
rect 1650 6875 1651 7370
rect 1644 6813 1645 6878
rect 1662 6877 1663 7370
rect 1626 6813 1627 6880
rect 1644 6879 1645 7370
rect 1500 6813 1501 6882
rect 1626 6881 1627 7370
rect 1494 6813 1495 6884
rect 1500 6883 1501 7370
rect 1674 6883 1675 7370
rect 1674 6813 1675 6884
rect 1680 6883 1681 7370
rect 1680 6813 1681 6884
rect 1686 6883 1687 7370
rect 1686 6813 1687 6884
rect 1698 6813 1699 6884
rect 1704 6883 1705 7370
rect 1692 6813 1693 6886
rect 1698 6885 1699 7370
rect 1431 6813 1432 6888
rect 1692 6887 1693 7370
rect 1430 6889 1431 7370
rect 1764 6813 1765 6890
rect 1722 6889 1723 7370
rect 1722 6813 1723 6890
rect 1749 6891 1750 7370
rect 2484 6813 2485 6892
rect 1764 6893 1765 7370
rect 1770 6813 1771 6894
rect 1433 6895 1434 7370
rect 1770 6895 1771 7370
rect 1836 6813 1837 6896
rect 3327 6895 3328 7370
rect 1836 6897 1837 7370
rect 1872 6813 1873 6898
rect 1740 6813 1741 6900
rect 1872 6899 1873 7370
rect 1423 6901 1424 7370
rect 1740 6901 1741 7370
rect 1866 6813 1867 6902
rect 1914 6901 1915 7370
rect 1806 6813 1807 6904
rect 1866 6903 1867 7370
rect 1788 6813 1789 6906
rect 1806 6905 1807 7370
rect 1776 6813 1777 6908
rect 1788 6907 1789 7370
rect 1758 6813 1759 6910
rect 1776 6909 1777 7370
rect 1746 6813 1747 6912
rect 1758 6911 1759 7370
rect 1887 6813 1888 6912
rect 1959 6911 1960 7370
rect 1905 6813 1906 6914
rect 1971 6913 1972 7370
rect 1656 6813 1657 6916
rect 1905 6915 1906 7370
rect 1920 6915 1921 7370
rect 2442 6813 2443 6916
rect 1950 6813 1951 6918
rect 1992 6917 1993 7370
rect 1878 6813 1879 6920
rect 1950 6919 1951 7370
rect 1728 6813 1729 6922
rect 1878 6921 1879 7370
rect 1728 6923 1729 7370
rect 1734 6813 1735 6924
rect 1426 6925 1427 7370
rect 1734 6925 1735 7370
rect 1980 6813 1981 6926
rect 2010 6925 2011 7370
rect 1938 6813 1939 6928
rect 1980 6927 1981 7370
rect 1884 6813 1885 6930
rect 1938 6929 1939 7370
rect 1884 6931 1885 7370
rect 3202 6813 3203 6932
rect 2001 6933 2002 7370
rect 2019 6813 2020 6934
rect 2025 6933 2026 7370
rect 2307 6813 2308 6934
rect 2034 6813 2035 6936
rect 2106 6935 2107 7370
rect 1962 6813 1963 6938
rect 2034 6937 2035 7370
rect 1902 6813 1903 6940
rect 1962 6939 1963 7370
rect 1848 6813 1849 6942
rect 1902 6941 1903 7370
rect 1812 6813 1813 6944
rect 1848 6943 1849 7370
rect 1800 6813 1801 6946
rect 1812 6945 1813 7370
rect 1800 6947 1801 7370
rect 3156 6813 3157 6948
rect 2043 6949 2044 7370
rect 2091 6813 2092 6950
rect 2058 6813 2059 6952
rect 2154 6951 2155 7370
rect 1974 6813 1975 6954
rect 2058 6953 2059 7370
rect 1974 6955 1975 7370
rect 2016 6813 2017 6956
rect 1944 6813 1945 6958
rect 2016 6957 2017 7370
rect 1944 6959 1945 7370
rect 2136 6813 2137 6960
rect 2040 6813 2041 6962
rect 2136 6961 2137 7370
rect 2040 6963 2041 7370
rect 2088 6813 2089 6964
rect 2064 6965 2065 7370
rect 3189 6965 3190 7370
rect 2070 6813 2071 6968
rect 2094 6967 2095 7370
rect 1986 6813 1987 6970
rect 2070 6969 2071 7370
rect 1908 6813 1909 6972
rect 1986 6971 1987 7370
rect 1437 6973 1438 7370
rect 1908 6973 1909 7370
rect 2100 6813 2101 6974
rect 2166 6973 2167 7370
rect 2004 6813 2005 6976
rect 2100 6975 2101 7370
rect 1932 6813 1933 6978
rect 2004 6977 2005 7370
rect 1890 6813 1891 6980
rect 1932 6979 1933 7370
rect 1854 6813 1855 6982
rect 1890 6981 1891 7370
rect 1440 6983 1441 7370
rect 1854 6983 1855 7370
rect 2112 6813 2113 6984
rect 3286 6813 3287 6984
rect 2022 6813 2023 6986
rect 2112 6985 2113 7370
rect 1451 6987 1452 7370
rect 2022 6987 2023 7370
rect 2130 6813 2131 6988
rect 2160 6987 2161 7370
rect 2046 6813 2047 6990
rect 2130 6989 2131 7370
rect 1420 6813 1421 6992
rect 2046 6991 2047 7370
rect 2181 6813 2182 6992
rect 2193 6991 2194 7370
rect 2184 6813 2185 6994
rect 2226 6993 2227 7370
rect 1485 6995 1486 7370
rect 2184 6995 2185 7370
rect 2235 6995 2236 7370
rect 3236 6813 3237 6996
rect 2280 6813 2281 6998
rect 3266 6997 3267 7370
rect 2280 6999 2281 7370
rect 2322 6813 2323 7000
rect 2286 6813 2287 7002
rect 2322 7001 2323 7370
rect 2250 6813 2251 7004
rect 2286 7003 2287 7370
rect 2190 6813 2191 7006
rect 2250 7005 2251 7370
rect 2178 6813 2179 7008
rect 2190 7007 2191 7370
rect 2178 7009 2179 7370
rect 3289 6813 3290 7010
rect 2310 6813 2311 7012
rect 3331 7011 3332 7370
rect 2262 6813 2263 7014
rect 2310 7013 2311 7370
rect 2214 6813 2215 7016
rect 2262 7015 2263 7370
rect 1515 6813 1516 7018
rect 2214 7017 2215 7370
rect 2316 6813 2317 7018
rect 3334 7017 3335 7370
rect 2274 6813 2275 7020
rect 2316 7019 2317 7370
rect 2274 7021 2275 7370
rect 2298 6813 2299 7022
rect 2244 6813 2245 7024
rect 2298 7023 2299 7370
rect 2232 6813 2233 7026
rect 2244 7025 2245 7370
rect 2220 6813 2221 7028
rect 2232 7027 2233 7370
rect 2142 6813 2143 7030
rect 2220 7029 2221 7370
rect 2052 6813 2053 7032
rect 2142 7031 2143 7370
rect 1968 6813 1969 7034
rect 2052 7033 2053 7370
rect 1896 6813 1897 7036
rect 1968 7035 1969 7370
rect 1842 6813 1843 7038
rect 1896 7037 1897 7370
rect 1842 7039 1843 7370
rect 2304 6813 2305 7040
rect 2268 6813 2269 7042
rect 2304 7041 2305 7370
rect 2268 7043 2269 7370
rect 2868 6813 2869 7044
rect 2337 6813 2338 7046
rect 2769 7045 2770 7370
rect 2358 6813 2359 7048
rect 3199 6813 3200 7048
rect 2340 6813 2341 7050
rect 2358 7049 2359 7370
rect 1827 6813 1828 7052
rect 2340 7051 2341 7370
rect 2391 7051 2392 7370
rect 2427 6813 2428 7052
rect 2406 6813 2407 7054
rect 2442 7053 2443 7370
rect 2376 6813 2377 7056
rect 2406 7055 2407 7370
rect 2352 6813 2353 7058
rect 2376 7057 2377 7370
rect 2328 6813 2329 7060
rect 2352 7059 2353 7370
rect 2292 6813 2293 7062
rect 2328 7061 2329 7370
rect 2256 6813 2257 7064
rect 2292 7063 2293 7370
rect 2238 6813 2239 7066
rect 2256 7065 2257 7370
rect 2208 6813 2209 7068
rect 2238 7067 2239 7370
rect 2118 6813 2119 7070
rect 2208 7069 2209 7370
rect 2118 7071 2119 7370
rect 2202 6813 2203 7072
rect 2124 6813 2125 7074
rect 2202 7073 2203 7370
rect 2028 6813 2029 7076
rect 2124 7075 2125 7370
rect 2028 7077 2029 7370
rect 2082 6813 2083 7078
rect 1998 6813 1999 7080
rect 2082 7079 2083 7370
rect 1926 6813 1927 7082
rect 1998 7081 1999 7370
rect 1926 7083 1927 7370
rect 3300 6813 3301 7084
rect 2448 6813 2449 7086
rect 3276 7085 3277 7370
rect 2418 6813 2419 7088
rect 2448 7087 2449 7370
rect 2394 6813 2395 7090
rect 2418 7089 2419 7370
rect 2364 6813 2365 7092
rect 2394 7091 2395 7370
rect 2364 7093 2365 7370
rect 2370 6813 2371 7094
rect 2346 6813 2347 7096
rect 2370 7095 2371 7370
rect 2334 6813 2335 7098
rect 2346 7097 2347 7370
rect 1824 6813 1825 7100
rect 2334 7099 2335 7370
rect 1824 7101 1825 7370
rect 1830 6813 1831 7102
rect 1521 7103 1522 7370
rect 1830 7103 1831 7370
rect 2472 6813 2473 7104
rect 2490 7103 2491 7370
rect 2454 6813 2455 7106
rect 2472 7105 2473 7370
rect 2436 6813 2437 7108
rect 2454 7107 2455 7370
rect 2412 6813 2413 7110
rect 2436 7109 2437 7370
rect 2382 6813 2383 7112
rect 2412 7111 2413 7370
rect 2382 7113 2383 7370
rect 3303 6813 3304 7114
rect 2478 6813 2479 7116
rect 3159 6813 3160 7116
rect 2478 7117 2479 7370
rect 2520 6813 2521 7118
rect 2484 7119 2485 7370
rect 3273 7119 3274 7370
rect 2496 7121 2497 7370
rect 2538 6813 2539 7122
rect 2502 6813 2503 7124
rect 2520 7123 2521 7370
rect 1584 6813 1585 7126
rect 2502 7125 2503 7370
rect 1572 6813 1573 7128
rect 1584 7127 1585 7370
rect 1560 6813 1561 7130
rect 1572 7129 1573 7370
rect 2514 7129 2515 7370
rect 2514 6813 2515 7130
rect 2526 6813 2527 7130
rect 2538 7129 2539 7370
rect 2526 7131 2527 7370
rect 2562 6813 2563 7132
rect 2466 6813 2467 7134
rect 2562 7133 2563 7370
rect 1746 7135 1747 7370
rect 2466 7135 2467 7370
rect 2568 6813 2569 7136
rect 3163 6813 3164 7136
rect 2568 7137 2569 7370
rect 3288 7137 3289 7370
rect 2574 6813 2575 7140
rect 3285 7139 3286 7370
rect 2556 6813 2557 7142
rect 2574 7141 2575 7370
rect 1587 6813 1588 7144
rect 2556 7143 2557 7370
rect 2586 7143 2587 7370
rect 2586 6813 2587 7144
rect 2616 6813 2617 7144
rect 3302 7143 3303 7370
rect 2616 7145 2617 7370
rect 2628 6813 2629 7146
rect 2628 7147 2629 7370
rect 2646 6813 2647 7148
rect 2646 7149 2647 7370
rect 2664 6813 2665 7150
rect 2658 7149 2659 7370
rect 2658 6813 2659 7150
rect 2664 7151 2665 7370
rect 2682 6813 2683 7152
rect 2676 6813 2677 7154
rect 3268 6813 3269 7154
rect 2676 7155 2677 7370
rect 3317 7155 3318 7370
rect 2688 7155 2689 7370
rect 2688 6813 2689 7156
rect 2694 7157 2695 7370
rect 3264 6813 3265 7158
rect 2712 6813 2713 7160
rect 2790 7159 2791 7370
rect 2712 7161 2713 7370
rect 2724 6813 2725 7162
rect 2706 6813 2707 7164
rect 2724 7163 2725 7370
rect 2706 7165 2707 7370
rect 3320 7165 3321 7370
rect 2748 7165 2749 7370
rect 2748 6813 2749 7166
rect 2754 7165 2755 7370
rect 2754 6813 2755 7166
rect 2760 7167 2761 7370
rect 3117 6813 3118 7168
rect 2808 7167 2809 7370
rect 2808 6813 2809 7168
rect 2838 6813 2839 7170
rect 2868 7169 2869 7370
rect 1447 7171 1448 7370
rect 2838 7171 2839 7370
rect 2859 6813 2860 7172
rect 2889 7171 2890 7370
rect 2862 6813 2863 7174
rect 3296 6813 3297 7174
rect 2832 6813 2833 7176
rect 2862 7175 2863 7370
rect 2778 6813 2779 7178
rect 2832 7177 2833 7370
rect 2772 6813 2773 7180
rect 2778 7179 2779 7370
rect 2766 6813 2767 7182
rect 2772 7181 2773 7370
rect 1860 6813 1861 7184
rect 2766 7183 2767 7370
rect 1818 6813 1819 7186
rect 1860 7185 1861 7370
rect 1518 7187 1519 7370
rect 1818 7187 1819 7370
rect 2877 6813 2878 7188
rect 2907 7187 2908 7370
rect 2886 6813 2887 7190
rect 3224 6813 3225 7190
rect 2856 6813 2857 7192
rect 2886 7191 2887 7370
rect 2826 6813 2827 7194
rect 2856 7193 2857 7370
rect 2718 6813 2719 7196
rect 2826 7195 2827 7370
rect 2544 6813 2545 7198
rect 2718 7197 2719 7370
rect 2532 6813 2533 7200
rect 2544 7199 2545 7370
rect 2508 6813 2509 7202
rect 2532 7201 2533 7370
rect 2508 7203 2509 7370
rect 2550 6813 2551 7204
rect 1444 7205 1445 7370
rect 2550 7205 2551 7370
rect 2895 7205 2896 7370
rect 2913 6813 2914 7206
rect 2904 6813 2905 7208
rect 2934 7207 2935 7370
rect 2874 6813 2875 7210
rect 2904 7209 2905 7370
rect 2844 6813 2845 7212
rect 2874 7211 2875 7370
rect 2784 6813 2785 7214
rect 2844 7213 2845 7370
rect 2580 6813 2581 7216
rect 2784 7215 2785 7370
rect 2580 7217 2581 7370
rect 2592 6813 2593 7218
rect 2592 7219 2593 7370
rect 2598 6813 2599 7220
rect 2598 7221 2599 7370
rect 2610 6813 2611 7222
rect 2610 7223 2611 7370
rect 2622 6813 2623 7224
rect 2622 7225 2623 7370
rect 2640 6813 2641 7226
rect 2640 7227 2641 7370
rect 2652 6813 2653 7228
rect 2652 7229 2653 7370
rect 2670 6813 2671 7230
rect 2670 7231 2671 7370
rect 2700 6813 2701 7232
rect 2700 7233 2701 7370
rect 2730 6813 2731 7234
rect 2730 7235 2731 7370
rect 2736 6813 2737 7236
rect 2736 7237 2737 7370
rect 2742 6813 2743 7238
rect 1539 6813 1540 7240
rect 2742 7239 2743 7370
rect 2940 6813 2941 7240
rect 3295 7239 3296 7370
rect 2898 6813 2899 7242
rect 2940 7241 2941 7370
rect 2892 6813 2893 7244
rect 2898 7243 2899 7370
rect 2892 7245 2893 7370
rect 2910 6813 2911 7246
rect 2880 6813 2881 7248
rect 2910 7247 2911 7370
rect 2850 6813 2851 7250
rect 2880 7249 2881 7370
rect 2820 6813 2821 7252
rect 2850 7251 2851 7370
rect 2802 6813 2803 7254
rect 2820 7253 2821 7370
rect 2796 6813 2797 7256
rect 2802 7255 2803 7370
rect 2796 7257 2797 7370
rect 3261 6813 3262 7258
rect 2964 6813 2965 7260
rect 2991 7259 2992 7370
rect 2946 6813 2947 7262
rect 2964 7261 2965 7370
rect 2916 6813 2917 7264
rect 2946 7263 2947 7370
rect 2916 7265 2917 7370
rect 3262 7265 3263 7370
rect 3006 6813 3007 7268
rect 3042 7267 3043 7370
rect 3006 7269 3007 7370
rect 3012 6813 3013 7270
rect 2982 6813 2983 7272
rect 3012 7271 3013 7370
rect 3009 7273 3010 7370
rect 3015 6813 3016 7274
rect 3030 6813 3031 7274
rect 3072 7273 3073 7370
rect 3030 7275 3031 7370
rect 3299 7275 3300 7370
rect 3036 6813 3037 7278
rect 3141 7277 3142 7370
rect 3000 6813 3001 7280
rect 3036 7279 3037 7370
rect 2958 6813 2959 7282
rect 3000 7281 3001 7370
rect 3048 6813 3049 7282
rect 3084 7281 3085 7370
rect 2976 6813 2977 7284
rect 3048 7283 3049 7370
rect 2922 6813 2923 7286
rect 2976 7285 2977 7370
rect 3066 6813 3067 7286
rect 3096 7285 3097 7370
rect 3024 6813 3025 7288
rect 3066 7287 3067 7370
rect 2994 6813 2995 7290
rect 3024 7289 3025 7370
rect 2994 7291 2995 7370
rect 3081 6813 3082 7292
rect 3078 6813 3079 7294
rect 3156 7293 3157 7370
rect 3105 6813 3106 7296
rect 3135 7295 3136 7370
rect 3108 6813 3109 7298
rect 3138 7297 3139 7370
rect 3111 6813 3112 7300
rect 3239 6813 3240 7300
rect 3123 6813 3124 7302
rect 3153 7301 3154 7370
rect 3132 6813 3133 7304
rect 3162 7303 3163 7370
rect 3102 6813 3103 7306
rect 3132 7305 3133 7370
rect 3102 7307 3103 7370
rect 3233 6813 3234 7308
rect 3144 6813 3145 7310
rect 3174 7309 3175 7370
rect 3147 6813 3148 7312
rect 3177 7311 3178 7370
rect 3159 7313 3160 7370
rect 3227 6813 3228 7314
rect 3166 6813 3167 7316
rect 3311 7315 3312 7370
rect 3169 6813 3170 7318
rect 3199 7317 3200 7370
rect 3181 6813 3182 7320
rect 3223 7319 3224 7370
rect 3150 6813 3151 7322
rect 3180 7321 3181 7370
rect 3120 6813 3121 7324
rect 3150 7323 3151 7370
rect 3090 6813 3091 7326
rect 3120 7325 3121 7370
rect 3060 6813 3061 7328
rect 3090 7327 3091 7370
rect 3054 6813 3055 7330
rect 3060 7329 3061 7370
rect 3018 6813 3019 7332
rect 3054 7331 3055 7370
rect 2988 6813 2989 7334
rect 3018 7333 3019 7370
rect 2970 6813 2971 7336
rect 2988 7335 2989 7370
rect 2952 6813 2953 7338
rect 2970 7337 2971 7370
rect 2928 6813 2929 7340
rect 2952 7339 2953 7370
rect 3193 6813 3194 7340
rect 3235 7339 3236 7370
rect 2922 7341 2923 7370
rect 3193 7341 3194 7370
rect 3196 6813 3197 7342
rect 3238 7341 3239 7370
rect 2928 7343 2929 7370
rect 3196 7343 3197 7370
rect 3205 7343 3206 7370
rect 3243 6813 3244 7344
rect 3114 6813 3115 7346
rect 3244 7345 3245 7370
rect 3211 6813 3212 7348
rect 3253 7347 3254 7370
rect 3217 6813 3218 7350
rect 3241 7349 3242 7370
rect 3220 6813 3221 7352
rect 3269 7351 3270 7370
rect 3255 6813 3256 7354
rect 3324 7353 3325 7370
rect 3214 6813 3215 7356
rect 3256 7355 3257 7370
rect 3258 6813 3259 7356
rect 3271 6813 3272 7356
rect 3126 6813 3127 7358
rect 3259 7357 3260 7370
rect 3280 6813 3281 7358
rect 3293 6813 3294 7358
rect 2958 7359 2959 7370
rect 3292 7359 3293 7370
rect 3230 6813 3231 7362
rect 3279 7361 3280 7370
rect 3187 6813 3188 7364
rect 3229 7363 3230 7370
rect 2088 7365 2089 7370
rect 3186 7365 3187 7370
rect 3283 6813 3284 7366
rect 3314 7365 3315 7370
rect 3246 6813 3247 7368
rect 3282 7367 3283 7370
rect 1423 7374 1424 7377
rect 1728 7374 1729 7377
rect 1423 7378 1424 8007
rect 1848 7374 1849 7379
rect 1430 7374 1431 7381
rect 1776 7374 1777 7381
rect 1433 7374 1434 7383
rect 1644 7374 1645 7383
rect 1437 7374 1438 7385
rect 1463 7374 1464 7385
rect 1438 7386 1439 8007
rect 1986 7374 1987 7387
rect 1444 7374 1445 7389
rect 1469 7374 1470 7389
rect 1445 7390 1446 8007
rect 1572 7374 1573 7391
rect 1447 7374 1448 7393
rect 2760 7374 2761 7393
rect 1449 7394 1450 8007
rect 1536 7374 1537 7395
rect 1451 7374 1452 7397
rect 2106 7374 2107 7397
rect 1452 7398 1453 8007
rect 1530 7374 1531 7399
rect 1454 7374 1455 7401
rect 1794 7374 1795 7401
rect 1461 7402 1462 8007
rect 1728 7402 1729 8007
rect 1464 7404 1465 8007
rect 1806 7374 1807 7405
rect 1468 7406 1469 8007
rect 1752 7374 1753 7407
rect 1475 7374 1476 7409
rect 1571 7408 1572 8007
rect 1478 7374 1479 7411
rect 2190 7374 2191 7411
rect 1480 7412 1481 8007
rect 1500 7374 1501 7413
rect 1482 7374 1483 7415
rect 1980 7374 1981 7415
rect 1485 7374 1486 7417
rect 2895 7374 2896 7417
rect 1492 7418 1493 8007
rect 3081 7418 3082 8007
rect 1504 7420 1505 8007
rect 1512 7374 1513 7421
rect 1510 7422 1511 8007
rect 1554 7374 1555 7423
rect 1442 7424 1443 8007
rect 1553 7424 1554 8007
rect 1513 7426 1514 8007
rect 2214 7374 2215 7427
rect 1518 7374 1519 7429
rect 2994 7374 2995 7429
rect 1517 7430 1518 8007
rect 1638 7374 1639 7431
rect 1521 7374 1522 7433
rect 1524 7374 1525 7433
rect 1523 7434 1524 8007
rect 1620 7374 1621 7435
rect 1551 7374 1552 7437
rect 2532 7374 2533 7437
rect 1559 7438 1560 8007
rect 1578 7374 1579 7439
rect 1580 7438 1581 8007
rect 2880 7374 2881 7439
rect 1589 7440 1590 8007
rect 1608 7374 1609 7441
rect 1599 7374 1600 7443
rect 2160 7374 2161 7443
rect 1602 7444 1603 8007
rect 2298 7374 2299 7445
rect 1605 7446 1606 8007
rect 2256 7374 2257 7447
rect 1614 7448 1615 8007
rect 1626 7374 1627 7449
rect 1623 7374 1624 7451
rect 2478 7374 2479 7451
rect 1626 7452 1627 8007
rect 1662 7374 1663 7453
rect 1644 7454 1645 8007
rect 3000 7374 3001 7455
rect 1656 7456 1657 8007
rect 2268 7374 2269 7457
rect 1662 7458 1663 8007
rect 2562 7374 2563 7459
rect 1520 7460 1521 8007
rect 2562 7460 2563 8007
rect 1668 7462 1669 8007
rect 1716 7374 1717 7463
rect 1692 7374 1693 7465
rect 1752 7464 1753 8007
rect 1710 7374 1711 7467
rect 2367 7466 2368 8007
rect 1686 7374 1687 7469
rect 1710 7468 1711 8007
rect 1650 7374 1651 7471
rect 1686 7470 1687 8007
rect 1650 7472 1651 8007
rect 3006 7374 3007 7473
rect 1716 7474 1717 8007
rect 3090 7374 3091 7475
rect 1746 7374 1747 7477
rect 2634 7374 2635 7477
rect 1746 7478 1747 8007
rect 2916 7374 2917 7479
rect 1749 7374 1750 7481
rect 2910 7374 2911 7481
rect 1776 7482 1777 8007
rect 2784 7374 2785 7483
rect 1782 7374 1783 7485
rect 1848 7484 1849 8007
rect 1782 7486 1783 8007
rect 2868 7374 2869 7487
rect 1794 7488 1795 8007
rect 2862 7374 2863 7489
rect 1806 7490 1807 8007
rect 2718 7374 2719 7491
rect 1824 7374 1825 7493
rect 1986 7492 1987 8007
rect 1722 7374 1723 7495
rect 1824 7494 1825 8007
rect 1722 7496 1723 8007
rect 2940 7374 2941 7497
rect 1896 7374 1897 7499
rect 2106 7498 2107 8007
rect 1788 7374 1789 7501
rect 1896 7500 1897 8007
rect 1471 7502 1472 8007
rect 1788 7502 1789 8007
rect 1905 7374 1906 7503
rect 2115 7502 2116 8007
rect 1959 7374 1960 7505
rect 2283 7504 2284 8007
rect 1974 7374 1975 7507
rect 2160 7506 2161 8007
rect 1974 7508 1975 8007
rect 2832 7374 2833 7509
rect 1980 7510 1981 8007
rect 2850 7374 2851 7511
rect 2001 7374 2002 7513
rect 2277 7512 2278 8007
rect 2016 7374 2017 7515
rect 2298 7514 2299 8007
rect 2016 7516 2017 8007
rect 2466 7374 2467 7517
rect 2025 7374 2026 7519
rect 2313 7518 2314 8007
rect 2028 7374 2029 7521
rect 2256 7520 2257 8007
rect 2028 7522 2029 8007
rect 2736 7374 2737 7523
rect 2043 7374 2044 7525
rect 2289 7524 2290 8007
rect 2100 7374 2101 7527
rect 3184 7526 3185 8007
rect 2100 7528 2101 8007
rect 2388 7374 2389 7529
rect 2088 7374 2089 7531
rect 2388 7530 2389 8007
rect 1890 7374 1891 7533
rect 2088 7532 2089 8007
rect 1764 7374 1765 7535
rect 1890 7534 1891 8007
rect 2190 7534 2191 8007
rect 2358 7374 2359 7535
rect 2064 7374 2065 7537
rect 2358 7536 2359 8007
rect 2064 7538 2065 8007
rect 2640 7374 2641 7539
rect 2193 7374 2194 7541
rect 2295 7540 2296 8007
rect 2208 7374 2209 7543
rect 2478 7542 2479 8007
rect 1950 7374 1951 7545
rect 2208 7544 2209 8007
rect 1812 7374 1813 7547
rect 1950 7546 1951 8007
rect 1812 7548 1813 8007
rect 1878 7374 1879 7549
rect 1818 7374 1819 7551
rect 1878 7550 1879 8007
rect 1548 7374 1549 7553
rect 1818 7552 1819 8007
rect 1547 7554 1548 8007
rect 1566 7374 1567 7555
rect 1565 7556 1566 8007
rect 1584 7374 1585 7557
rect 2214 7556 2215 8007
rect 2550 7374 2551 7557
rect 2235 7374 2236 7559
rect 2355 7558 2356 8007
rect 1971 7374 1972 7561
rect 2235 7560 2236 8007
rect 2238 7374 2239 7561
rect 2466 7560 2467 8007
rect 1992 7374 1993 7563
rect 2238 7562 2239 8007
rect 1836 7374 1837 7565
rect 1992 7564 1993 8007
rect 1598 7566 1599 8007
rect 1836 7566 1837 8007
rect 2244 7374 2245 7567
rect 3186 7374 3187 7567
rect 1440 7374 1441 7569
rect 2244 7568 2245 8007
rect 2268 7568 2269 8007
rect 2274 7374 2275 7569
rect 1998 7374 1999 7571
rect 2274 7570 2275 8007
rect 1842 7374 1843 7573
rect 1998 7572 1999 8007
rect 1758 7374 1759 7575
rect 1842 7574 1843 8007
rect 1698 7374 1699 7577
rect 1758 7576 1759 8007
rect 1698 7578 1699 8007
rect 1704 7374 1705 7579
rect 2286 7374 2287 7579
rect 2532 7578 2533 8007
rect 2004 7374 2005 7581
rect 2286 7580 2287 8007
rect 2004 7582 2005 8007
rect 2724 7374 2725 7583
rect 2316 7374 2317 7585
rect 3189 7374 3190 7585
rect 2316 7586 2317 8007
rect 2352 7374 2353 7587
rect 2052 7374 2053 7589
rect 2352 7588 2353 8007
rect 1854 7374 1855 7591
rect 2052 7590 2053 8007
rect 1426 7374 1427 7593
rect 1854 7592 1855 8007
rect 1426 7594 1427 8007
rect 1866 7374 1867 7595
rect 1740 7374 1741 7597
rect 1866 7596 1867 8007
rect 1680 7374 1681 7599
rect 1740 7598 1741 8007
rect 1680 7600 1681 8007
rect 2892 7374 2893 7601
rect 2337 7602 2338 8007
rect 2391 7374 2392 7603
rect 2361 7604 2362 8007
rect 2769 7374 2770 7605
rect 2406 7374 2407 7607
rect 3276 7374 3277 7607
rect 2166 7374 2167 7609
rect 2406 7608 2407 8007
rect 2166 7610 2167 8007
rect 2280 7374 2281 7611
rect 2280 7612 2281 8007
rect 3187 7612 3188 8007
rect 2412 7374 2413 7615
rect 3212 7614 3213 8007
rect 2124 7374 2125 7617
rect 2412 7616 2413 8007
rect 1926 7374 1927 7619
rect 2124 7618 2125 8007
rect 1926 7620 1927 8007
rect 2556 7374 2557 7621
rect 2394 7374 2395 7623
rect 2556 7622 2557 8007
rect 2130 7374 2131 7625
rect 2394 7624 2395 8007
rect 2076 7374 2077 7627
rect 2130 7626 2131 8007
rect 1914 7374 1915 7629
rect 2076 7628 2077 8007
rect 1914 7630 1915 8007
rect 2742 7374 2743 7631
rect 2454 7374 2455 7633
rect 2550 7632 2551 8007
rect 2322 7374 2323 7635
rect 2454 7634 2455 8007
rect 2034 7374 2035 7637
rect 2322 7636 2323 8007
rect 2034 7638 2035 8007
rect 3170 7638 3171 8007
rect 2460 7374 2461 7641
rect 3266 7374 3267 7641
rect 2172 7374 2173 7643
rect 2460 7642 2461 8007
rect 1938 7374 1939 7645
rect 2172 7644 2173 8007
rect 1938 7646 1939 8007
rect 2790 7374 2791 7647
rect 2472 7374 2473 7649
rect 3262 7374 3263 7649
rect 2202 7374 2203 7651
rect 2472 7650 2473 8007
rect 1956 7374 1957 7653
rect 2202 7652 2203 8007
rect 1920 7374 1921 7655
rect 1956 7654 1957 8007
rect 1920 7656 1921 8007
rect 2502 7374 2503 7657
rect 2340 7374 2341 7659
rect 2502 7658 2503 8007
rect 2046 7374 2047 7661
rect 2340 7660 2341 8007
rect 1435 7662 1436 8007
rect 2046 7662 2047 8007
rect 2490 7374 2491 7663
rect 2640 7662 2641 8007
rect 2262 7374 2263 7665
rect 2490 7664 2491 8007
rect 2040 7374 2041 7667
rect 2262 7666 2263 8007
rect 2040 7668 2041 8007
rect 2526 7374 2527 7669
rect 2508 7374 2509 7671
rect 3166 7670 3167 8007
rect 2304 7374 2305 7673
rect 2508 7672 2509 8007
rect 2094 7374 2095 7675
rect 2304 7674 2305 8007
rect 1908 7374 1909 7677
rect 2094 7676 2095 8007
rect 1770 7374 1771 7679
rect 1908 7678 1909 8007
rect 1770 7680 1771 8007
rect 2874 7374 2875 7681
rect 2514 7374 2515 7683
rect 3144 7682 3145 8007
rect 2514 7684 2515 8007
rect 2544 7374 2545 7685
rect 2310 7374 2311 7687
rect 2544 7686 2545 8007
rect 2022 7374 2023 7689
rect 2310 7688 2311 8007
rect 2022 7690 2023 8007
rect 2496 7374 2497 7691
rect 2250 7374 2251 7693
rect 2496 7692 2497 8007
rect 2010 7374 2011 7695
rect 2250 7694 2251 8007
rect 2010 7696 2011 8007
rect 2838 7374 2839 7697
rect 2526 7698 2527 8007
rect 3269 7374 3270 7699
rect 2538 7374 2539 7701
rect 2634 7700 2635 8007
rect 2292 7374 2293 7703
rect 2538 7702 2539 8007
rect 2184 7374 2185 7705
rect 2292 7704 2293 8007
rect 2184 7706 2185 8007
rect 2232 7374 2233 7707
rect 1968 7374 1969 7709
rect 2232 7708 2233 8007
rect 1968 7710 1969 8007
rect 3273 7374 3274 7711
rect 2610 7374 2611 7713
rect 3299 7374 3300 7713
rect 2424 7374 2425 7715
rect 2610 7714 2611 8007
rect 2136 7374 2137 7717
rect 2424 7716 2425 8007
rect 2118 7374 2119 7719
rect 2136 7718 2137 8007
rect 2118 7720 2119 8007
rect 2364 7374 2365 7721
rect 1596 7374 1597 7723
rect 2364 7722 2365 8007
rect 1595 7724 1596 8007
rect 2832 7724 2833 8007
rect 2616 7374 2617 7727
rect 3302 7374 3303 7727
rect 2436 7374 2437 7729
rect 2616 7728 2617 8007
rect 2196 7374 2197 7731
rect 2436 7730 2437 8007
rect 2196 7732 2197 8007
rect 2580 7374 2581 7733
rect 2370 7374 2371 7735
rect 2580 7734 2581 8007
rect 2646 7374 2647 7735
rect 2724 7734 2725 8007
rect 2664 7374 2665 7737
rect 2736 7736 2737 8007
rect 2568 7374 2569 7739
rect 2664 7738 2665 8007
rect 2568 7740 2569 8007
rect 3327 7374 3328 7741
rect 2670 7374 2671 7743
rect 2742 7742 2743 8007
rect 2670 7744 2671 8007
rect 3288 7374 3289 7745
rect 2682 7746 2683 8007
rect 3324 7374 3325 7747
rect 2688 7374 2689 7749
rect 3320 7374 3321 7749
rect 2574 7374 2575 7751
rect 2688 7750 2689 8007
rect 2520 7374 2521 7753
rect 2574 7752 2575 8007
rect 2484 7374 2485 7755
rect 2520 7754 2521 8007
rect 2220 7374 2221 7757
rect 2484 7756 2485 8007
rect 2148 7374 2149 7759
rect 2220 7758 2221 8007
rect 1932 7374 1933 7761
rect 2148 7760 2149 8007
rect 1932 7762 1933 8007
rect 2400 7374 2401 7763
rect 2142 7374 2143 7765
rect 2400 7764 2401 8007
rect 2142 7766 2143 8007
rect 3334 7374 3335 7767
rect 2694 7374 2695 7769
rect 3147 7768 3148 8007
rect 2604 7374 2605 7771
rect 2694 7770 2695 8007
rect 2604 7772 2605 8007
rect 3209 7772 3210 8007
rect 2700 7374 2701 7775
rect 2718 7774 2719 8007
rect 2622 7374 2623 7777
rect 2700 7776 2701 8007
rect 2442 7374 2443 7779
rect 2622 7778 2623 8007
rect 2334 7374 2335 7781
rect 2442 7780 2443 8007
rect 2058 7374 2059 7783
rect 2334 7782 2335 8007
rect 1860 7374 1861 7785
rect 2058 7784 2059 8007
rect 1734 7374 1735 7787
rect 1860 7786 1861 8007
rect 1674 7374 1675 7789
rect 1734 7788 1735 8007
rect 1577 7790 1578 8007
rect 1674 7790 1675 8007
rect 2706 7374 2707 7791
rect 2760 7790 2761 8007
rect 2628 7374 2629 7793
rect 2706 7792 2707 8007
rect 2448 7374 2449 7795
rect 2628 7794 2629 8007
rect 2178 7374 2179 7797
rect 2448 7796 2449 8007
rect 2178 7798 2179 8007
rect 2346 7374 2347 7799
rect 2070 7374 2071 7801
rect 2346 7800 2347 8007
rect 1884 7374 1885 7803
rect 2070 7802 2071 8007
rect 1800 7374 1801 7805
rect 1884 7804 1885 8007
rect 1800 7806 1801 8007
rect 2856 7374 2857 7807
rect 2754 7374 2755 7809
rect 3015 7808 3016 8007
rect 2784 7810 2785 8007
rect 2844 7374 2845 7811
rect 2790 7812 2791 8007
rect 2796 7374 2797 7813
rect 2772 7374 2773 7815
rect 2796 7814 2797 8007
rect 2748 7374 2749 7817
rect 2772 7816 2773 8007
rect 2676 7374 2677 7819
rect 2748 7818 2749 8007
rect 2586 7374 2587 7821
rect 2676 7820 2677 8007
rect 2376 7374 2377 7823
rect 2586 7822 2587 8007
rect 2112 7374 2113 7825
rect 2376 7824 2377 8007
rect 1902 7374 1903 7827
rect 2112 7826 2113 8007
rect 1830 7374 1831 7829
rect 1902 7828 1903 8007
rect 1830 7830 1831 8007
rect 1872 7374 1873 7831
rect 1872 7832 1873 8007
rect 2766 7374 2767 7833
rect 2712 7374 2713 7835
rect 2766 7834 2767 8007
rect 2658 7374 2659 7837
rect 2712 7836 2713 8007
rect 2592 7374 2593 7839
rect 2658 7838 2659 8007
rect 2418 7374 2419 7841
rect 2592 7840 2593 8007
rect 2328 7374 2329 7843
rect 2418 7842 2419 8007
rect 2226 7374 2227 7845
rect 2328 7844 2329 8007
rect 1962 7374 1963 7847
rect 2226 7846 2227 8007
rect 1962 7848 1963 8007
rect 3331 7374 3332 7849
rect 2814 7850 2815 8007
rect 2820 7374 2821 7851
rect 2835 7850 2836 8007
rect 3009 7374 3010 7851
rect 2838 7852 2839 8007
rect 2946 7374 2947 7853
rect 2844 7854 2845 8007
rect 2976 7374 2977 7855
rect 2850 7856 2851 8007
rect 2898 7374 2899 7857
rect 2856 7858 2857 8007
rect 2922 7374 2923 7859
rect 2862 7860 2863 8007
rect 2886 7374 2887 7861
rect 2865 7862 2866 8007
rect 2889 7374 2890 7863
rect 2868 7864 2869 8007
rect 2928 7374 2929 7865
rect 2874 7866 2875 8007
rect 3096 7374 3097 7867
rect 2880 7868 2881 8007
rect 2904 7374 2905 7869
rect 2883 7870 2884 8007
rect 2907 7374 2908 7871
rect 2886 7872 2887 8007
rect 3129 7872 3130 8007
rect 2892 7874 2893 8007
rect 3156 7374 3157 7875
rect 2895 7876 2896 8007
rect 3159 7374 3160 7877
rect 2898 7878 2899 8007
rect 3012 7374 3013 7879
rect 2904 7880 2905 8007
rect 2958 7374 2959 7881
rect 2910 7882 2911 8007
rect 2952 7374 2953 7883
rect 2916 7884 2917 8007
rect 3295 7374 3296 7885
rect 2922 7886 2923 8007
rect 2970 7374 2971 7887
rect 2928 7888 2929 8007
rect 3018 7374 3019 7889
rect 2934 7374 2935 7891
rect 3196 7374 3197 7891
rect 2940 7892 2941 8007
rect 2988 7374 2989 7893
rect 2943 7894 2944 8007
rect 2991 7374 2992 7895
rect 2946 7896 2947 8007
rect 3030 7374 3031 7897
rect 2952 7898 2953 8007
rect 3259 7374 3260 7899
rect 2958 7900 2959 8007
rect 3024 7374 3025 7901
rect 2964 7374 2965 7903
rect 3292 7374 3293 7903
rect 2964 7904 2965 8007
rect 3317 7374 3318 7905
rect 2970 7906 2971 8007
rect 3036 7374 3037 7907
rect 2976 7908 2977 8007
rect 3042 7374 3043 7909
rect 2982 7910 2983 8007
rect 3066 7374 3067 7911
rect 2370 7912 2371 8007
rect 3066 7912 3067 8007
rect 2988 7914 2989 8007
rect 3072 7374 3073 7915
rect 2994 7916 2995 8007
rect 3141 7374 3142 7917
rect 3000 7918 3001 8007
rect 3084 7374 3085 7919
rect 3006 7920 3007 8007
rect 3150 7374 3151 7921
rect 3009 7922 3010 8007
rect 3054 7374 3055 7923
rect 3012 7924 3013 8007
rect 3244 7374 3245 7925
rect 3018 7926 3019 8007
rect 3102 7374 3103 7927
rect 3030 7928 3031 8007
rect 3138 7374 3139 7929
rect 3033 7930 3034 8007
rect 3069 7930 3070 8007
rect 3036 7932 3037 8007
rect 3120 7374 3121 7933
rect 3048 7374 3049 7935
rect 3126 7934 3127 8007
rect 3048 7936 3049 8007
rect 3132 7374 3133 7937
rect 3051 7938 3052 8007
rect 3135 7374 3136 7939
rect 3054 7940 3055 8007
rect 3162 7374 3163 7941
rect 3060 7374 3061 7943
rect 3163 7942 3164 8007
rect 3060 7944 3061 8007
rect 3177 7374 3178 7945
rect 3063 7946 3064 8007
rect 3174 7374 3175 7947
rect 2730 7374 2731 7949
rect 3173 7948 3174 8007
rect 2652 7374 2653 7951
rect 2730 7950 2731 8007
rect 2652 7952 2653 8007
rect 3202 7952 3203 8007
rect 3072 7954 3073 8007
rect 3180 7374 3181 7955
rect 2646 7956 2647 8007
rect 3180 7956 3181 8007
rect 3078 7958 3079 8007
rect 3153 7374 3154 7959
rect 3084 7960 3085 8007
rect 3199 7374 3200 7961
rect 3096 7962 3097 8007
rect 3205 7374 3206 7963
rect 2382 7374 2383 7965
rect 3205 7964 3206 8007
rect 2082 7374 2083 7967
rect 2382 7966 2383 8007
rect 2082 7968 2083 8007
rect 2598 7374 2599 7969
rect 2430 7374 2431 7971
rect 2598 7970 2599 8007
rect 2154 7374 2155 7973
rect 2430 7972 2431 8007
rect 1944 7374 1945 7975
rect 2154 7974 2155 8007
rect 1944 7976 1945 8007
rect 2826 7374 2827 7977
rect 2808 7374 2809 7979
rect 2826 7978 2827 8007
rect 2802 7374 2803 7981
rect 2808 7980 2809 8007
rect 2778 7374 2779 7983
rect 2802 7982 2803 8007
rect 3108 7982 3109 8007
rect 3223 7374 3224 7983
rect 3114 7984 3115 8007
rect 3229 7374 3230 7985
rect 3120 7986 3121 8007
rect 3235 7374 3236 7987
rect 3123 7988 3124 8007
rect 3238 7374 3239 7989
rect 3138 7990 3139 8007
rect 3253 7374 3254 7991
rect 3141 7992 3142 8007
rect 3151 7992 3152 8007
rect 3154 7992 3155 8007
rect 3256 7374 3257 7993
rect 3157 7994 3158 8007
rect 3279 7374 3280 7995
rect 3160 7996 3161 8007
rect 3282 7374 3283 7997
rect 3177 7998 3178 8007
rect 3241 7374 3242 7999
rect 3193 7374 3194 8001
rect 3285 7374 3286 8001
rect 3196 8002 3197 8007
rect 3311 7374 3312 8003
rect 3199 8004 3200 8007
rect 3314 7374 3315 8005
rect 1423 8011 1424 8014
rect 1440 8013 1441 8586
rect 1423 8015 1424 8586
rect 2208 8011 2209 8016
rect 1426 8011 1427 8018
rect 2046 8011 2047 8018
rect 1430 8019 1431 8586
rect 1488 8019 1489 8586
rect 1433 8021 1434 8586
rect 1492 8011 1493 8022
rect 1438 8011 1439 8024
rect 1926 8011 1927 8024
rect 1445 8011 1446 8026
rect 2289 8011 2290 8026
rect 1444 8027 1445 8586
rect 2322 8011 2323 8028
rect 1452 8011 1453 8030
rect 1523 8011 1524 8030
rect 1454 8031 1455 8586
rect 1890 8011 1891 8032
rect 1461 8011 1462 8034
rect 1830 8011 1831 8034
rect 1464 8011 1465 8036
rect 1812 8011 1813 8036
rect 1463 8037 1464 8586
rect 1896 8011 1897 8038
rect 1437 8039 1438 8586
rect 1896 8039 1897 8586
rect 1466 8041 1467 8586
rect 1812 8041 1813 8586
rect 1468 8011 1469 8044
rect 1547 8011 1548 8044
rect 1471 8011 1472 8046
rect 1575 8045 1576 8586
rect 1480 8011 1481 8048
rect 1494 8047 1495 8586
rect 1504 8011 1505 8048
rect 1506 8047 1507 8586
rect 1510 8011 1511 8048
rect 2370 8011 2371 8048
rect 1520 8011 1521 8050
rect 2358 8011 2359 8050
rect 1524 8051 1525 8586
rect 1764 8051 1765 8586
rect 1527 8053 1528 8586
rect 1914 8011 1915 8054
rect 1548 8055 1549 8586
rect 1553 8011 1554 8056
rect 1554 8057 1555 8586
rect 1559 8011 1560 8058
rect 1560 8059 1561 8586
rect 1565 8011 1566 8060
rect 1566 8061 1567 8586
rect 1571 8011 1572 8062
rect 1572 8063 1573 8586
rect 1650 8011 1651 8064
rect 1577 8011 1578 8066
rect 3051 8011 3052 8066
rect 1584 8067 1585 8586
rect 1589 8011 1590 8068
rect 1590 8069 1591 8586
rect 1626 8011 1627 8070
rect 1593 8071 1594 8586
rect 3054 8011 3055 8072
rect 1595 8011 1596 8074
rect 1800 8011 1801 8074
rect 1598 8011 1599 8076
rect 1794 8011 1795 8076
rect 1602 8011 1603 8078
rect 2454 8011 2455 8078
rect 1602 8079 1603 8586
rect 1614 8011 1615 8080
rect 1614 8081 1615 8586
rect 1674 8011 1675 8082
rect 1620 8083 1621 8586
rect 1686 8011 1687 8084
rect 1638 8085 1639 8586
rect 1698 8011 1699 8086
rect 1650 8087 1651 8586
rect 1734 8011 1735 8088
rect 1656 8011 1657 8090
rect 1692 8089 1693 8586
rect 1656 8091 1657 8586
rect 1740 8011 1741 8092
rect 1662 8011 1663 8094
rect 1698 8093 1699 8586
rect 1662 8095 1663 8586
rect 1668 8011 1669 8096
rect 1668 8097 1669 8586
rect 1752 8011 1753 8098
rect 1674 8099 1675 8586
rect 1758 8011 1759 8100
rect 1686 8101 1687 8586
rect 1728 8011 1729 8102
rect 1704 8103 1705 8586
rect 1788 8011 1789 8104
rect 1716 8011 1717 8106
rect 2778 8105 2779 8586
rect 1716 8107 1717 8586
rect 1776 8011 1777 8108
rect 1722 8011 1723 8110
rect 2745 8109 2746 8586
rect 1722 8111 1723 8586
rect 1806 8011 1807 8112
rect 1451 8113 1452 8586
rect 1806 8113 1807 8586
rect 1728 8115 1729 8586
rect 1818 8011 1819 8116
rect 1734 8117 1735 8586
rect 1824 8011 1825 8118
rect 1740 8119 1741 8586
rect 1782 8011 1783 8120
rect 1752 8121 1753 8586
rect 1842 8011 1843 8122
rect 1758 8123 1759 8586
rect 1848 8011 1849 8124
rect 1776 8125 1777 8586
rect 1854 8011 1855 8126
rect 1782 8127 1783 8586
rect 1860 8011 1861 8128
rect 1788 8129 1789 8586
rect 1866 8011 1867 8130
rect 1794 8131 1795 8586
rect 1902 8011 1903 8132
rect 1800 8133 1801 8586
rect 1884 8011 1885 8134
rect 1818 8135 1819 8586
rect 1878 8011 1879 8136
rect 1824 8137 1825 8586
rect 1920 8011 1921 8138
rect 1830 8139 1831 8586
rect 1944 8011 1945 8140
rect 1842 8141 1843 8586
rect 1908 8011 1909 8142
rect 1836 8011 1837 8144
rect 1908 8143 1909 8586
rect 1836 8145 1837 8586
rect 1932 8011 1933 8146
rect 1848 8147 1849 8586
rect 1974 8011 1975 8148
rect 1854 8149 1855 8586
rect 1980 8011 1981 8150
rect 1860 8151 1861 8586
rect 2010 8011 2011 8152
rect 1866 8153 1867 8586
rect 2784 8011 2785 8154
rect 1878 8155 1879 8586
rect 1962 8011 1963 8156
rect 1884 8157 1885 8586
rect 1968 8011 1969 8158
rect 1890 8159 1891 8586
rect 1950 8011 1951 8160
rect 1902 8161 1903 8586
rect 2004 8011 2005 8162
rect 1473 8163 1474 8586
rect 2004 8163 2005 8586
rect 1914 8165 1915 8586
rect 2772 8011 2773 8166
rect 1926 8167 1927 8586
rect 2034 8011 2035 8168
rect 1932 8169 1933 8586
rect 3184 8011 3185 8170
rect 1944 8171 1945 8586
rect 1992 8011 1993 8172
rect 1950 8173 1951 8586
rect 1998 8011 1999 8174
rect 1962 8175 1963 8586
rect 2016 8011 2017 8176
rect 1968 8177 1969 8586
rect 2022 8011 2023 8178
rect 1974 8179 1975 8586
rect 2760 8011 2761 8180
rect 1980 8181 1981 8586
rect 2040 8011 2041 8182
rect 1992 8183 1993 8586
rect 2052 8011 2053 8184
rect 1998 8185 1999 8586
rect 2058 8011 2059 8186
rect 2010 8187 2011 8586
rect 2082 8011 2083 8188
rect 2016 8189 2017 8586
rect 2070 8011 2071 8190
rect 2022 8191 2023 8586
rect 2076 8011 2077 8192
rect 2028 8011 2029 8194
rect 3170 8011 3171 8194
rect 2028 8195 2029 8586
rect 2682 8011 2683 8196
rect 2034 8197 2035 8586
rect 2100 8011 2101 8198
rect 2040 8199 2041 8586
rect 2088 8011 2089 8200
rect 2046 8201 2047 8586
rect 2106 8011 2107 8202
rect 2052 8203 2053 8586
rect 2112 8011 2113 8204
rect 2055 8205 2056 8586
rect 2115 8011 2116 8206
rect 2058 8207 2059 8586
rect 2094 8011 2095 8208
rect 2064 8011 2065 8210
rect 3041 8209 3042 8586
rect 2064 8211 2065 8586
rect 2118 8011 2119 8212
rect 1447 8213 1448 8586
rect 2118 8213 2119 8586
rect 2070 8215 2071 8586
rect 2142 8011 2143 8216
rect 2076 8217 2077 8586
rect 2124 8011 2125 8218
rect 2082 8219 2083 8586
rect 2130 8011 2131 8220
rect 2088 8221 2089 8586
rect 2136 8011 2137 8222
rect 2094 8223 2095 8586
rect 2154 8011 2155 8224
rect 2100 8225 2101 8586
rect 2148 8011 2149 8226
rect 2106 8227 2107 8586
rect 2178 8011 2179 8228
rect 2112 8229 2113 8586
rect 2160 8011 2161 8230
rect 1580 8011 1581 8232
rect 2160 8231 2161 8586
rect 2124 8233 2125 8586
rect 2196 8011 2197 8234
rect 2130 8235 2131 8586
rect 2184 8011 2185 8236
rect 2136 8237 2137 8586
rect 3023 8237 3024 8586
rect 2142 8239 2143 8586
rect 2190 8011 2191 8240
rect 1426 8241 1427 8586
rect 2190 8241 2191 8586
rect 2148 8243 2149 8586
rect 2172 8011 2173 8244
rect 2154 8245 2155 8586
rect 2652 8011 2653 8246
rect 2166 8011 2167 8248
rect 3202 8011 3203 8248
rect 2166 8249 2167 8586
rect 2268 8011 2269 8250
rect 2172 8251 2173 8586
rect 2214 8011 2215 8252
rect 1435 8011 1436 8254
rect 2214 8253 2215 8586
rect 2178 8255 2179 8586
rect 2520 8011 2521 8256
rect 2184 8257 2185 8586
rect 2202 8011 2203 8258
rect 2196 8259 2197 8586
rect 2220 8011 2221 8260
rect 2202 8261 2203 8586
rect 2514 8011 2515 8262
rect 2208 8263 2209 8586
rect 2292 8011 2293 8264
rect 2220 8265 2221 8586
rect 2226 8011 2227 8266
rect 2226 8267 2227 8586
rect 2232 8011 2233 8268
rect 2229 8269 2230 8586
rect 2235 8011 2236 8270
rect 2232 8271 2233 8586
rect 2238 8011 2239 8272
rect 2238 8273 2239 8586
rect 2244 8011 2245 8274
rect 2244 8275 2245 8586
rect 2250 8011 2251 8276
rect 2250 8277 2251 8586
rect 2256 8011 2257 8278
rect 2256 8279 2257 8586
rect 2262 8011 2263 8280
rect 2262 8281 2263 8586
rect 2502 8011 2503 8282
rect 2268 8283 2269 8586
rect 2274 8011 2275 8284
rect 2271 8285 2272 8586
rect 2277 8011 2278 8286
rect 1442 8011 1443 8288
rect 2277 8287 2278 8586
rect 2274 8289 2275 8586
rect 2286 8011 2287 8290
rect 2280 8011 2281 8292
rect 2286 8291 2287 8586
rect 1515 8293 1516 8586
rect 2280 8293 2281 8586
rect 2283 8011 2284 8294
rect 2289 8293 2290 8586
rect 2292 8293 2293 8586
rect 2304 8011 2305 8294
rect 2298 8011 2299 8296
rect 2304 8295 2305 8586
rect 2298 8297 2299 8586
rect 2418 8011 2419 8298
rect 2313 8011 2314 8300
rect 2331 8299 2332 8586
rect 2316 8011 2317 8302
rect 3069 8011 3070 8302
rect 2316 8303 2317 8586
rect 2364 8011 2365 8304
rect 2319 8305 2320 8586
rect 3075 8305 3076 8586
rect 2322 8307 2323 8586
rect 2442 8011 2443 8308
rect 1605 8011 1606 8310
rect 2442 8309 2443 8586
rect 2337 8011 2338 8312
rect 2349 8311 2350 8586
rect 2295 8011 2296 8314
rect 2337 8313 2338 8586
rect 2346 8011 2347 8314
rect 2358 8313 2359 8586
rect 2334 8011 2335 8316
rect 2346 8315 2347 8586
rect 1470 8317 1471 8586
rect 2334 8317 2335 8586
rect 2352 8011 2353 8318
rect 2364 8317 2365 8586
rect 2340 8011 2341 8320
rect 2352 8319 2353 8586
rect 2340 8321 2341 8586
rect 2376 8011 2377 8322
rect 2361 8321 2362 8586
rect 2361 8011 2362 8322
rect 2370 8323 2371 8586
rect 2394 8011 2395 8324
rect 2376 8325 2377 8586
rect 2400 8011 2401 8326
rect 2382 8011 2383 8328
rect 2394 8327 2395 8586
rect 2382 8329 2383 8586
rect 2550 8011 2551 8330
rect 2400 8331 2401 8586
rect 2490 8011 2491 8332
rect 2418 8333 2419 8586
rect 2430 8011 2431 8334
rect 2424 8011 2425 8336
rect 2430 8335 2431 8586
rect 2412 8011 2413 8338
rect 2424 8337 2425 8586
rect 2412 8339 2413 8586
rect 3147 8011 3148 8340
rect 2448 8339 2449 8586
rect 2448 8011 2449 8340
rect 2454 8341 2455 8586
rect 2466 8011 2467 8342
rect 2460 8341 2461 8586
rect 2460 8011 2461 8342
rect 2466 8343 2467 8586
rect 2556 8011 2557 8344
rect 2472 8343 2473 8586
rect 2472 8011 2473 8344
rect 2478 8343 2479 8586
rect 2478 8011 2479 8344
rect 2484 8343 2485 8586
rect 2484 8011 2485 8344
rect 2490 8345 2491 8586
rect 2508 8011 2509 8346
rect 2496 8011 2497 8348
rect 2956 8347 2957 8586
rect 2496 8349 2497 8586
rect 2562 8011 2563 8350
rect 2502 8351 2503 8586
rect 2574 8011 2575 8352
rect 2508 8353 2509 8586
rect 2526 8011 2527 8354
rect 2514 8355 2515 8586
rect 2568 8011 2569 8356
rect 2520 8357 2521 8586
rect 2532 8011 2533 8358
rect 2526 8359 2527 8586
rect 2538 8011 2539 8360
rect 2532 8361 2533 8586
rect 2598 8011 2599 8362
rect 2538 8363 2539 8586
rect 3180 8011 3181 8364
rect 2544 8011 2545 8366
rect 3020 8365 3021 8586
rect 2544 8367 2545 8586
rect 2592 8011 2593 8368
rect 2550 8369 2551 8586
rect 2616 8011 2617 8370
rect 2556 8371 2557 8586
rect 2610 8011 2611 8372
rect 2562 8373 2563 8586
rect 2580 8011 2581 8374
rect 2568 8375 2569 8586
rect 2586 8011 2587 8376
rect 2574 8377 2575 8586
rect 2622 8011 2623 8378
rect 2586 8379 2587 8586
rect 2604 8011 2605 8380
rect 2592 8381 2593 8586
rect 2628 8011 2629 8382
rect 2604 8383 2605 8586
rect 2640 8011 2641 8384
rect 2610 8385 2611 8586
rect 2646 8011 2647 8386
rect 2616 8387 2617 8586
rect 2658 8011 2659 8388
rect 2622 8389 2623 8586
rect 2670 8011 2671 8390
rect 2628 8391 2629 8586
rect 2664 8011 2665 8392
rect 2640 8393 2641 8586
rect 2694 8011 2695 8394
rect 2646 8395 2647 8586
rect 2700 8011 2701 8396
rect 2652 8397 2653 8586
rect 2706 8011 2707 8398
rect 2658 8399 2659 8586
rect 2736 8011 2737 8400
rect 2664 8401 2665 8586
rect 2742 8011 2743 8402
rect 1746 8011 1747 8404
rect 2742 8403 2743 8586
rect 1746 8405 1747 8586
rect 1872 8011 1873 8406
rect 1872 8407 1873 8586
rect 1956 8011 1957 8408
rect 1956 8409 1957 8586
rect 2718 8011 2719 8410
rect 2670 8411 2671 8586
rect 2724 8011 2725 8412
rect 2682 8413 2683 8586
rect 2748 8011 2749 8414
rect 2694 8415 2695 8586
rect 2796 8011 2797 8416
rect 2700 8417 2701 8586
rect 2802 8011 2803 8418
rect 2706 8419 2707 8586
rect 2808 8011 2809 8420
rect 2724 8421 2725 8586
rect 2826 8011 2827 8422
rect 2733 8423 2734 8586
rect 2835 8011 2836 8424
rect 2736 8425 2737 8586
rect 2850 8011 2851 8426
rect 1517 8011 1518 8428
rect 2850 8427 2851 8586
rect 1449 8011 1450 8430
rect 1518 8429 1519 8586
rect 2748 8429 2749 8586
rect 2862 8011 2863 8430
rect 2751 8431 2752 8586
rect 2865 8011 2866 8432
rect 2754 8433 2755 8586
rect 2868 8011 2869 8434
rect 2769 8435 2770 8586
rect 3209 8011 3210 8436
rect 2772 8437 2773 8586
rect 2844 8011 2845 8438
rect 2775 8439 2776 8586
rect 2838 8011 2839 8440
rect 2784 8441 2785 8586
rect 2886 8011 2887 8442
rect 2796 8443 2797 8586
rect 2910 8011 2911 8444
rect 2802 8445 2803 8586
rect 3126 8011 3127 8446
rect 2808 8447 2809 8586
rect 2922 8011 2923 8448
rect 2826 8449 2827 8586
rect 2940 8011 2941 8450
rect 2829 8451 2830 8586
rect 2943 8011 2944 8452
rect 2832 8011 2833 8454
rect 3173 8011 3174 8454
rect 2832 8455 2833 8586
rect 2970 8011 2971 8456
rect 2838 8457 2839 8586
rect 2946 8011 2947 8458
rect 2856 8011 2857 8460
rect 3066 8011 3067 8460
rect 2856 8461 2857 8586
rect 2976 8011 2977 8462
rect 2862 8463 2863 8586
rect 2874 8011 2875 8464
rect 2874 8465 2875 8586
rect 3000 8011 3001 8466
rect 2883 8011 2884 8468
rect 3205 8011 3206 8468
rect 2892 8467 2893 8586
rect 2892 8011 2893 8468
rect 2895 8467 2896 8586
rect 2895 8011 2896 8468
rect 2898 8011 2899 8470
rect 3166 8011 3167 8470
rect 2898 8471 2899 8586
rect 3012 8011 3013 8472
rect 2598 8473 2599 8586
rect 3011 8473 3012 8586
rect 2901 8475 2902 8586
rect 3015 8011 3016 8476
rect 2910 8477 2911 8586
rect 3018 8011 3019 8478
rect 2916 8011 2917 8480
rect 3177 8011 3178 8480
rect 2916 8481 2917 8586
rect 3033 8011 3034 8482
rect 2712 8011 2713 8484
rect 3034 8483 3035 8586
rect 2712 8485 2713 8586
rect 2814 8011 2815 8486
rect 2814 8487 2815 8586
rect 2928 8011 2929 8488
rect 2919 8489 2920 8586
rect 2994 8011 2995 8490
rect 2928 8491 2929 8586
rect 3048 8011 3049 8492
rect 2931 8493 2932 8586
rect 2964 8011 2965 8494
rect 2934 8495 2935 8586
rect 3063 8011 3064 8496
rect 2937 8497 2938 8586
rect 2949 8497 2950 8586
rect 2940 8499 2941 8586
rect 3072 8011 3073 8500
rect 2730 8011 2731 8502
rect 3072 8501 3073 8586
rect 1644 8011 1645 8504
rect 2730 8503 2731 8586
rect 1644 8505 1645 8586
rect 1710 8011 1711 8506
rect 1680 8011 1681 8508
rect 1710 8507 1711 8586
rect 1680 8509 1681 8586
rect 2367 8011 2368 8510
rect 2355 8011 2356 8512
rect 2367 8511 2368 8586
rect 2946 8511 2947 8586
rect 3060 8011 3061 8512
rect 2952 8011 2953 8514
rect 3068 8513 3069 8586
rect 2406 8011 2407 8516
rect 2953 8515 2954 8586
rect 2388 8011 2389 8518
rect 2406 8517 2407 8586
rect 2388 8519 2389 8586
rect 2436 8011 2437 8520
rect 2436 8521 2437 8586
rect 3144 8011 3145 8522
rect 2958 8011 2959 8524
rect 3065 8523 3066 8586
rect 2959 8525 2960 8586
rect 3084 8011 3085 8526
rect 2971 8527 2972 8586
rect 3123 8011 3124 8528
rect 2986 8529 2987 8586
rect 3001 8529 3002 8586
rect 2995 8531 2996 8586
rect 3151 8011 3152 8532
rect 2998 8533 2999 8586
rect 3141 8011 3142 8534
rect 3004 8535 3005 8586
rect 3120 8011 3121 8536
rect 3006 8011 3007 8538
rect 3081 8011 3082 8538
rect 2982 8011 2983 8540
rect 3082 8539 3083 8586
rect 3009 8011 3010 8542
rect 3129 8011 3130 8542
rect 2634 8011 2635 8544
rect 3008 8543 3009 8586
rect 2634 8545 2635 8586
rect 2676 8011 2677 8546
rect 1770 8011 1771 8548
rect 2676 8547 2677 8586
rect 1770 8549 1771 8586
rect 1938 8011 1939 8550
rect 1938 8551 1939 8586
rect 1986 8011 1987 8552
rect 1986 8553 1987 8586
rect 2766 8011 2767 8554
rect 2766 8555 2767 8586
rect 2880 8011 2881 8556
rect 2880 8557 2881 8586
rect 2988 8011 2989 8558
rect 3014 8557 3015 8586
rect 3157 8011 3158 8558
rect 3017 8559 3018 8586
rect 3160 8011 3161 8560
rect 3027 8561 3028 8586
rect 3096 8011 3097 8562
rect 3030 8561 3031 8586
rect 3030 8011 3031 8562
rect 3036 8011 3037 8564
rect 3212 8011 3213 8564
rect 2983 8565 2984 8586
rect 3037 8565 3038 8586
rect 3044 8565 3045 8586
rect 3114 8011 3115 8566
rect 3047 8567 3048 8586
rect 3199 8011 3200 8568
rect 3059 8569 3060 8586
rect 3078 8011 3079 8570
rect 2688 8011 2689 8572
rect 3079 8571 3080 8586
rect 2688 8573 2689 8586
rect 2790 8011 2791 8574
rect 2790 8575 2791 8586
rect 2904 8011 2905 8576
rect 2904 8577 2905 8586
rect 3163 8011 3164 8578
rect 3062 8579 3063 8586
rect 3196 8011 3197 8580
rect 3108 8011 3109 8582
rect 3187 8011 3188 8582
rect 3138 8011 3139 8584
rect 3154 8011 3155 8584
rect 1423 8590 1424 8593
rect 2184 8590 2185 8593
rect 1423 8594 1424 9129
rect 2004 8590 2005 8595
rect 1426 8590 1427 8597
rect 1680 8590 1681 8597
rect 1426 8598 1427 9129
rect 1998 8590 1999 8599
rect 1430 8590 1431 8601
rect 2188 8600 2189 9129
rect 1430 8602 1431 9129
rect 2226 8590 2227 8603
rect 1433 8590 1434 8605
rect 2229 8590 2230 8605
rect 1437 8590 1438 8607
rect 2232 8590 2233 8607
rect 1440 8590 1441 8609
rect 1444 8590 1445 8609
rect 1444 8610 1445 9129
rect 1656 8590 1657 8611
rect 1447 8590 1448 8613
rect 1758 8590 1759 8613
rect 1433 8614 1434 9129
rect 1447 8614 1448 9129
rect 1451 8590 1452 8615
rect 1692 8590 1693 8615
rect 1451 8616 1452 9129
rect 1770 8590 1771 8617
rect 1454 8590 1455 8619
rect 1693 8618 1694 9129
rect 1454 8620 1455 9129
rect 1776 8590 1777 8621
rect 1461 8622 1462 9129
rect 2733 8590 2734 8623
rect 1466 8590 1467 8625
rect 1800 8590 1801 8625
rect 1470 8590 1471 8627
rect 2358 8590 2359 8627
rect 1470 8628 1471 9129
rect 1938 8590 1939 8629
rect 1473 8590 1474 8631
rect 1939 8630 1940 9129
rect 1473 8632 1474 9129
rect 2244 8590 2245 8633
rect 1458 8634 1459 9129
rect 2245 8634 2246 9129
rect 1494 8590 1495 8637
rect 1500 8636 1501 9129
rect 1488 8590 1489 8639
rect 1494 8638 1495 9129
rect 1512 8590 1513 8639
rect 1980 8590 1981 8639
rect 1506 8590 1507 8641
rect 1512 8640 1513 9129
rect 1506 8642 1507 9129
rect 3037 8590 3038 8643
rect 1515 8590 1516 8645
rect 1534 8644 1535 9129
rect 1518 8644 1519 9129
rect 1518 8590 1519 8645
rect 1524 8590 1525 8647
rect 1746 8590 1747 8647
rect 1531 8648 1532 9129
rect 1962 8590 1963 8649
rect 1543 8650 1544 9129
rect 1566 8590 1567 8651
rect 1552 8652 1553 9129
rect 1884 8590 1885 8653
rect 1560 8590 1561 8655
rect 1567 8654 1568 9129
rect 1554 8590 1555 8657
rect 1561 8656 1562 9129
rect 1584 8590 1585 8657
rect 1597 8656 1598 9129
rect 1588 8658 1589 9129
rect 1627 8658 1628 9129
rect 1602 8590 1603 8661
rect 1609 8660 1610 9129
rect 1620 8590 1621 8661
rect 2266 8660 2267 9129
rect 1614 8590 1615 8663
rect 1621 8662 1622 9129
rect 1644 8590 1645 8663
rect 1657 8662 1658 9129
rect 1638 8590 1639 8665
rect 1645 8664 1646 9129
rect 1674 8590 1675 8665
rect 1681 8664 1682 9129
rect 1668 8590 1669 8667
rect 1675 8666 1676 9129
rect 1662 8590 1663 8669
rect 1669 8668 1670 9129
rect 1650 8590 1651 8671
rect 1663 8670 1664 9129
rect 1585 8672 1586 9129
rect 1651 8672 1652 9129
rect 1686 8590 1687 8673
rect 1687 8672 1688 9129
rect 1722 8590 1723 8673
rect 1747 8672 1748 9129
rect 1723 8674 1724 9129
rect 1734 8590 1735 8675
rect 1716 8590 1717 8677
rect 1735 8676 1736 9129
rect 1717 8678 1718 9129
rect 1728 8590 1729 8679
rect 1729 8680 1730 9129
rect 2730 8590 2731 8681
rect 1740 8590 1741 8683
rect 1801 8682 1802 9129
rect 1741 8684 1742 9129
rect 1752 8590 1753 8685
rect 1527 8590 1528 8687
rect 1753 8686 1754 9129
rect 1527 8688 1528 9129
rect 2289 8590 2290 8689
rect 1759 8690 1760 9129
rect 1782 8590 1783 8691
rect 1764 8590 1765 8693
rect 1771 8692 1772 9129
rect 1765 8694 1766 9129
rect 1788 8590 1789 8695
rect 1463 8590 1464 8697
rect 1789 8696 1790 9129
rect 1777 8698 1778 9129
rect 1794 8590 1795 8699
rect 1783 8700 1784 9129
rect 1806 8590 1807 8701
rect 1795 8702 1796 9129
rect 1818 8590 1819 8703
rect 1807 8704 1808 9129
rect 1824 8590 1825 8705
rect 1819 8706 1820 9129
rect 1830 8590 1831 8707
rect 1825 8708 1826 9129
rect 1854 8590 1855 8709
rect 1831 8710 1832 9129
rect 1908 8590 1909 8711
rect 1848 8590 1849 8713
rect 2975 8712 2976 9129
rect 1849 8714 1850 9129
rect 1866 8590 1867 8715
rect 1855 8716 1856 9129
rect 1878 8590 1879 8717
rect 1867 8718 1868 9129
rect 1896 8590 1897 8719
rect 1872 8590 1873 8721
rect 1873 8720 1874 9129
rect 1879 8720 1880 9129
rect 1902 8590 1903 8721
rect 1894 8722 1895 9129
rect 1914 8590 1915 8723
rect 1897 8724 1898 9129
rect 2676 8590 2677 8725
rect 1903 8726 1904 9129
rect 1926 8590 1927 8727
rect 1909 8728 1910 9129
rect 1932 8590 1933 8729
rect 1915 8730 1916 9129
rect 1944 8590 1945 8731
rect 1921 8732 1922 9129
rect 1950 8590 1951 8733
rect 1927 8734 1928 9129
rect 1956 8590 1957 8735
rect 1933 8736 1934 9129
rect 1974 8590 1975 8737
rect 1945 8738 1946 9129
rect 1968 8590 1969 8739
rect 1951 8740 1952 9129
rect 2010 8590 2011 8741
rect 1957 8742 1958 9129
rect 1992 8590 1993 8743
rect 1963 8744 1964 9129
rect 2028 8590 2029 8745
rect 1969 8746 1970 9129
rect 2016 8590 2017 8747
rect 1975 8748 1976 9129
rect 2022 8590 2023 8749
rect 1981 8750 1982 9129
rect 2923 8750 2924 9129
rect 1993 8752 1994 9129
rect 2064 8590 2065 8753
rect 1572 8590 1573 8755
rect 2065 8754 2066 9129
rect 1548 8590 1549 8757
rect 1573 8756 1574 9129
rect 1549 8758 1550 9129
rect 1812 8590 1813 8759
rect 1813 8760 1814 9129
rect 1842 8590 1843 8761
rect 1843 8762 1844 9129
rect 1860 8590 1861 8763
rect 1861 8764 1862 9129
rect 1890 8590 1891 8765
rect 1999 8764 2000 9129
rect 2040 8590 2041 8765
rect 2005 8766 2006 9129
rect 2046 8590 2047 8767
rect 2011 8768 2012 9129
rect 2052 8590 2053 8769
rect 2014 8770 2015 9129
rect 2055 8590 2056 8771
rect 2017 8772 2018 9129
rect 2058 8590 2059 8773
rect 2023 8774 2024 9129
rect 2034 8590 2035 8775
rect 2029 8776 2030 9129
rect 2106 8590 2107 8777
rect 2032 8778 2033 9129
rect 2361 8590 2362 8779
rect 2035 8780 2036 9129
rect 2076 8590 2077 8781
rect 2041 8782 2042 9129
rect 2082 8590 2083 8783
rect 2047 8784 2048 9129
rect 2094 8590 2095 8785
rect 2053 8786 2054 9129
rect 2100 8590 2101 8787
rect 2059 8788 2060 9129
rect 2088 8590 2089 8789
rect 2070 8590 2071 8791
rect 2101 8790 2102 9129
rect 2071 8792 2072 9129
rect 2112 8590 2113 8793
rect 2077 8794 2078 9129
rect 2118 8590 2119 8795
rect 2083 8796 2084 9129
rect 2646 8590 2647 8797
rect 2089 8798 2090 9129
rect 2130 8590 2131 8799
rect 2095 8800 2096 9129
rect 2136 8590 2137 8801
rect 1440 8802 1441 9129
rect 2137 8802 2138 9129
rect 2107 8804 2108 9129
rect 2142 8590 2143 8805
rect 2113 8806 2114 9129
rect 2160 8590 2161 8807
rect 2119 8808 2120 9129
rect 2166 8590 2167 8809
rect 2124 8590 2125 8811
rect 2131 8810 2132 9129
rect 2125 8812 2126 9129
rect 2148 8590 2149 8813
rect 2143 8814 2144 9129
rect 2178 8590 2179 8815
rect 2149 8816 2150 9129
rect 2616 8590 2617 8817
rect 2161 8818 2162 9129
rect 2196 8590 2197 8819
rect 2167 8820 2168 9129
rect 2190 8590 2191 8821
rect 2179 8822 2180 9129
rect 2322 8590 2323 8823
rect 2185 8824 2186 9129
rect 2214 8590 2215 8825
rect 2191 8826 2192 9129
rect 2208 8590 2209 8827
rect 2197 8828 2198 9129
rect 2256 8590 2257 8829
rect 2202 8590 2203 8831
rect 3011 8590 3012 8831
rect 2203 8832 2204 9129
rect 2280 8590 2281 8833
rect 2209 8834 2210 9129
rect 2298 8590 2299 8835
rect 2215 8836 2216 9129
rect 2466 8590 2467 8837
rect 2227 8838 2228 9129
rect 2310 8590 2311 8839
rect 2233 8840 2234 9129
rect 2292 8590 2293 8841
rect 1593 8590 1594 8843
rect 2293 8842 2294 9129
rect 2250 8590 2251 8845
rect 3044 8590 3045 8845
rect 2251 8846 2252 9129
rect 2268 8590 2269 8847
rect 2254 8848 2255 9129
rect 2271 8590 2272 8849
rect 2257 8850 2258 9129
rect 2274 8590 2275 8851
rect 2260 8852 2261 9129
rect 2277 8590 2278 8853
rect 2262 8590 2263 8855
rect 2852 8854 2853 9129
rect 2263 8856 2264 9129
rect 2286 8590 2287 8857
rect 2269 8858 2270 9129
rect 2502 8590 2503 8859
rect 2275 8860 2276 9129
rect 2442 8590 2443 8861
rect 2281 8862 2282 9129
rect 2316 8590 2317 8863
rect 1575 8590 1576 8865
rect 2317 8864 2318 9129
rect 2287 8866 2288 9129
rect 2304 8590 2305 8867
rect 2299 8868 2300 9129
rect 2956 8590 2957 8869
rect 2305 8870 2306 9129
rect 2334 8590 2335 8871
rect 2308 8872 2309 9129
rect 2337 8590 2338 8873
rect 2311 8874 2312 9129
rect 2328 8590 2329 8875
rect 2314 8876 2315 9129
rect 2331 8590 2332 8877
rect 2319 8590 2320 8879
rect 2356 8878 2357 9129
rect 2323 8880 2324 9129
rect 2346 8590 2347 8881
rect 2326 8882 2327 9129
rect 2349 8590 2350 8883
rect 2329 8884 2330 9129
rect 2340 8590 2341 8885
rect 2335 8886 2336 9129
rect 2352 8590 2353 8887
rect 2341 8888 2342 9129
rect 2364 8590 2365 8889
rect 2344 8890 2345 9129
rect 2367 8590 2368 8891
rect 2347 8892 2348 9129
rect 2388 8590 2389 8893
rect 2353 8894 2354 9129
rect 2961 8894 2962 9129
rect 2359 8896 2360 9129
rect 2370 8590 2371 8897
rect 2365 8898 2366 9129
rect 2376 8590 2377 8899
rect 2371 8900 2372 9129
rect 2394 8590 2395 8901
rect 2377 8902 2378 9129
rect 2490 8590 2491 8903
rect 2389 8904 2390 9129
rect 2454 8590 2455 8905
rect 2395 8906 2396 9129
rect 2412 8590 2413 8907
rect 2400 8590 2401 8909
rect 2953 8590 2954 8909
rect 2401 8910 2402 9129
rect 2418 8590 2419 8911
rect 2413 8912 2414 9129
rect 2430 8590 2431 8913
rect 2419 8914 2420 9129
rect 2436 8590 2437 8915
rect 2431 8916 2432 9129
rect 2448 8590 2449 8917
rect 2437 8918 2438 9129
rect 2460 8590 2461 8919
rect 2443 8920 2444 9129
rect 2514 8590 2515 8921
rect 2449 8922 2450 9129
rect 2508 8590 2509 8923
rect 2455 8924 2456 9129
rect 2484 8590 2485 8925
rect 2461 8926 2462 9129
rect 2472 8590 2473 8927
rect 2467 8928 2468 9129
rect 2478 8590 2479 8929
rect 2473 8930 2474 9129
rect 2544 8590 2545 8931
rect 2479 8932 2480 9129
rect 2532 8590 2533 8933
rect 2485 8934 2486 9129
rect 2550 8590 2551 8935
rect 2491 8936 2492 9129
rect 2520 8590 2521 8937
rect 2496 8590 2497 8939
rect 3008 8590 3009 8939
rect 2497 8940 2498 9129
rect 2526 8590 2527 8941
rect 2503 8942 2504 9129
rect 2538 8590 2539 8943
rect 2509 8944 2510 9129
rect 2556 8590 2557 8945
rect 2515 8946 2516 9129
rect 2592 8590 2593 8947
rect 2521 8948 2522 9129
rect 2562 8590 2563 8949
rect 2527 8950 2528 9129
rect 2568 8590 2569 8951
rect 2533 8952 2534 9129
rect 2598 8590 2599 8953
rect 2536 8954 2537 9129
rect 2901 8590 2902 8955
rect 2539 8956 2540 9129
rect 2769 8590 2770 8957
rect 2545 8958 2546 9129
rect 2586 8590 2587 8959
rect 2551 8960 2552 9129
rect 2604 8590 2605 8961
rect 2557 8962 2558 9129
rect 2610 8590 2611 8963
rect 2563 8964 2564 9129
rect 2622 8590 2623 8965
rect 2569 8966 2570 9129
rect 2628 8590 2629 8967
rect 2574 8590 2575 8969
rect 3034 8590 3035 8969
rect 2575 8970 2576 9129
rect 2634 8590 2635 8971
rect 2581 8972 2582 9129
rect 2652 8590 2653 8973
rect 2593 8974 2594 9129
rect 2664 8590 2665 8975
rect 2605 8976 2606 9129
rect 3079 8590 3080 8977
rect 2611 8978 2612 9129
rect 2670 8590 2671 8979
rect 2617 8980 2618 9129
rect 2800 8980 2801 9129
rect 2620 8982 2621 9129
rect 2895 8590 2896 8983
rect 2623 8984 2624 9129
rect 2688 8590 2689 8985
rect 2629 8986 2630 9129
rect 2694 8590 2695 8987
rect 2635 8988 2636 9129
rect 2700 8590 2701 8989
rect 2653 8990 2654 9129
rect 2751 8590 2752 8991
rect 2656 8992 2657 9129
rect 2724 8590 2725 8993
rect 2658 8590 2659 8995
rect 3072 8590 3073 8995
rect 2659 8996 2660 9129
rect 2848 8996 2849 9129
rect 2665 8998 2666 9129
rect 2736 8590 2737 8999
rect 2671 9000 2672 9129
rect 2742 8590 2743 9001
rect 2677 9002 2678 9129
rect 2754 8590 2755 9003
rect 2695 9004 2696 9129
rect 2766 8590 2767 9005
rect 2698 9006 2699 9129
rect 3082 8590 3083 9007
rect 2701 9008 2702 9129
rect 2772 8590 2773 9009
rect 2704 9010 2705 9129
rect 2775 8590 2776 9011
rect 2719 9012 2720 9129
rect 2796 8590 2797 9013
rect 2722 9014 2723 9129
rect 2901 9014 2902 9129
rect 2725 9016 2726 9129
rect 2862 8590 2863 9017
rect 2731 9018 2732 9129
rect 2968 9018 2969 9129
rect 2737 9020 2738 9129
rect 2808 8590 2809 9021
rect 2743 9022 2744 9129
rect 2784 8590 2785 9023
rect 2761 9024 2762 9129
rect 2826 8590 2827 9025
rect 2764 9026 2765 9129
rect 2829 8590 2830 9027
rect 2767 9028 2768 9129
rect 2832 8590 2833 9029
rect 2773 9030 2774 9129
rect 2850 8590 2851 9031
rect 2785 9032 2786 9129
rect 2802 8590 2803 9033
rect 2797 9034 2798 9129
rect 2892 8590 2893 9035
rect 2818 9036 2819 9129
rect 2919 8590 2920 9037
rect 2332 9038 2333 9129
rect 2920 9038 2921 9129
rect 2821 9040 2822 9129
rect 2904 8590 2905 9041
rect 2682 8590 2683 9043
rect 2904 9042 2905 9129
rect 2683 9044 2684 9129
rect 2745 8590 2746 9045
rect 2827 9044 2828 9129
rect 2910 8590 2911 9045
rect 2833 9046 2834 9129
rect 2949 8590 2950 9047
rect 2836 9048 2837 9129
rect 2937 8590 2938 9049
rect 2790 8590 2791 9051
rect 2937 9050 2938 9129
rect 2838 8590 2839 9053
rect 3065 8590 3066 9053
rect 2839 9054 2840 9129
rect 2940 8590 2941 9055
rect 2845 9056 2846 9129
rect 3075 8590 3076 9057
rect 2856 8590 2857 9059
rect 2891 9058 2892 9129
rect 2220 8590 2221 9061
rect 2855 9060 2856 9129
rect 2221 9062 2222 9129
rect 2238 8590 2239 9063
rect 1524 9064 1525 9129
rect 2239 9064 2240 9129
rect 2858 9064 2859 9129
rect 2959 8590 2960 9065
rect 2748 8590 2749 9067
rect 2958 9066 2959 9129
rect 2749 9068 2750 9129
rect 2814 8590 2815 9069
rect 2815 9070 2816 9129
rect 3030 8590 3031 9071
rect 2870 9072 2871 9129
rect 2971 8590 2972 9073
rect 2712 8590 2713 9075
rect 2972 9074 2973 9129
rect 2880 8590 2881 9077
rect 3020 8590 3021 9077
rect 2882 9078 2883 9129
rect 3001 8590 3002 9079
rect 2885 9080 2886 9129
rect 2986 8590 2987 9081
rect 2888 9082 2889 9129
rect 2995 8590 2996 9083
rect 2894 9084 2895 9129
rect 2898 8590 2899 9085
rect 1836 8590 1837 9087
rect 2897 9086 2898 9129
rect 1437 9088 1438 9129
rect 1837 9088 1838 9129
rect 2907 9088 2908 9129
rect 3014 8590 3015 9089
rect 2910 9090 2911 9129
rect 3017 8590 3018 9091
rect 2913 9092 2914 9129
rect 3023 8590 3024 9093
rect 2916 8590 2917 9095
rect 3027 8590 3028 9095
rect 2154 8590 2155 9097
rect 2916 9096 2917 9129
rect 2155 9098 2156 9129
rect 2172 8590 2173 9099
rect 2173 9100 2174 9129
rect 2382 8590 2383 9101
rect 2383 9102 2384 9129
rect 2406 8590 2407 9103
rect 2407 9104 2408 9129
rect 2424 8590 2425 9105
rect 1590 8590 1591 9107
rect 2425 9106 2426 9129
rect 2928 8590 2929 9107
rect 3041 8590 3042 9107
rect 1986 8590 1987 9109
rect 2927 9108 2928 9129
rect 1987 9110 1988 9129
rect 2640 8590 2641 9111
rect 2641 9112 2642 9129
rect 2706 8590 2707 9113
rect 2707 9114 2708 9129
rect 2778 8590 2779 9115
rect 2931 8590 2932 9115
rect 3068 8590 3069 9115
rect 2587 9116 2588 9129
rect 2930 9116 2931 9129
rect 2934 8590 2935 9117
rect 2946 8590 2947 9117
rect 2874 8590 2875 9119
rect 2934 9118 2935 9129
rect 2940 9118 2941 9129
rect 3047 8590 3048 9119
rect 2952 9120 2953 9129
rect 3059 8590 3060 9121
rect 2955 9122 2956 9129
rect 3062 8590 3063 9123
rect 2965 9124 2966 9129
rect 2998 8590 2999 9125
rect 2983 8590 2984 9127
rect 3004 8590 3005 9127
rect 1426 9133 1427 9136
rect 1957 9133 1958 9136
rect 1426 9137 1427 9632
rect 2263 9133 2264 9138
rect 1430 9133 1431 9140
rect 1783 9133 1784 9140
rect 1430 9141 1431 9632
rect 2185 9133 2186 9142
rect 1437 9133 1438 9144
rect 2260 9133 2261 9144
rect 1440 9133 1441 9146
rect 1813 9133 1814 9146
rect 1444 9133 1445 9148
rect 2521 9133 2522 9148
rect 1444 9149 1445 9632
rect 2257 9133 2258 9150
rect 1451 9133 1452 9152
rect 2617 9133 2618 9152
rect 1458 9133 1459 9154
rect 2593 9133 2594 9154
rect 1458 9155 1459 9632
rect 2209 9133 2210 9156
rect 1461 9133 1462 9158
rect 2305 9133 2306 9158
rect 1461 9159 1462 9632
rect 1795 9133 1796 9160
rect 1470 9133 1471 9162
rect 1534 9133 1535 9162
rect 1470 9163 1471 9632
rect 2059 9133 2060 9164
rect 1473 9133 1474 9166
rect 2341 9133 2342 9166
rect 1473 9167 1474 9632
rect 2041 9133 2042 9168
rect 1494 9167 1495 9632
rect 1494 9133 1495 9168
rect 1506 9167 1507 9632
rect 1506 9133 1507 9168
rect 1512 9167 1513 9632
rect 1512 9133 1513 9168
rect 1518 9167 1519 9632
rect 1518 9133 1519 9168
rect 1531 9133 1532 9170
rect 1891 9169 1892 9632
rect 1531 9171 1532 9632
rect 2125 9133 2126 9172
rect 1534 9173 1535 9632
rect 1573 9133 1574 9174
rect 1537 9175 1538 9632
rect 1561 9133 1562 9176
rect 1543 9133 1544 9178
rect 1555 9177 1556 9632
rect 1543 9179 1544 9632
rect 1567 9133 1568 9180
rect 1549 9133 1550 9182
rect 1873 9133 1874 9182
rect 1552 9133 1553 9184
rect 1597 9133 1598 9184
rect 1564 9185 1565 9632
rect 1699 9133 1700 9186
rect 1576 9187 1577 9632
rect 2855 9133 2856 9188
rect 1585 9133 1586 9190
rect 2548 9189 2549 9632
rect 1588 9133 1589 9192
rect 2332 9133 2333 9192
rect 1603 9193 1604 9632
rect 1657 9133 1658 9194
rect 1609 9133 1610 9196
rect 1633 9195 1634 9632
rect 1609 9197 1610 9632
rect 1663 9133 1664 9198
rect 1437 9199 1438 9632
rect 1663 9199 1664 9632
rect 1615 9201 1616 9632
rect 1645 9133 1646 9202
rect 1621 9133 1622 9204
rect 1858 9203 1859 9632
rect 1621 9205 1622 9632
rect 1675 9133 1676 9206
rect 1627 9133 1628 9208
rect 2521 9207 2522 9632
rect 1627 9209 1628 9632
rect 1681 9133 1682 9210
rect 1639 9211 1640 9632
rect 1693 9133 1694 9212
rect 1645 9213 1646 9632
rect 1687 9133 1688 9214
rect 1657 9215 1658 9632
rect 1717 9133 1718 9216
rect 1675 9217 1676 9632
rect 1765 9133 1766 9218
rect 1681 9219 1682 9632
rect 1723 9133 1724 9220
rect 1687 9221 1688 9632
rect 1741 9133 1742 9222
rect 1693 9223 1694 9632
rect 1711 9133 1712 9224
rect 1423 9133 1424 9226
rect 1711 9225 1712 9632
rect 1423 9227 1424 9632
rect 2293 9133 2294 9228
rect 1717 9229 1718 9632
rect 2005 9133 2006 9230
rect 1723 9231 1724 9632
rect 2011 9133 2012 9232
rect 1726 9233 1727 9632
rect 2014 9133 2015 9234
rect 1741 9235 1742 9632
rect 1999 9133 2000 9236
rect 1747 9133 1748 9238
rect 2257 9237 2258 9632
rect 1747 9239 1748 9632
rect 2053 9133 2054 9240
rect 1765 9241 1766 9632
rect 2065 9133 2066 9242
rect 1777 9133 1778 9244
rect 2209 9243 2210 9632
rect 1777 9245 1778 9632
rect 2137 9133 2138 9246
rect 1783 9247 1784 9632
rect 1915 9133 1916 9248
rect 1795 9249 1796 9632
rect 2167 9133 2168 9250
rect 1798 9251 1799 9632
rect 2266 9133 2267 9252
rect 1813 9253 1814 9632
rect 2191 9133 2192 9254
rect 1825 9133 1826 9256
rect 2341 9255 2342 9632
rect 1825 9257 1826 9632
rect 2089 9133 2090 9258
rect 1846 9259 1847 9632
rect 2254 9133 2255 9260
rect 1852 9261 1853 9632
rect 2188 9133 2189 9262
rect 1873 9263 1874 9632
rect 2311 9133 2312 9264
rect 1885 9265 1886 9632
rect 2335 9133 2336 9266
rect 1888 9267 1889 9632
rect 2344 9133 2345 9268
rect 1894 9133 1895 9270
rect 2386 9269 2387 9632
rect 1903 9133 1904 9272
rect 2897 9133 2898 9272
rect 1524 9133 1525 9274
rect 1903 9273 1904 9632
rect 1440 9275 1441 9632
rect 1524 9275 1525 9632
rect 1915 9275 1916 9632
rect 2371 9133 2372 9276
rect 1927 9133 1928 9278
rect 2930 9133 2931 9278
rect 1927 9279 1928 9632
rect 2383 9133 2384 9280
rect 1933 9133 1934 9282
rect 2927 9133 2928 9282
rect 1933 9283 1934 9632
rect 2233 9133 2234 9284
rect 1957 9285 1958 9632
rect 2407 9133 2408 9286
rect 1999 9287 2000 9632
rect 2347 9133 2348 9288
rect 2005 9289 2006 9632
rect 2437 9133 2438 9290
rect 1735 9133 1736 9292
rect 2437 9291 2438 9632
rect 1735 9293 1736 9632
rect 2017 9133 2018 9294
rect 2011 9295 2012 9632
rect 2299 9133 2300 9296
rect 2017 9297 2018 9632
rect 2431 9133 2432 9298
rect 2023 9133 2024 9300
rect 2191 9299 2192 9632
rect 1433 9133 1434 9302
rect 2023 9301 2024 9632
rect 2032 9133 2033 9302
rect 2416 9301 2417 9632
rect 2041 9303 2042 9632
rect 2461 9133 2462 9304
rect 2053 9305 2054 9632
rect 2675 9305 2676 9632
rect 2059 9307 2060 9632
rect 2113 9133 2114 9308
rect 2029 9133 2030 9310
rect 2113 9309 2114 9632
rect 2029 9311 2030 9632
rect 2389 9133 2390 9312
rect 1849 9133 1850 9314
rect 2389 9313 2390 9632
rect 1849 9315 1850 9632
rect 2961 9133 2962 9316
rect 2065 9317 2066 9632
rect 2449 9133 2450 9318
rect 1897 9133 1898 9320
rect 2449 9319 2450 9632
rect 1897 9321 1898 9632
rect 2323 9133 2324 9322
rect 1819 9133 1820 9324
rect 2323 9323 2324 9632
rect 1819 9325 1820 9632
rect 2197 9133 2198 9326
rect 1789 9133 1790 9328
rect 2197 9327 2198 9632
rect 1789 9329 1790 9632
rect 2047 9133 2048 9330
rect 2083 9133 2084 9330
rect 2734 9329 2735 9632
rect 2083 9331 2084 9632
rect 2491 9133 2492 9332
rect 2089 9333 2090 9632
rect 2497 9133 2498 9334
rect 2098 9335 2099 9632
rect 2455 9133 2456 9336
rect 2101 9133 2102 9338
rect 2916 9133 2917 9338
rect 1969 9133 1970 9340
rect 2101 9339 2102 9632
rect 1969 9341 1970 9632
rect 2119 9133 2120 9342
rect 2119 9343 2120 9632
rect 2527 9133 2528 9344
rect 2125 9345 2126 9632
rect 2509 9133 2510 9346
rect 2131 9133 2132 9348
rect 2913 9133 2914 9348
rect 2095 9133 2096 9350
rect 2131 9349 2132 9632
rect 2095 9351 2096 9632
rect 2503 9133 2504 9352
rect 2137 9353 2138 9632
rect 2545 9133 2546 9354
rect 1651 9133 1652 9356
rect 2545 9355 2546 9632
rect 1651 9357 1652 9632
rect 1669 9133 1670 9358
rect 1669 9359 1670 9632
rect 1759 9133 1760 9360
rect 1759 9361 1760 9632
rect 2071 9133 2072 9362
rect 2071 9363 2072 9632
rect 2443 9133 2444 9364
rect 1573 9365 1574 9632
rect 2443 9365 2444 9632
rect 2143 9133 2144 9368
rect 2626 9367 2627 9632
rect 2143 9369 2144 9632
rect 2473 9133 2474 9370
rect 2149 9133 2150 9372
rect 2920 9133 2921 9372
rect 2107 9133 2108 9374
rect 2149 9373 2150 9632
rect 1939 9133 1940 9376
rect 2107 9375 2108 9632
rect 1939 9377 1940 9632
rect 2227 9133 2228 9378
rect 1945 9133 1946 9380
rect 2227 9379 2228 9632
rect 1945 9381 1946 9632
rect 2329 9133 2330 9382
rect 1951 9133 1952 9384
rect 2329 9383 2330 9632
rect 1951 9385 1952 9632
rect 2179 9133 2180 9386
rect 1993 9133 1994 9388
rect 2179 9387 2180 9632
rect 1993 9389 1994 9632
rect 2395 9133 2396 9390
rect 1843 9133 1844 9392
rect 2395 9391 2396 9632
rect 1843 9393 1844 9632
rect 2251 9133 2252 9394
rect 1771 9133 1772 9396
rect 2251 9395 2252 9632
rect 1454 9133 1455 9398
rect 1771 9397 1772 9632
rect 1454 9399 1455 9632
rect 1500 9133 1501 9400
rect 1451 9401 1452 9632
rect 1500 9401 1501 9632
rect 2161 9133 2162 9402
rect 2778 9401 2779 9632
rect 1921 9133 1922 9404
rect 2161 9403 2162 9632
rect 1921 9405 1922 9632
rect 2239 9133 2240 9406
rect 1561 9407 1562 9632
rect 2239 9407 2240 9632
rect 2164 9409 2165 9632
rect 2314 9133 2315 9410
rect 2167 9411 2168 9632
rect 2515 9133 2516 9412
rect 2173 9133 2174 9414
rect 2185 9413 2186 9632
rect 1837 9133 1838 9416
rect 2173 9415 2174 9632
rect 1837 9417 1838 9632
rect 2245 9133 2246 9418
rect 2200 9419 2201 9632
rect 2308 9133 2309 9420
rect 2212 9421 2213 9632
rect 2326 9133 2327 9422
rect 2215 9133 2216 9424
rect 2901 9133 2902 9424
rect 1855 9133 1856 9426
rect 2215 9425 2216 9632
rect 2233 9425 2234 9632
rect 2269 9133 2270 9426
rect 2155 9133 2156 9428
rect 2269 9427 2270 9632
rect 2155 9429 2156 9632
rect 2425 9133 2426 9430
rect 2245 9431 2246 9632
rect 2533 9133 2534 9432
rect 2293 9433 2294 9632
rect 2563 9133 2564 9434
rect 2299 9435 2300 9632
rect 2569 9133 2570 9436
rect 2305 9437 2306 9632
rect 2575 9133 2576 9438
rect 2311 9439 2312 9632
rect 2715 9439 2716 9632
rect 2317 9133 2318 9442
rect 2894 9133 2895 9442
rect 1801 9133 1802 9444
rect 2317 9443 2318 9632
rect 1433 9445 1434 9632
rect 1801 9445 1802 9632
rect 2335 9445 2336 9632
rect 2581 9133 2582 9446
rect 2347 9447 2348 9632
rect 2611 9133 2612 9448
rect 2356 9133 2357 9450
rect 2470 9449 2471 9632
rect 2359 9133 2360 9452
rect 2668 9451 2669 9632
rect 1831 9133 1832 9454
rect 2359 9453 2360 9632
rect 1831 9455 1832 9632
rect 2221 9133 2222 9456
rect 1753 9133 1754 9458
rect 2221 9457 2222 9632
rect 1753 9459 1754 9632
rect 2077 9133 2078 9460
rect 1527 9133 1528 9462
rect 2077 9461 2078 9632
rect 1527 9463 1528 9632
rect 2785 9133 2786 9464
rect 2371 9465 2372 9632
rect 2587 9133 2588 9466
rect 2383 9467 2384 9632
rect 2536 9133 2537 9468
rect 2407 9469 2408 9632
rect 2635 9133 2636 9470
rect 2419 9133 2420 9472
rect 2711 9471 2712 9632
rect 2419 9473 2420 9632
rect 2623 9133 2624 9474
rect 2425 9475 2426 9632
rect 2641 9133 2642 9476
rect 2431 9477 2432 9632
rect 2904 9133 2905 9478
rect 2455 9479 2456 9632
rect 2659 9133 2660 9480
rect 2461 9481 2462 9632
rect 2848 9133 2849 9482
rect 2467 9133 2468 9484
rect 2972 9133 2973 9484
rect 1705 9133 1706 9486
rect 2467 9485 2468 9632
rect 1705 9487 1706 9632
rect 1867 9133 1868 9488
rect 1867 9489 1868 9632
rect 2287 9133 2288 9490
rect 2473 9489 2474 9632
rect 2695 9133 2696 9490
rect 2476 9491 2477 9632
rect 2698 9133 2699 9492
rect 2485 9133 2486 9494
rect 2741 9493 2742 9632
rect 2485 9495 2486 9632
rect 2671 9133 2672 9496
rect 2497 9497 2498 9632
rect 2719 9133 2720 9498
rect 1963 9133 1964 9500
rect 2718 9499 2719 9632
rect 1963 9501 1964 9632
rect 2281 9133 2282 9502
rect 1981 9133 1982 9504
rect 2281 9503 2282 9632
rect 1447 9133 1448 9506
rect 1981 9505 1982 9632
rect 1447 9507 1448 9632
rect 1855 9507 1856 9632
rect 2500 9507 2501 9632
rect 2722 9133 2723 9508
rect 2515 9509 2516 9632
rect 2701 9133 2702 9510
rect 2518 9511 2519 9632
rect 2704 9133 2705 9512
rect 2527 9513 2528 9632
rect 2731 9133 2732 9514
rect 2263 9515 2264 9632
rect 2730 9515 2731 9632
rect 2533 9517 2534 9632
rect 2965 9133 2966 9518
rect 2539 9133 2540 9520
rect 2852 9133 2853 9520
rect 1729 9133 1730 9522
rect 2539 9521 2540 9632
rect 1729 9523 1730 9632
rect 1861 9133 1862 9524
rect 1861 9525 1862 9632
rect 2035 9133 2036 9526
rect 2035 9527 2036 9632
rect 2377 9133 2378 9528
rect 1909 9133 1910 9530
rect 2377 9529 2378 9632
rect 1909 9531 1910 9632
rect 2353 9133 2354 9532
rect 1879 9133 1880 9534
rect 2353 9533 2354 9632
rect 1879 9535 1880 9632
rect 2203 9133 2204 9536
rect 2551 9133 2552 9536
rect 2672 9535 2673 9632
rect 2551 9537 2552 9632
rect 2751 9537 2752 9632
rect 2557 9133 2558 9540
rect 2727 9539 2728 9632
rect 2563 9541 2564 9632
rect 2761 9133 2762 9542
rect 2566 9543 2567 9632
rect 2764 9133 2765 9544
rect 2569 9545 2570 9632
rect 2749 9133 2750 9546
rect 2575 9547 2576 9632
rect 2767 9133 2768 9548
rect 2581 9549 2582 9632
rect 2773 9133 2774 9550
rect 2593 9551 2594 9632
rect 2743 9133 2744 9552
rect 2479 9133 2480 9554
rect 2744 9553 2745 9632
rect 2479 9555 2480 9632
rect 2677 9133 2678 9556
rect 2599 9557 2600 9632
rect 2707 9133 2708 9558
rect 2401 9133 2402 9560
rect 2708 9559 2709 9632
rect 2401 9561 2402 9632
rect 2629 9133 2630 9562
rect 2605 9133 2606 9564
rect 2748 9563 2749 9632
rect 2605 9565 2606 9632
rect 2725 9133 2726 9566
rect 2611 9567 2612 9632
rect 2800 9133 2801 9568
rect 2614 9569 2615 9632
rect 2683 9133 2684 9570
rect 2620 9133 2621 9572
rect 2797 9133 2798 9572
rect 2635 9573 2636 9632
rect 2815 9133 2816 9574
rect 2638 9575 2639 9632
rect 2818 9133 2819 9576
rect 2641 9577 2642 9632
rect 2821 9133 2822 9578
rect 2647 9579 2648 9632
rect 2827 9133 2828 9580
rect 2653 9133 2654 9582
rect 2937 9133 2938 9582
rect 2653 9583 2654 9632
rect 2833 9133 2834 9584
rect 2656 9133 2657 9586
rect 2934 9133 2935 9586
rect 2656 9587 2657 9632
rect 2836 9133 2837 9588
rect 2659 9589 2660 9632
rect 2839 9133 2840 9590
rect 2665 9133 2666 9592
rect 2845 9133 2846 9592
rect 2365 9133 2366 9594
rect 2665 9593 2666 9632
rect 2678 9593 2679 9632
rect 2870 9133 2871 9594
rect 2696 9595 2697 9632
rect 2882 9133 2883 9596
rect 2699 9597 2700 9632
rect 2885 9133 2886 9598
rect 2702 9599 2703 9632
rect 2888 9133 2889 9600
rect 2705 9601 2706 9632
rect 2891 9133 2892 9602
rect 2721 9603 2722 9632
rect 2907 9133 2908 9604
rect 2724 9605 2725 9632
rect 2910 9133 2911 9606
rect 2737 9133 2738 9608
rect 2968 9133 2969 9608
rect 1987 9133 1988 9610
rect 2737 9609 2738 9632
rect 1987 9611 1988 9632
rect 2275 9133 2276 9612
rect 1807 9133 1808 9614
rect 2275 9613 2276 9632
rect 1807 9615 1808 9632
rect 1975 9133 1976 9616
rect 1975 9617 1976 9632
rect 2413 9133 2414 9618
rect 2413 9619 2414 9632
rect 2623 9619 2624 9632
rect 2754 9619 2755 9632
rect 2940 9133 2941 9620
rect 2760 9621 2761 9632
rect 2955 9133 2956 9622
rect 2772 9623 2773 9632
rect 2958 9133 2959 9624
rect 2775 9625 2776 9632
rect 2952 9133 2953 9626
rect 2781 9627 2782 9632
rect 2975 9133 2976 9628
rect 2858 9133 2859 9630
rect 2923 9133 2924 9630
rect 1423 9636 1424 9639
rect 1518 9636 1519 9639
rect 1423 9640 1424 10093
rect 1615 9636 1616 9641
rect 1426 9636 1427 9643
rect 1831 9636 1832 9643
rect 1426 9644 1427 10093
rect 2263 9636 2264 9645
rect 1430 9636 1431 9647
rect 1777 9636 1778 9647
rect 1430 9648 1431 10093
rect 2059 9636 2060 9649
rect 1433 9636 1434 9651
rect 2527 9636 2528 9651
rect 1433 9652 1434 10093
rect 2275 9636 2276 9653
rect 1437 9636 1438 9655
rect 1603 9636 1604 9655
rect 1437 9656 1438 10093
rect 1633 9636 1634 9657
rect 1440 9636 1441 9659
rect 1602 9658 1603 10093
rect 1440 9660 1441 10093
rect 2699 9636 2700 9661
rect 1444 9636 1445 9663
rect 1711 9636 1712 9663
rect 1444 9664 1445 10093
rect 2212 9636 2213 9665
rect 1447 9636 1448 9667
rect 1698 9666 1699 10093
rect 1447 9668 1448 10093
rect 1609 9636 1610 9669
rect 1451 9636 1452 9671
rect 1899 9670 1900 10093
rect 1454 9636 1455 9673
rect 2164 9636 2165 9673
rect 1456 9674 1457 10093
rect 1879 9636 1880 9675
rect 1458 9636 1459 9677
rect 1537 9636 1538 9677
rect 1459 9678 1460 10093
rect 2098 9636 2099 9679
rect 1463 9680 1464 10093
rect 1639 9636 1640 9681
rect 1466 9682 1467 10093
rect 1645 9636 1646 9683
rect 1473 9636 1474 9685
rect 1861 9636 1862 9685
rect 1481 9686 1482 10093
rect 1494 9636 1495 9687
rect 1487 9688 1488 10093
rect 1500 9636 1501 9689
rect 1493 9690 1494 10093
rect 1512 9636 1513 9691
rect 1496 9692 1497 10093
rect 1506 9636 1507 9693
rect 1499 9694 1500 10093
rect 1543 9636 1544 9695
rect 1511 9696 1512 10093
rect 2386 9636 2387 9697
rect 1518 9698 1519 10093
rect 2413 9636 2414 9699
rect 1524 9636 1525 9701
rect 2545 9636 2546 9701
rect 1527 9636 1528 9703
rect 1632 9702 1633 10093
rect 1554 9704 1555 10093
rect 1555 9636 1556 9705
rect 1566 9704 1567 10093
rect 1627 9636 1628 9705
rect 1573 9636 1574 9707
rect 2449 9636 2450 9707
rect 1572 9708 1573 10093
rect 1626 9708 1627 10093
rect 1578 9710 1579 10093
rect 1651 9636 1652 9711
rect 1590 9712 1591 10093
rect 1657 9636 1658 9713
rect 1521 9714 1522 10093
rect 1656 9714 1657 10093
rect 1596 9716 1597 10093
rect 1681 9636 1682 9717
rect 1611 9718 1612 10093
rect 2065 9636 2066 9719
rect 1614 9720 1615 10093
rect 1669 9636 1670 9721
rect 1638 9722 1639 10093
rect 1687 9636 1688 9723
rect 1644 9724 1645 10093
rect 1771 9636 1772 9725
rect 1650 9726 1651 10093
rect 2197 9636 2198 9727
rect 1663 9636 1664 9729
rect 2665 9636 2666 9729
rect 1662 9730 1663 10093
rect 1729 9636 1730 9731
rect 1668 9732 1669 10093
rect 1705 9636 1706 9733
rect 1680 9734 1681 10093
rect 1783 9636 1784 9735
rect 1686 9736 1687 10093
rect 2161 9636 2162 9737
rect 1693 9636 1694 9739
rect 2633 9738 2634 10093
rect 1692 9740 1693 10093
rect 2107 9636 2108 9741
rect 1704 9742 1705 10093
rect 1801 9636 1802 9743
rect 1710 9744 1711 10093
rect 2173 9636 2174 9745
rect 1726 9636 1727 9747
rect 1743 9746 1744 10093
rect 1728 9748 1729 10093
rect 2718 9636 2719 9749
rect 1753 9636 1754 9751
rect 1776 9750 1777 10093
rect 1747 9636 1748 9753
rect 1752 9752 1753 10093
rect 1741 9636 1742 9755
rect 1746 9754 1747 10093
rect 1723 9636 1724 9757
rect 1740 9756 1741 10093
rect 1722 9758 1723 10093
rect 1807 9636 1808 9759
rect 1759 9636 1760 9761
rect 1770 9760 1771 10093
rect 1735 9636 1736 9763
rect 1758 9762 1759 10093
rect 1717 9636 1718 9765
rect 1734 9764 1735 10093
rect 1716 9766 1717 10093
rect 2101 9636 2102 9767
rect 1764 9768 1765 10093
rect 1765 9636 1766 9769
rect 1798 9636 1799 9769
rect 1827 9768 1828 10093
rect 1800 9770 1801 10093
rect 2179 9636 2180 9771
rect 1806 9772 1807 10093
rect 2077 9636 2078 9773
rect 1830 9774 1831 10093
rect 1969 9636 1970 9775
rect 1843 9636 1844 9777
rect 1860 9776 1861 10093
rect 1819 9636 1820 9779
rect 1842 9778 1843 10093
rect 1461 9636 1462 9781
rect 1818 9780 1819 10093
rect 1846 9636 1847 9781
rect 1863 9780 1864 10093
rect 1858 9636 1859 9783
rect 1869 9782 1870 10093
rect 1867 9636 1868 9785
rect 1878 9784 1879 10093
rect 1855 9636 1856 9787
rect 1866 9786 1867 10093
rect 1837 9636 1838 9789
rect 1854 9788 1855 10093
rect 1836 9790 1837 10093
rect 2053 9636 2054 9791
rect 1888 9636 1889 9793
rect 1923 9792 1924 10093
rect 1852 9636 1853 9795
rect 1887 9794 1888 10093
rect 1851 9796 1852 10093
rect 2200 9636 2201 9797
rect 1921 9636 1922 9799
rect 2616 9798 2617 10093
rect 1885 9636 1886 9801
rect 1920 9800 1921 10093
rect 1849 9636 1850 9803
rect 1884 9802 1885 10093
rect 1813 9636 1814 9805
rect 1848 9804 1849 10093
rect 1812 9806 1813 10093
rect 1825 9636 1826 9807
rect 1795 9636 1796 9809
rect 1824 9808 1825 10093
rect 1789 9636 1790 9811
rect 1794 9810 1795 10093
rect 1470 9636 1471 9813
rect 1788 9812 1789 10093
rect 1932 9812 1933 10093
rect 1933 9636 1934 9813
rect 1968 9812 1969 10093
rect 2113 9636 2114 9813
rect 1981 9636 1982 9815
rect 2708 9636 2709 9815
rect 1980 9816 1981 10093
rect 2011 9636 2012 9817
rect 1987 9636 1988 9819
rect 2052 9818 2053 10093
rect 1957 9636 1958 9821
rect 1986 9820 1987 10093
rect 1927 9636 1928 9823
rect 1956 9822 1957 10093
rect 1903 9636 1904 9825
rect 1926 9824 1927 10093
rect 1902 9826 1903 10093
rect 2023 9636 2024 9827
rect 1993 9636 1994 9829
rect 2010 9828 2011 10093
rect 1992 9830 1993 10093
rect 2711 9636 2712 9831
rect 2005 9636 2006 9833
rect 2022 9832 2023 10093
rect 1951 9636 1952 9835
rect 2004 9834 2005 10093
rect 1915 9636 1916 9837
rect 1950 9836 1951 10093
rect 1897 9636 1898 9839
rect 1914 9838 1915 10093
rect 1873 9636 1874 9841
rect 1896 9840 1897 10093
rect 1531 9636 1532 9843
rect 1872 9842 1873 10093
rect 2029 9636 2030 9843
rect 2046 9842 2047 10093
rect 2035 9636 2036 9845
rect 2058 9844 2059 10093
rect 2041 9636 2042 9847
rect 2109 9846 2110 10093
rect 2017 9636 2018 9849
rect 2040 9848 2041 10093
rect 1999 9636 2000 9851
rect 2016 9850 2017 10093
rect 1975 9636 1976 9853
rect 1998 9852 1999 10093
rect 1963 9636 1964 9855
rect 1974 9854 1975 10093
rect 1945 9636 1946 9857
rect 1962 9856 1963 10093
rect 1939 9636 1940 9859
rect 1944 9858 1945 10093
rect 1909 9636 1910 9861
rect 1938 9860 1939 10093
rect 1891 9636 1892 9863
rect 1908 9862 1909 10093
rect 1534 9636 1535 9865
rect 1890 9864 1891 10093
rect 2071 9636 2072 9865
rect 2112 9864 2113 10093
rect 2070 9866 2071 10093
rect 2191 9636 2192 9867
rect 2073 9868 2074 10093
rect 2209 9636 2210 9869
rect 2076 9870 2077 10093
rect 2131 9636 2132 9871
rect 2083 9636 2084 9873
rect 2619 9872 2620 10093
rect 2082 9874 2083 10093
rect 2668 9636 2669 9875
rect 2095 9636 2096 9877
rect 2106 9876 2107 10093
rect 2089 9636 2090 9879
rect 2094 9878 2095 10093
rect 2088 9880 2089 10093
rect 2149 9636 2150 9881
rect 2100 9882 2101 10093
rect 2672 9636 2673 9883
rect 2125 9636 2126 9885
rect 2751 9636 2752 9885
rect 2124 9886 2125 10093
rect 2215 9636 2216 9887
rect 2130 9888 2131 10093
rect 2251 9636 2252 9889
rect 2133 9890 2134 10093
rect 2416 9636 2417 9891
rect 2142 9892 2143 10093
rect 2143 9636 2144 9893
rect 2148 9892 2149 10093
rect 2239 9636 2240 9893
rect 2155 9636 2156 9895
rect 2741 9636 2742 9895
rect 2137 9636 2138 9897
rect 2154 9896 2155 10093
rect 2119 9636 2120 9899
rect 2136 9898 2137 10093
rect 2118 9900 2119 10093
rect 2650 9900 2651 10093
rect 2160 9902 2161 10093
rect 2185 9636 2186 9903
rect 1564 9636 1565 9905
rect 2184 9904 2185 10093
rect 2167 9636 2168 9907
rect 2172 9906 2173 10093
rect 1561 9636 1562 9909
rect 2166 9908 2167 10093
rect 1560 9910 1561 10093
rect 1621 9636 1622 9911
rect 1620 9912 1621 10093
rect 1675 9636 1676 9913
rect 1608 9914 1609 10093
rect 1674 9914 1675 10093
rect 2178 9914 2179 10093
rect 2227 9636 2228 9915
rect 2190 9916 2191 10093
rect 2317 9636 2318 9917
rect 2196 9918 2197 10093
rect 2233 9636 2234 9919
rect 2202 9920 2203 10093
rect 2245 9636 2246 9921
rect 2208 9922 2209 10093
rect 2323 9636 2324 9923
rect 2214 9924 2215 10093
rect 2281 9636 2282 9925
rect 2221 9636 2222 9927
rect 2623 9636 2624 9927
rect 2034 9928 2035 10093
rect 2623 9928 2624 10093
rect 2220 9930 2221 10093
rect 2341 9636 2342 9931
rect 2226 9932 2227 10093
rect 2293 9636 2294 9933
rect 2232 9934 2233 10093
rect 2305 9636 2306 9935
rect 2238 9936 2239 10093
rect 2630 9936 2631 10093
rect 2250 9938 2251 10093
rect 2335 9636 2336 9939
rect 2257 9636 2258 9941
rect 2781 9636 2782 9941
rect 2256 9942 2257 10093
rect 2359 9636 2360 9943
rect 1514 9944 1515 10093
rect 2358 9944 2359 10093
rect 2262 9946 2263 10093
rect 2437 9636 2438 9947
rect 2269 9636 2270 9949
rect 2727 9636 2728 9949
rect 2268 9950 2269 10093
rect 2347 9636 2348 9951
rect 2274 9952 2275 10093
rect 2607 9952 2608 10093
rect 2280 9954 2281 10093
rect 2371 9636 2372 9955
rect 2286 9956 2287 10093
rect 2395 9636 2396 9957
rect 2299 9636 2300 9959
rect 2553 9958 2554 10093
rect 2298 9960 2299 10093
rect 2383 9636 2384 9961
rect 2301 9962 2302 10093
rect 2353 9636 2354 9963
rect 2304 9964 2305 10093
rect 2377 9636 2378 9965
rect 2311 9636 2312 9967
rect 2626 9636 2627 9967
rect 2310 9968 2311 10093
rect 2443 9636 2444 9969
rect 2316 9970 2317 10093
rect 2425 9636 2426 9971
rect 2322 9972 2323 10093
rect 2419 9636 2420 9973
rect 2329 9636 2330 9975
rect 2734 9636 2735 9975
rect 1576 9636 1577 9977
rect 2328 9976 2329 10093
rect 1575 9978 1576 10093
rect 2431 9636 2432 9979
rect 2334 9980 2335 10093
rect 2401 9636 2402 9981
rect 2346 9982 2347 10093
rect 2455 9636 2456 9983
rect 2352 9984 2353 10093
rect 2461 9636 2462 9985
rect 2364 9986 2365 10093
rect 2479 9636 2480 9987
rect 2370 9988 2371 10093
rect 2485 9636 2486 9989
rect 2382 9990 2383 10093
rect 2473 9636 2474 9991
rect 2385 9992 2386 10093
rect 2476 9636 2477 9993
rect 2394 9994 2395 10093
rect 2497 9636 2498 9995
rect 2397 9996 2398 10093
rect 2407 9636 2408 9997
rect 2400 9998 2401 10093
rect 2583 9998 2584 10093
rect 2412 10000 2413 10093
rect 2533 9636 2534 10001
rect 2418 10002 2419 10093
rect 2515 9636 2516 10003
rect 2421 10004 2422 10093
rect 2518 9636 2519 10005
rect 2424 10006 2425 10093
rect 2467 9636 2468 10007
rect 2427 10008 2428 10093
rect 2470 9636 2471 10009
rect 2430 10010 2431 10093
rect 2551 9636 2552 10011
rect 2028 10012 2029 10093
rect 2550 10012 2551 10093
rect 2442 10014 2443 10093
rect 2563 9636 2564 10015
rect 2445 10016 2446 10093
rect 2566 9636 2567 10017
rect 2454 10018 2455 10093
rect 2548 9636 2549 10019
rect 2457 10020 2458 10093
rect 2539 9636 2540 10021
rect 2460 10022 2461 10093
rect 2569 9636 2570 10023
rect 2466 10024 2467 10093
rect 2575 9636 2576 10025
rect 2472 10026 2473 10093
rect 2737 9636 2738 10027
rect 2478 10028 2479 10093
rect 2581 9636 2582 10029
rect 2490 10030 2491 10093
rect 2593 9636 2594 10031
rect 2496 10032 2497 10093
rect 2599 9636 2600 10033
rect 2500 9636 2501 10035
rect 2643 10034 2644 10093
rect 2502 10036 2503 10093
rect 2568 10036 2569 10093
rect 2508 10038 2509 10093
rect 2571 10038 2572 10093
rect 2526 10040 2527 10093
rect 2611 9636 2612 10041
rect 2529 10042 2530 10093
rect 2614 9636 2615 10043
rect 2532 10044 2533 10093
rect 2635 9636 2636 10045
rect 2535 10046 2536 10093
rect 2638 9636 2639 10047
rect 2544 10048 2545 10093
rect 2647 9636 2648 10049
rect 2521 9636 2522 10051
rect 2646 10050 2647 10093
rect 2556 10052 2557 10093
rect 2656 9636 2657 10053
rect 2559 10054 2560 10093
rect 2605 9636 2606 10055
rect 2389 9636 2390 10057
rect 2604 10056 2605 10093
rect 2388 10058 2389 10093
rect 2580 10058 2581 10093
rect 2574 10060 2575 10093
rect 2659 9636 2660 10061
rect 2592 10062 2593 10093
rect 2696 9636 2697 10063
rect 2595 10064 2596 10093
rect 2678 9636 2679 10065
rect 2598 10066 2599 10093
rect 2724 9636 2725 10067
rect 2601 10068 2602 10093
rect 2778 9636 2779 10069
rect 2610 10070 2611 10093
rect 2702 9636 2703 10071
rect 2613 10072 2614 10093
rect 2705 9636 2706 10073
rect 2626 10074 2627 10093
rect 2683 10074 2684 10093
rect 2637 10076 2638 10093
rect 2641 9636 2642 10077
rect 2538 10078 2539 10093
rect 2640 10078 2641 10093
rect 2653 10078 2654 10093
rect 2653 9636 2654 10079
rect 2656 10078 2657 10093
rect 2754 9636 2755 10079
rect 2662 10080 2663 10093
rect 2760 9636 2761 10081
rect 2668 10082 2669 10093
rect 2775 9636 2776 10083
rect 2675 9636 2676 10085
rect 2715 9636 2716 10085
rect 2680 10086 2681 10093
rect 2772 9636 2773 10087
rect 2721 9636 2722 10089
rect 2744 9636 2745 10089
rect 2730 9636 2731 10091
rect 2748 9636 2749 10091
rect 1423 10097 1424 10100
rect 1878 10097 1879 10100
rect 1426 10097 1427 10102
rect 1644 10097 1645 10102
rect 1430 10097 1431 10104
rect 2130 10097 2131 10104
rect 1429 10105 1430 10510
rect 1788 10097 1789 10106
rect 1433 10097 1434 10108
rect 1998 10097 1999 10108
rect 1432 10109 1433 10510
rect 1602 10097 1603 10110
rect 1437 10097 1438 10112
rect 1596 10097 1597 10112
rect 1436 10113 1437 10510
rect 1743 10097 1744 10114
rect 1440 10097 1441 10116
rect 1590 10097 1591 10116
rect 1439 10117 1440 10510
rect 1560 10097 1561 10118
rect 1447 10097 1448 10120
rect 1794 10097 1795 10120
rect 1446 10121 1447 10510
rect 1899 10097 1900 10122
rect 1459 10097 1460 10124
rect 2388 10097 2389 10124
rect 1463 10097 1464 10126
rect 2454 10097 2455 10126
rect 1462 10127 1463 10510
rect 1626 10097 1627 10128
rect 1466 10097 1467 10130
rect 2328 10097 2329 10130
rect 1465 10131 1466 10510
rect 1674 10097 1675 10132
rect 1481 10097 1482 10134
rect 2030 10133 2031 10510
rect 1480 10135 1481 10510
rect 1499 10097 1500 10136
rect 1487 10097 1488 10138
rect 2042 10137 2043 10510
rect 1486 10139 1487 10510
rect 1974 10097 1975 10140
rect 1489 10141 1490 10510
rect 1956 10097 1957 10142
rect 1493 10097 1494 10144
rect 2066 10143 2067 10510
rect 1496 10097 1497 10146
rect 1923 10097 1924 10146
rect 1498 10147 1499 10510
rect 2298 10097 2299 10148
rect 1501 10149 1502 10510
rect 2352 10097 2353 10150
rect 1505 10151 1506 10510
rect 1926 10097 1927 10152
rect 1508 10153 1509 10510
rect 2162 10153 2163 10510
rect 1511 10097 1512 10156
rect 1800 10097 1801 10156
rect 1514 10097 1515 10158
rect 2070 10097 2071 10158
rect 1518 10097 1519 10160
rect 1595 10159 1596 10510
rect 1521 10097 1522 10162
rect 1887 10097 1888 10162
rect 1523 10163 1524 10510
rect 1611 10097 1612 10164
rect 1535 10165 1536 10510
rect 1578 10097 1579 10166
rect 1541 10167 1542 10510
rect 1554 10097 1555 10168
rect 1553 10169 1554 10510
rect 2526 10097 2527 10170
rect 1556 10171 1557 10510
rect 2198 10171 2199 10510
rect 1566 10097 1567 10174
rect 1577 10173 1578 10510
rect 1568 10175 1569 10510
rect 2136 10097 2137 10176
rect 1572 10097 1573 10178
rect 2358 10097 2359 10178
rect 1458 10179 1459 10510
rect 1571 10179 1572 10510
rect 1575 10097 1576 10180
rect 2424 10097 2425 10180
rect 1583 10181 1584 10510
rect 1728 10097 1729 10182
rect 1589 10183 1590 10510
rect 2262 10097 2263 10184
rect 1601 10185 1602 10510
rect 1656 10097 1657 10186
rect 1620 10097 1621 10188
rect 1643 10187 1644 10510
rect 1619 10189 1620 10510
rect 1638 10097 1639 10190
rect 1614 10097 1615 10192
rect 1637 10191 1638 10510
rect 1613 10193 1614 10510
rect 1632 10097 1633 10194
rect 1650 10097 1651 10194
rect 1655 10193 1656 10510
rect 1649 10195 1650 10510
rect 2256 10097 2257 10196
rect 1664 10197 1665 10510
rect 2190 10097 2191 10198
rect 1673 10199 1674 10510
rect 2208 10097 2209 10200
rect 1680 10097 1681 10202
rect 2387 10201 2388 10510
rect 1679 10203 1680 10510
rect 2220 10097 2221 10204
rect 1686 10097 1687 10206
rect 1727 10205 1728 10510
rect 1722 10097 1723 10208
rect 1781 10207 1782 10510
rect 1721 10209 1722 10510
rect 2124 10097 2125 10210
rect 1734 10097 1735 10212
rect 1808 10211 1809 10510
rect 1733 10213 1734 10510
rect 2166 10097 2167 10214
rect 1787 10215 1788 10510
rect 2274 10097 2275 10216
rect 1793 10217 1794 10510
rect 2346 10097 2347 10218
rect 1827 10097 1828 10220
rect 1940 10219 1941 10510
rect 1832 10221 1833 10510
rect 2370 10097 2371 10222
rect 1836 10097 1837 10224
rect 1877 10223 1878 10510
rect 1764 10097 1765 10226
rect 1835 10225 1836 10510
rect 1698 10097 1699 10228
rect 1763 10227 1764 10510
rect 1697 10229 1698 10510
rect 2184 10097 2185 10230
rect 1848 10097 1849 10232
rect 1955 10231 1956 10510
rect 1776 10097 1777 10234
rect 1847 10233 1848 10510
rect 1716 10097 1717 10236
rect 1775 10235 1776 10510
rect 1668 10097 1669 10238
rect 1715 10237 1716 10510
rect 1851 10097 1852 10238
rect 1958 10237 1959 10510
rect 1854 10097 1855 10240
rect 1973 10239 1974 10510
rect 1853 10241 1854 10510
rect 2178 10097 2179 10242
rect 1863 10097 1864 10244
rect 1982 10243 1983 10510
rect 1869 10097 1870 10246
rect 2012 10245 2013 10510
rect 1920 10097 1921 10248
rect 2063 10247 2064 10510
rect 1925 10249 1926 10510
rect 2196 10097 2197 10250
rect 1932 10097 1933 10252
rect 2619 10097 2620 10252
rect 1931 10253 1932 10510
rect 2028 10097 2029 10254
rect 1884 10097 1885 10256
rect 2027 10255 2028 10510
rect 1883 10257 1884 10510
rect 1902 10097 1903 10258
rect 1901 10259 1902 10510
rect 2076 10097 2077 10260
rect 1938 10097 1939 10262
rect 2075 10261 2076 10510
rect 1824 10097 1825 10264
rect 1937 10263 1938 10510
rect 1752 10097 1753 10266
rect 1823 10265 1824 10510
rect 1444 10097 1445 10268
rect 1751 10267 1752 10510
rect 1443 10269 1444 10510
rect 2088 10097 2089 10270
rect 1950 10097 1951 10272
rect 2222 10271 2223 10510
rect 1872 10097 1873 10274
rect 1949 10273 1950 10510
rect 1812 10097 1813 10276
rect 1871 10275 1872 10510
rect 1746 10097 1747 10278
rect 1811 10277 1812 10510
rect 1704 10097 1705 10280
rect 1745 10279 1746 10510
rect 1703 10281 1704 10510
rect 2148 10097 2149 10282
rect 1952 10283 1953 10510
rect 2133 10097 2134 10284
rect 1997 10285 1998 10510
rect 2052 10097 2053 10286
rect 1914 10097 1915 10288
rect 2051 10287 2052 10510
rect 1818 10097 1819 10290
rect 1913 10289 1914 10510
rect 1758 10097 1759 10292
rect 1817 10291 1818 10510
rect 1757 10293 1758 10510
rect 2318 10293 2319 10510
rect 2016 10097 2017 10296
rect 2087 10295 2088 10510
rect 1908 10097 1909 10298
rect 2015 10297 2016 10510
rect 1907 10299 1908 10510
rect 2550 10097 2551 10300
rect 2024 10301 2025 10510
rect 2529 10097 2530 10302
rect 2034 10097 2035 10304
rect 2135 10303 2136 10510
rect 2033 10305 2034 10510
rect 2202 10097 2203 10306
rect 2040 10097 2041 10308
rect 2626 10097 2627 10308
rect 1896 10097 1897 10310
rect 2039 10309 2040 10510
rect 1895 10311 1896 10510
rect 2316 10097 2317 10312
rect 2046 10097 2047 10314
rect 2204 10313 2205 10510
rect 1608 10097 1609 10316
rect 2045 10315 2046 10510
rect 1565 10317 1566 10510
rect 1607 10317 1608 10510
rect 2054 10317 2055 10510
rect 2073 10097 2074 10318
rect 2058 10097 2059 10320
rect 2616 10097 2617 10320
rect 1962 10097 1963 10322
rect 2057 10321 2058 10510
rect 1842 10097 1843 10324
rect 1961 10323 1962 10510
rect 1770 10097 1771 10326
rect 1841 10325 1842 10510
rect 1769 10327 1770 10510
rect 2315 10327 2316 10510
rect 2060 10329 2061 10510
rect 2310 10097 2311 10330
rect 2069 10331 2070 10510
rect 2100 10097 2101 10332
rect 2078 10333 2079 10510
rect 2427 10097 2428 10334
rect 2082 10097 2083 10336
rect 2147 10335 2148 10510
rect 2081 10337 2082 10510
rect 2112 10097 2113 10338
rect 2010 10097 2011 10340
rect 2111 10339 2112 10510
rect 1456 10097 1457 10342
rect 2009 10341 2010 10510
rect 1455 10343 1456 10510
rect 1625 10343 1626 10510
rect 2094 10097 2095 10344
rect 2165 10343 2166 10510
rect 2093 10345 2094 10510
rect 2219 10345 2220 10510
rect 2106 10097 2107 10348
rect 2650 10097 2651 10348
rect 1992 10097 1993 10350
rect 2105 10349 2106 10510
rect 1991 10351 1992 10510
rect 2623 10097 2624 10352
rect 2118 10097 2119 10354
rect 2123 10353 2124 10510
rect 1986 10097 1987 10356
rect 2117 10355 2118 10510
rect 1866 10097 1867 10358
rect 1985 10357 1986 10510
rect 1806 10097 1807 10360
rect 1865 10359 1866 10510
rect 1740 10097 1741 10362
rect 1805 10361 1806 10510
rect 1692 10097 1693 10364
rect 1739 10363 1740 10510
rect 1691 10365 1692 10510
rect 1710 10097 1711 10366
rect 1662 10097 1663 10368
rect 1709 10367 1710 10510
rect 2129 10367 2130 10510
rect 2160 10097 2161 10368
rect 2141 10369 2142 10510
rect 2142 10097 2143 10370
rect 2154 10097 2155 10370
rect 2186 10369 2187 10510
rect 2153 10371 2154 10510
rect 2390 10371 2391 10510
rect 2159 10373 2160 10510
rect 2214 10097 2215 10374
rect 2168 10375 2169 10510
rect 2322 10097 2323 10376
rect 2172 10097 2173 10378
rect 2630 10097 2631 10378
rect 2174 10379 2175 10510
rect 2226 10097 2227 10380
rect 2180 10381 2181 10510
rect 2232 10097 2233 10382
rect 2192 10383 2193 10510
rect 2250 10097 2251 10384
rect 2201 10385 2202 10510
rect 2400 10097 2401 10386
rect 2207 10387 2208 10510
rect 2304 10097 2305 10388
rect 2225 10389 2226 10510
rect 2268 10097 2269 10390
rect 2231 10391 2232 10510
rect 2502 10097 2503 10392
rect 2238 10097 2239 10394
rect 2424 10393 2425 10510
rect 2243 10395 2244 10510
rect 2460 10097 2461 10396
rect 2249 10397 2250 10510
rect 2382 10097 2383 10398
rect 2252 10399 2253 10510
rect 2385 10097 2386 10400
rect 2255 10401 2256 10510
rect 2434 10401 2435 10510
rect 2261 10403 2262 10510
rect 2462 10403 2463 10510
rect 2267 10405 2268 10510
rect 2412 10097 2413 10406
rect 2273 10407 2274 10510
rect 2472 10097 2473 10408
rect 2286 10097 2287 10410
rect 2607 10097 2608 10410
rect 2291 10411 2292 10510
rect 2442 10097 2443 10412
rect 2294 10413 2295 10510
rect 2445 10097 2446 10414
rect 2022 10097 2023 10416
rect 2445 10415 2446 10510
rect 1980 10097 1981 10418
rect 2021 10417 2022 10510
rect 1860 10097 1861 10420
rect 1979 10419 1980 10510
rect 1859 10421 1860 10510
rect 1968 10097 1969 10422
rect 1967 10423 1968 10510
rect 2004 10097 2005 10424
rect 1944 10097 1945 10426
rect 2003 10425 2004 10510
rect 1890 10097 1891 10428
rect 1943 10427 1944 10510
rect 1830 10097 1831 10430
rect 1889 10429 1890 10510
rect 2297 10429 2298 10510
rect 2478 10097 2479 10430
rect 2301 10097 2302 10432
rect 2553 10097 2554 10432
rect 2309 10433 2310 10510
rect 2556 10097 2557 10434
rect 2312 10435 2313 10510
rect 2508 10097 2509 10436
rect 2321 10437 2322 10510
rect 2405 10437 2406 10510
rect 2334 10097 2335 10440
rect 2452 10439 2453 10510
rect 2333 10441 2334 10510
rect 2532 10097 2533 10442
rect 2336 10443 2337 10510
rect 2535 10097 2536 10444
rect 2339 10445 2340 10510
rect 2640 10097 2641 10446
rect 2345 10447 2346 10510
rect 2408 10447 2409 10510
rect 2351 10449 2352 10510
rect 2438 10449 2439 10510
rect 2357 10451 2358 10510
rect 2441 10451 2442 10510
rect 2364 10097 2365 10454
rect 2643 10097 2644 10454
rect 2369 10455 2370 10510
rect 2574 10097 2575 10456
rect 2375 10457 2376 10510
rect 2633 10097 2634 10458
rect 2381 10459 2382 10510
rect 2598 10097 2599 10460
rect 2384 10461 2385 10510
rect 2601 10097 2602 10462
rect 2394 10097 2395 10464
rect 2646 10097 2647 10464
rect 2397 10097 2398 10466
rect 2455 10465 2456 10510
rect 2399 10467 2400 10510
rect 2592 10097 2593 10468
rect 2402 10469 2403 10510
rect 2595 10097 2596 10470
rect 2411 10471 2412 10510
rect 2610 10097 2611 10472
rect 2414 10473 2415 10510
rect 2613 10097 2614 10474
rect 2418 10097 2419 10476
rect 2583 10097 2584 10476
rect 2109 10097 2110 10478
rect 2417 10477 2418 10510
rect 2421 10097 2422 10478
rect 2580 10097 2581 10478
rect 2280 10097 2281 10480
rect 2420 10479 2421 10510
rect 2279 10481 2280 10510
rect 2430 10097 2431 10482
rect 2427 10483 2428 10510
rect 2538 10097 2539 10484
rect 2431 10485 2432 10510
rect 2466 10097 2467 10486
rect 2448 10487 2449 10510
rect 2604 10097 2605 10488
rect 2457 10097 2458 10490
rect 2568 10097 2569 10490
rect 2459 10491 2460 10510
rect 2496 10097 2497 10492
rect 2465 10493 2466 10510
rect 2656 10097 2657 10494
rect 2471 10495 2472 10510
rect 2662 10097 2663 10496
rect 2477 10497 2478 10510
rect 2668 10097 2669 10498
rect 2490 10097 2491 10500
rect 2653 10097 2654 10500
rect 2489 10501 2490 10510
rect 2680 10097 2681 10502
rect 2492 10503 2493 10510
rect 2683 10097 2684 10504
rect 2544 10097 2545 10506
rect 2637 10097 2638 10506
rect 2559 10097 2560 10508
rect 2571 10097 2572 10508
rect 1429 10514 1430 10517
rect 1535 10514 1536 10517
rect 1432 10514 1433 10519
rect 2027 10514 2028 10519
rect 1436 10514 1437 10521
rect 1769 10514 1770 10521
rect 1439 10514 1440 10523
rect 1664 10514 1665 10523
rect 1441 10524 1442 10851
rect 1649 10514 1650 10525
rect 1443 10514 1444 10527
rect 2009 10514 2010 10527
rect 1444 10528 1445 10851
rect 1480 10514 1481 10529
rect 1448 10530 1449 10851
rect 1733 10514 1734 10531
rect 1451 10532 1452 10851
rect 1781 10514 1782 10533
rect 1455 10514 1456 10535
rect 1619 10514 1620 10535
rect 1455 10536 1456 10851
rect 1745 10514 1746 10537
rect 1458 10514 1459 10539
rect 1613 10514 1614 10539
rect 1465 10514 1466 10541
rect 1691 10514 1692 10541
rect 1467 10542 1468 10851
rect 1534 10542 1535 10851
rect 1470 10544 1471 10851
rect 2030 10514 2031 10545
rect 1479 10546 1480 10851
rect 1883 10514 1884 10547
rect 1482 10548 1483 10851
rect 1819 10548 1820 10851
rect 1486 10514 1487 10551
rect 2411 10514 2412 10551
rect 1486 10552 1487 10851
rect 1958 10514 1959 10553
rect 1489 10514 1490 10555
rect 1889 10514 1890 10555
rect 1489 10556 1490 10851
rect 1565 10514 1566 10557
rect 1498 10514 1499 10559
rect 2015 10514 2016 10559
rect 1498 10560 1499 10851
rect 1952 10514 1953 10561
rect 1505 10514 1506 10563
rect 1985 10514 1986 10563
rect 1504 10564 1505 10851
rect 1541 10514 1542 10565
rect 1510 10566 1511 10851
rect 1633 10566 1634 10851
rect 1523 10514 1524 10569
rect 1528 10568 1529 10851
rect 1462 10514 1463 10571
rect 1522 10570 1523 10851
rect 1537 10570 1538 10851
rect 1963 10570 1964 10851
rect 1553 10514 1554 10573
rect 1901 10514 1902 10573
rect 1552 10574 1553 10851
rect 2434 10514 2435 10575
rect 1556 10514 1557 10577
rect 2180 10514 2181 10577
rect 1558 10578 1559 10851
rect 2045 10514 2046 10579
rect 1561 10580 1562 10851
rect 1757 10514 1758 10581
rect 1568 10514 1569 10583
rect 2345 10514 2346 10583
rect 1577 10514 1578 10585
rect 1777 10584 1778 10851
rect 1576 10586 1577 10851
rect 1832 10514 1833 10587
rect 1612 10588 1613 10851
rect 1637 10514 1638 10589
rect 1618 10590 1619 10851
rect 1643 10514 1644 10591
rect 1630 10592 1631 10851
rect 2021 10514 2022 10593
rect 1651 10594 1652 10851
rect 1673 10514 1674 10595
rect 1655 10514 1656 10597
rect 2219 10514 2220 10597
rect 1654 10598 1655 10851
rect 2231 10514 2232 10599
rect 1660 10600 1661 10851
rect 1793 10514 1794 10601
rect 1666 10602 1667 10851
rect 2315 10514 2316 10603
rect 1672 10604 1673 10851
rect 1709 10514 1710 10605
rect 1684 10606 1685 10851
rect 1703 10514 1704 10607
rect 1446 10514 1447 10609
rect 1702 10608 1703 10851
rect 1690 10610 1691 10851
rect 1751 10514 1752 10611
rect 1708 10612 1709 10851
rect 1763 10514 1764 10613
rect 1720 10614 1721 10851
rect 1721 10514 1722 10615
rect 1727 10514 1728 10615
rect 2390 10514 2391 10615
rect 1697 10514 1698 10617
rect 1726 10616 1727 10851
rect 1732 10616 1733 10851
rect 1775 10514 1776 10617
rect 1735 10618 1736 10851
rect 2042 10514 2043 10619
rect 1750 10620 1751 10851
rect 1805 10514 1806 10621
rect 1753 10622 1754 10851
rect 1808 10514 1809 10623
rect 1756 10624 1757 10851
rect 1811 10514 1812 10625
rect 1762 10626 1763 10851
rect 1817 10514 1818 10627
rect 1774 10628 1775 10851
rect 1823 10514 1824 10629
rect 1780 10630 1781 10851
rect 2201 10514 2202 10631
rect 1789 10632 1790 10851
rect 1841 10514 1842 10633
rect 1795 10634 1796 10851
rect 1847 10514 1848 10635
rect 1801 10636 1802 10851
rect 1853 10514 1854 10637
rect 1807 10638 1808 10851
rect 1865 10514 1866 10639
rect 1813 10640 1814 10851
rect 1877 10514 1878 10641
rect 1831 10642 1832 10851
rect 2168 10514 2169 10643
rect 1835 10514 1836 10645
rect 1888 10644 1889 10851
rect 1843 10646 1844 10851
rect 1925 10514 1926 10647
rect 1849 10648 1850 10851
rect 1937 10514 1938 10649
rect 1852 10650 1853 10851
rect 1940 10514 1941 10651
rect 1855 10652 1856 10851
rect 1913 10514 1914 10653
rect 1859 10514 1860 10655
rect 2176 10654 2177 10851
rect 1861 10656 1862 10851
rect 1991 10514 1992 10657
rect 1867 10658 1868 10851
rect 2033 10514 2034 10659
rect 1871 10514 1872 10661
rect 2101 10660 2102 10851
rect 1873 10662 1874 10851
rect 1961 10514 1962 10663
rect 1876 10664 1877 10851
rect 2012 10514 2013 10665
rect 1879 10666 1880 10851
rect 1973 10514 1974 10667
rect 1885 10668 1886 10851
rect 1979 10514 1980 10669
rect 1891 10670 1892 10851
rect 1955 10514 1956 10671
rect 1895 10514 1896 10673
rect 2131 10672 2132 10851
rect 1739 10514 1740 10675
rect 1894 10674 1895 10851
rect 1738 10676 1739 10851
rect 1787 10514 1788 10677
rect 1897 10676 1898 10851
rect 2159 10514 2160 10677
rect 1903 10678 1904 10851
rect 1943 10514 1944 10679
rect 1907 10514 1908 10681
rect 2424 10514 2425 10681
rect 1458 10682 1459 10851
rect 1906 10682 1907 10851
rect 1909 10682 1910 10851
rect 2003 10514 2004 10683
rect 1915 10684 1916 10851
rect 1931 10514 1932 10685
rect 1921 10686 1922 10851
rect 1967 10514 1968 10687
rect 1924 10688 1925 10851
rect 2024 10514 2025 10689
rect 1927 10690 1928 10851
rect 2051 10514 2052 10691
rect 1930 10692 1931 10851
rect 2054 10514 2055 10693
rect 1936 10694 1937 10851
rect 2312 10514 2313 10695
rect 1939 10696 1940 10851
rect 2063 10514 2064 10697
rect 1942 10698 1943 10851
rect 2066 10514 2067 10699
rect 1945 10700 1946 10851
rect 2057 10514 2058 10701
rect 1501 10514 1502 10703
rect 2056 10702 2057 10851
rect 1949 10514 1950 10705
rect 2196 10704 2197 10851
rect 1679 10514 1680 10707
rect 1948 10706 1949 10851
rect 1678 10708 1679 10851
rect 1715 10514 1716 10709
rect 1508 10514 1509 10711
rect 1714 10710 1715 10851
rect 1951 10710 1952 10851
rect 2075 10514 2076 10711
rect 1954 10712 1955 10851
rect 2078 10514 2079 10713
rect 1957 10714 1958 10851
rect 2179 10714 2180 10851
rect 1969 10716 1970 10851
rect 2093 10514 2094 10717
rect 1972 10718 1973 10851
rect 2309 10514 2310 10719
rect 1975 10720 1976 10851
rect 2081 10514 2082 10721
rect 1982 10514 1983 10723
rect 2455 10514 2456 10723
rect 1981 10724 1982 10851
rect 2123 10514 2124 10725
rect 1987 10726 1988 10851
rect 2069 10514 2070 10727
rect 1993 10728 1994 10851
rect 2117 10514 2118 10729
rect 1997 10514 1998 10731
rect 2098 10730 2099 10851
rect 1999 10732 2000 10851
rect 2111 10514 2112 10733
rect 2002 10734 2003 10851
rect 2162 10514 2163 10735
rect 2005 10736 2006 10851
rect 2427 10514 2428 10737
rect 2011 10738 2012 10851
rect 2135 10514 2136 10739
rect 2017 10740 2018 10851
rect 2147 10514 2148 10741
rect 2029 10742 2030 10851
rect 2141 10514 2142 10743
rect 2039 10514 2040 10745
rect 2140 10744 2141 10851
rect 2041 10746 2042 10851
rect 2192 10514 2193 10747
rect 2047 10748 2048 10851
rect 2198 10514 2199 10749
rect 2060 10514 2061 10751
rect 2420 10514 2421 10751
rect 2062 10752 2063 10851
rect 2207 10514 2208 10753
rect 2068 10754 2069 10851
rect 2252 10514 2253 10755
rect 2071 10756 2072 10851
rect 2186 10514 2187 10757
rect 1601 10514 1602 10759
rect 2186 10758 2187 10851
rect 1600 10760 1601 10851
rect 1625 10514 1626 10761
rect 1607 10514 1608 10763
rect 1624 10762 1625 10851
rect 1595 10514 1596 10765
rect 1606 10764 1607 10851
rect 1589 10514 1590 10767
rect 1594 10766 1595 10851
rect 1583 10514 1584 10769
rect 1588 10768 1589 10851
rect 1571 10514 1572 10771
rect 1582 10770 1583 10851
rect 2074 10770 2075 10851
rect 2273 10514 2274 10771
rect 2080 10772 2081 10851
rect 2452 10514 2453 10773
rect 2083 10774 2084 10851
rect 2165 10514 2166 10775
rect 2087 10514 2088 10777
rect 2448 10514 2449 10777
rect 2086 10778 2087 10851
rect 2243 10514 2244 10779
rect 2092 10780 2093 10851
rect 2414 10514 2415 10781
rect 2095 10782 2096 10851
rect 2297 10514 2298 10783
rect 2105 10514 2106 10785
rect 2143 10784 2144 10851
rect 2110 10786 2111 10851
rect 2279 10514 2280 10787
rect 2122 10788 2123 10851
rect 2291 10514 2292 10789
rect 2125 10790 2126 10851
rect 2294 10514 2295 10791
rect 2129 10514 2130 10793
rect 2202 10792 2203 10851
rect 2128 10794 2129 10851
rect 2333 10514 2334 10795
rect 2134 10796 2135 10851
rect 2339 10514 2340 10797
rect 2146 10798 2147 10851
rect 2351 10514 2352 10799
rect 2153 10514 2154 10801
rect 2190 10800 2191 10851
rect 2158 10802 2159 10851
rect 2399 10514 2400 10803
rect 2161 10804 2162 10851
rect 2321 10514 2322 10805
rect 2164 10806 2165 10851
rect 2336 10514 2337 10807
rect 2167 10808 2168 10851
rect 2193 10808 2194 10851
rect 2170 10810 2171 10851
rect 2381 10514 2382 10811
rect 2174 10514 2175 10813
rect 2199 10812 2200 10851
rect 2173 10814 2174 10851
rect 2357 10514 2358 10815
rect 2183 10816 2184 10851
rect 2402 10514 2403 10817
rect 2204 10514 2205 10819
rect 2387 10514 2388 10819
rect 2205 10820 2206 10851
rect 2438 10514 2439 10821
rect 2208 10822 2209 10851
rect 2465 10514 2466 10823
rect 2220 10824 2221 10851
rect 2489 10514 2490 10825
rect 2222 10514 2223 10827
rect 2249 10514 2250 10827
rect 2223 10828 2224 10851
rect 2492 10514 2493 10829
rect 2225 10514 2226 10831
rect 2462 10514 2463 10831
rect 2226 10832 2227 10851
rect 2471 10514 2472 10833
rect 2229 10834 2230 10851
rect 2477 10514 2478 10835
rect 2255 10514 2256 10837
rect 2417 10514 2418 10837
rect 2261 10514 2262 10839
rect 2431 10514 2432 10839
rect 2267 10514 2268 10841
rect 2459 10514 2460 10841
rect 2318 10514 2319 10843
rect 2445 10514 2446 10843
rect 2369 10514 2370 10845
rect 2405 10514 2406 10845
rect 2375 10514 2376 10847
rect 2408 10514 2409 10847
rect 2384 10514 2385 10849
rect 2441 10514 2442 10849
rect 1423 10857 1424 11106
rect 1714 10855 1715 10858
rect 1426 10859 1427 11106
rect 1600 10855 1601 10860
rect 1430 10861 1431 11106
rect 1873 10855 1874 10862
rect 1433 10863 1434 11106
rect 1921 10855 1922 10864
rect 1437 10865 1438 11106
rect 1795 10855 1796 10866
rect 1441 10855 1442 10868
rect 1606 10855 1607 10868
rect 1440 10869 1441 11106
rect 1753 10855 1754 10870
rect 1444 10855 1445 10872
rect 1682 10871 1683 11106
rect 1444 10873 1445 11106
rect 1528 10855 1529 10874
rect 1451 10855 1452 10876
rect 1732 10855 1733 10876
rect 1450 10877 1451 11106
rect 1903 10855 1904 10878
rect 1453 10879 1454 11106
rect 2029 10855 2030 10880
rect 1458 10855 1459 10882
rect 1894 10855 1895 10882
rect 1448 10855 1449 10884
rect 1459 10883 1460 11106
rect 1447 10885 1448 11106
rect 1522 10855 1523 10886
rect 1462 10887 1463 11106
rect 1684 10855 1685 10888
rect 1467 10855 1468 10890
rect 1651 10855 1652 10890
rect 1470 10855 1471 10892
rect 1948 10855 1949 10892
rect 1477 10893 1478 11106
rect 2101 10855 2102 10894
rect 1479 10855 1480 10896
rect 1813 10855 1814 10896
rect 1482 10855 1483 10898
rect 1807 10855 1808 10898
rect 1486 10855 1487 10900
rect 1720 10855 1721 10900
rect 1489 10855 1490 10902
rect 1777 10855 1778 10902
rect 1489 10903 1490 11106
rect 1927 10855 1928 10904
rect 1496 10905 1497 11106
rect 1510 10855 1511 10906
rect 1498 10855 1499 10908
rect 1508 10907 1509 11106
rect 1499 10909 1500 11106
rect 1504 10855 1505 10910
rect 1511 10909 1512 11106
rect 1906 10855 1907 10910
rect 1514 10911 1515 11106
rect 1552 10855 1553 10912
rect 1520 10913 1521 11106
rect 1588 10855 1589 10914
rect 1526 10915 1527 11106
rect 1594 10855 1595 10916
rect 1532 10917 1533 11106
rect 1612 10855 1613 10918
rect 1537 10855 1538 10920
rect 1951 10855 1952 10920
rect 1538 10921 1539 11106
rect 1618 10855 1619 10922
rect 1544 10923 1545 11106
rect 1624 10855 1625 10924
rect 1550 10925 1551 11106
rect 1582 10855 1583 10926
rect 1558 10855 1559 10928
rect 1924 10855 1925 10928
rect 1561 10855 1562 10930
rect 1766 10929 1767 11106
rect 1568 10931 1569 11106
rect 1660 10855 1661 10932
rect 1586 10933 1587 11106
rect 1672 10855 1673 10934
rect 1592 10935 1593 11106
rect 1678 10855 1679 10936
rect 1595 10937 1596 11106
rect 1876 10855 1877 10938
rect 1598 10939 1599 11106
rect 1708 10855 1709 10940
rect 1604 10941 1605 11106
rect 1865 10941 1866 11106
rect 1622 10943 1623 11106
rect 1750 10855 1751 10944
rect 1625 10945 1626 11106
rect 1756 10855 1757 10946
rect 1630 10855 1631 10948
rect 2161 10855 2162 10948
rect 1631 10949 1632 11106
rect 1762 10855 1763 10950
rect 1576 10855 1577 10952
rect 1763 10951 1764 11106
rect 1577 10953 1578 11106
rect 1954 10855 1955 10954
rect 1633 10855 1634 10956
rect 2041 10855 2042 10956
rect 1534 10855 1535 10958
rect 1634 10957 1635 11106
rect 1637 10957 1638 11106
rect 1690 10855 1691 10958
rect 1643 10959 1644 11106
rect 1702 10855 1703 10960
rect 1661 10961 1662 11106
rect 1738 10855 1739 10962
rect 1673 10963 1674 11106
rect 1780 10855 1781 10964
rect 1455 10855 1456 10966
rect 1781 10965 1782 11106
rect 1456 10967 1457 11106
rect 1735 10855 1736 10968
rect 1676 10969 1677 11106
rect 2143 10855 2144 10970
rect 1688 10971 1689 11106
rect 1831 10855 1832 10972
rect 1694 10973 1695 11106
rect 1849 10855 1850 10974
rect 1697 10975 1698 11106
rect 1852 10855 1853 10976
rect 1712 10977 1713 11106
rect 1891 10855 1892 10978
rect 1715 10979 1716 11106
rect 1855 10855 1856 10980
rect 1724 10981 1725 11106
rect 1879 10855 1880 10982
rect 1726 10855 1727 10984
rect 1950 10983 1951 11106
rect 1730 10985 1731 11106
rect 1885 10855 1886 10986
rect 1733 10987 1734 11106
rect 1888 10855 1889 10988
rect 1736 10989 1737 11106
rect 1897 10855 1898 10990
rect 1742 10991 1743 11106
rect 1843 10855 1844 10992
rect 1748 10993 1749 11106
rect 1909 10855 1910 10994
rect 1654 10855 1655 10996
rect 1910 10995 1911 11106
rect 1655 10997 1656 11106
rect 1789 10855 1790 10998
rect 1754 10999 1755 11106
rect 1867 10855 1868 11000
rect 1760 11001 1761 11106
rect 1915 10855 1916 11002
rect 1769 11003 1770 11106
rect 1939 10855 1940 11004
rect 1666 10855 1667 11006
rect 1939 11005 1940 11106
rect 1772 11007 1773 11106
rect 1942 10855 1943 11008
rect 1774 10855 1775 11010
rect 2179 10855 2180 11010
rect 1492 11011 1493 11106
rect 1775 11011 1776 11106
rect 1778 11011 1779 11106
rect 1930 10855 1931 11012
rect 1787 11013 1788 11106
rect 1920 11013 1921 11106
rect 1790 11015 1791 11106
rect 2002 10855 2003 11016
rect 1793 11017 1794 11106
rect 1963 10855 1964 11018
rect 1799 11019 1800 11106
rect 1969 10855 1970 11020
rect 1801 10855 1802 11022
rect 1953 11021 1954 11106
rect 1805 11023 1806 11106
rect 2183 10855 2184 11024
rect 1811 11025 1812 11106
rect 1975 10855 1976 11026
rect 1817 11027 1818 11106
rect 1981 10855 1982 11028
rect 1819 10855 1820 11030
rect 2140 10855 2141 11030
rect 1823 11031 1824 11106
rect 1987 10855 1988 11032
rect 1829 11033 1830 11106
rect 2011 10855 2012 11034
rect 1835 11035 1836 11106
rect 2005 10855 2006 11036
rect 1841 11037 1842 11106
rect 2199 10855 2200 11038
rect 1847 11039 1848 11106
rect 2056 10855 2057 11040
rect 1859 11041 1860 11106
rect 2047 10855 2048 11042
rect 1861 10855 1862 11044
rect 1913 11043 1914 11106
rect 1574 11045 1575 11106
rect 1862 11045 1863 11106
rect 1868 11045 1869 11106
rect 2071 10855 2072 11046
rect 1877 11047 1878 11106
rect 2092 10855 2093 11048
rect 1880 11049 1881 11106
rect 2095 10855 2096 11050
rect 1883 11051 1884 11106
rect 1972 10855 1973 11052
rect 1886 11053 1887 11106
rect 1936 10855 1937 11054
rect 1889 11055 1890 11106
rect 2128 10855 2129 11056
rect 1892 11057 1893 11106
rect 2131 10855 2132 11058
rect 1895 11059 1896 11106
rect 2122 10855 2123 11060
rect 1904 11061 1905 11106
rect 2158 10855 2159 11062
rect 1907 11063 1908 11106
rect 2167 10855 2168 11064
rect 1917 11065 1918 11106
rect 1957 10855 1958 11066
rect 1923 11067 1924 11106
rect 2170 10855 2171 11068
rect 1926 11069 1927 11106
rect 2146 10855 2147 11070
rect 1929 11071 1930 11106
rect 2086 10855 2087 11072
rect 1932 11073 1933 11106
rect 2074 10855 2075 11074
rect 1936 11075 1937 11106
rect 1945 10855 1946 11076
rect 1853 11077 1854 11106
rect 1946 11077 1947 11106
rect 1943 11079 1944 11106
rect 2062 10855 2063 11080
rect 1956 11081 1957 11106
rect 2110 10855 2111 11082
rect 1959 11083 1960 11106
rect 2125 10855 2126 11084
rect 1993 10855 1994 11086
rect 2176 10855 2177 11086
rect 1999 10855 2000 11088
rect 2186 10855 2187 11088
rect 2017 10855 2018 11090
rect 2193 10855 2194 11090
rect 2068 10855 2069 11092
rect 2098 10855 2099 11092
rect 2080 10855 2081 11094
rect 2205 10855 2206 11094
rect 2083 10855 2084 11096
rect 2196 10855 2197 11096
rect 2134 10855 2135 11098
rect 2202 10855 2203 11098
rect 2164 10855 2165 11100
rect 2208 10855 2209 11100
rect 2173 10855 2174 11102
rect 2190 10855 2191 11102
rect 2220 10855 2221 11102
rect 2229 10855 2230 11102
rect 2223 10855 2224 11104
rect 2226 10855 2227 11104
rect 1423 11110 1424 11113
rect 1604 11110 1605 11113
rect 1426 11110 1427 11115
rect 1598 11110 1599 11115
rect 1430 11110 1431 11117
rect 1534 11116 1535 11265
rect 1429 11118 1430 11265
rect 1631 11110 1632 11119
rect 1433 11110 1434 11121
rect 1748 11110 1749 11121
rect 1432 11122 1433 11265
rect 1763 11110 1764 11123
rect 1437 11110 1438 11125
rect 1655 11110 1656 11125
rect 1436 11126 1437 11265
rect 1772 11110 1773 11127
rect 1440 11110 1441 11129
rect 1733 11110 1734 11129
rect 1439 11130 1440 11265
rect 1538 11110 1539 11131
rect 1444 11110 1445 11133
rect 1477 11110 1478 11133
rect 1443 11134 1444 11265
rect 1532 11110 1533 11135
rect 1447 11110 1448 11137
rect 1595 11110 1596 11137
rect 1446 11138 1447 11265
rect 1592 11110 1593 11139
rect 1450 11110 1451 11141
rect 1622 11110 1623 11141
rect 1450 11142 1451 11265
rect 1715 11110 1716 11143
rect 1453 11110 1454 11145
rect 1712 11110 1713 11145
rect 1453 11146 1454 11265
rect 1787 11110 1788 11147
rect 1456 11146 1457 11265
rect 1456 11110 1457 11147
rect 1459 11110 1460 11149
rect 1643 11110 1644 11149
rect 1462 11110 1463 11151
rect 1637 11110 1638 11151
rect 1465 11152 1466 11265
rect 1694 11110 1695 11153
rect 1468 11154 1469 11265
rect 1625 11110 1626 11155
rect 1471 11156 1472 11265
rect 1634 11110 1635 11157
rect 1474 11158 1475 11265
rect 1586 11110 1587 11159
rect 1483 11160 1484 11265
rect 1730 11110 1731 11161
rect 1486 11162 1487 11265
rect 1724 11110 1725 11163
rect 1489 11110 1490 11165
rect 1883 11110 1884 11165
rect 1489 11166 1490 11265
rect 1697 11110 1698 11167
rect 1492 11110 1493 11169
rect 1835 11110 1836 11169
rect 1492 11170 1493 11265
rect 1917 11110 1918 11171
rect 1496 11110 1497 11173
rect 1508 11110 1509 11173
rect 1495 11174 1496 11265
rect 1778 11110 1779 11175
rect 1499 11110 1500 11177
rect 1511 11110 1512 11177
rect 1498 11178 1499 11265
rect 1769 11110 1770 11179
rect 1501 11180 1502 11265
rect 1544 11110 1545 11181
rect 1504 11182 1505 11265
rect 1526 11110 1527 11183
rect 1507 11184 1508 11265
rect 1520 11110 1521 11185
rect 1514 11110 1515 11187
rect 1519 11186 1520 11265
rect 1513 11188 1514 11265
rect 1550 11110 1551 11189
rect 1525 11190 1526 11265
rect 1760 11110 1761 11191
rect 1546 11192 1547 11265
rect 1907 11110 1908 11193
rect 1555 11194 1556 11265
rect 1829 11110 1830 11195
rect 1561 11196 1562 11265
rect 1754 11110 1755 11197
rect 1564 11198 1565 11265
rect 1790 11110 1791 11199
rect 1568 11110 1569 11201
rect 1603 11200 1604 11265
rect 1574 11110 1575 11203
rect 1585 11202 1586 11265
rect 1573 11204 1574 11265
rect 1823 11110 1824 11205
rect 1577 11110 1578 11207
rect 1588 11206 1589 11265
rect 1576 11208 1577 11265
rect 1793 11110 1794 11209
rect 1579 11210 1580 11265
rect 1886 11110 1887 11211
rect 1582 11212 1583 11265
rect 1799 11110 1800 11213
rect 1597 11214 1598 11265
rect 1892 11110 1893 11215
rect 1600 11216 1601 11265
rect 1676 11110 1677 11217
rect 1606 11218 1607 11265
rect 1805 11110 1806 11219
rect 1609 11220 1610 11265
rect 1736 11110 1737 11221
rect 1612 11222 1613 11265
rect 1661 11110 1662 11223
rect 1616 11224 1617 11265
rect 1817 11110 1818 11225
rect 1619 11226 1620 11265
rect 1811 11110 1812 11227
rect 1623 11228 1624 11265
rect 1688 11110 1689 11229
rect 1626 11230 1627 11265
rect 1682 11110 1683 11231
rect 1629 11232 1630 11265
rect 1775 11110 1776 11233
rect 1632 11234 1633 11265
rect 1868 11110 1869 11235
rect 1673 11110 1674 11237
rect 1953 11110 1954 11237
rect 1742 11110 1743 11239
rect 1913 11110 1914 11239
rect 1766 11110 1767 11241
rect 1865 11110 1866 11241
rect 1781 11110 1782 11243
rect 1946 11110 1947 11243
rect 1841 11110 1842 11245
rect 1939 11110 1940 11245
rect 1847 11110 1848 11247
rect 1943 11110 1944 11247
rect 1853 11110 1854 11249
rect 1862 11110 1863 11249
rect 1859 11110 1860 11251
rect 1950 11110 1951 11251
rect 1877 11110 1878 11253
rect 1932 11110 1933 11253
rect 1880 11110 1881 11255
rect 1929 11110 1930 11255
rect 1889 11110 1890 11257
rect 1910 11110 1911 11257
rect 1895 11110 1896 11259
rect 1956 11110 1957 11259
rect 1904 11110 1905 11261
rect 1920 11110 1921 11261
rect 1923 11110 1924 11261
rect 1959 11110 1960 11261
rect 1926 11110 1927 11263
rect 1936 11110 1937 11263
rect 1429 11269 1430 11272
rect 1468 11269 1469 11272
rect 1432 11269 1433 11274
rect 1471 11269 1472 11274
rect 1436 11269 1437 11276
rect 1483 11269 1484 11276
rect 1439 11269 1440 11278
rect 1486 11269 1487 11278
rect 1443 11269 1444 11280
rect 1456 11269 1457 11280
rect 1446 11269 1447 11282
rect 1474 11269 1475 11282
rect 1450 11269 1451 11284
rect 1555 11269 1556 11284
rect 1453 11269 1454 11286
rect 1525 11269 1526 11286
rect 1465 11269 1466 11288
rect 1629 11269 1630 11288
rect 1477 11289 1478 11322
rect 1519 11269 1520 11290
rect 1480 11291 1481 11322
rect 1534 11269 1535 11292
rect 1489 11269 1490 11294
rect 1498 11269 1499 11294
rect 1489 11295 1490 11322
rect 1585 11269 1586 11296
rect 1492 11269 1493 11298
rect 1495 11269 1496 11298
rect 1492 11299 1493 11322
rect 1588 11269 1589 11300
rect 1501 11269 1502 11302
rect 1507 11269 1508 11302
rect 1504 11269 1505 11304
rect 1513 11269 1514 11304
rect 1546 11269 1547 11304
rect 1603 11269 1604 11304
rect 1561 11269 1562 11306
rect 1632 11269 1633 11306
rect 1564 11269 1565 11308
rect 1609 11269 1610 11308
rect 1573 11269 1574 11310
rect 1619 11269 1620 11310
rect 1576 11269 1577 11312
rect 1616 11269 1617 11312
rect 1579 11269 1580 11314
rect 1612 11269 1613 11314
rect 1582 11269 1583 11316
rect 1606 11269 1607 11316
rect 1597 11269 1598 11318
rect 1626 11269 1627 11318
rect 1600 11269 1601 11320
rect 1623 11269 1624 11320
rect 1477 11326 1478 11329
rect 1492 11326 1493 11329
rect 1480 11326 1481 11331
rect 1489 11326 1490 11331
<< via >>
rect 1423 683 1424 684
rect 1561 683 1562 684
rect 1426 685 1427 686
rect 1594 685 1595 686
rect 1430 687 1431 688
rect 1437 687 1438 688
rect 1433 689 1434 690
rect 1449 689 1450 690
rect 1440 691 1441 692
rect 1458 691 1459 692
rect 1443 693 1444 694
rect 1486 693 1487 694
rect 1446 695 1447 696
rect 1489 695 1490 696
rect 1452 697 1453 698
rect 1597 697 1598 698
rect 1455 699 1456 700
rect 1492 699 1493 700
rect 1461 701 1462 702
rect 1498 701 1499 702
rect 1464 703 1465 704
rect 1567 703 1568 704
rect 1468 705 1469 706
rect 1516 705 1517 706
rect 1471 707 1472 708
rect 1555 707 1556 708
rect 1495 709 1496 710
rect 1629 709 1630 710
rect 1507 711 1508 712
rect 1519 711 1520 712
rect 1510 713 1511 714
rect 1513 713 1514 714
rect 1525 713 1526 714
rect 1600 713 1601 714
rect 1543 715 1544 716
rect 1606 715 1607 716
rect 1546 717 1547 718
rect 1549 717 1550 718
rect 1552 717 1553 718
rect 1618 717 1619 718
rect 1558 719 1559 720
rect 1636 719 1637 720
rect 1564 721 1565 722
rect 1632 721 1633 722
rect 1579 723 1580 724
rect 1639 723 1640 724
rect 1582 725 1583 726
rect 1622 725 1623 726
rect 1603 727 1604 728
rect 1609 727 1610 728
rect 1612 727 1613 728
rect 1625 727 1626 728
rect 1615 729 1616 730
rect 1642 729 1643 730
rect 1423 739 1424 740
rect 1682 739 1683 740
rect 1423 741 1424 742
rect 1685 741 1686 742
rect 1426 743 1427 744
rect 1721 743 1722 744
rect 1426 745 1427 746
rect 1724 745 1725 746
rect 1430 747 1431 748
rect 1709 747 1710 748
rect 1430 749 1431 750
rect 1679 749 1680 750
rect 1433 751 1434 752
rect 1649 751 1650 752
rect 1433 753 1434 754
rect 1667 753 1668 754
rect 1437 755 1438 756
rect 1589 755 1590 756
rect 1436 757 1437 758
rect 2029 757 2030 758
rect 1440 759 1441 760
rect 1688 759 1689 760
rect 1439 761 1440 762
rect 1805 761 1806 762
rect 1443 763 1444 764
rect 1715 763 1716 764
rect 1443 765 1444 766
rect 1706 765 1707 766
rect 1446 767 1447 768
rect 1922 767 1923 768
rect 1446 769 1447 770
rect 1634 769 1635 770
rect 1455 771 1456 772
rect 1961 771 1962 772
rect 1464 773 1465 774
rect 1895 773 1896 774
rect 1465 775 1466 776
rect 1661 775 1662 776
rect 1468 777 1469 778
rect 1733 777 1734 778
rect 1471 779 1472 780
rect 1781 779 1782 780
rect 1474 781 1475 782
rect 1964 781 1965 782
rect 1481 783 1482 784
rect 1541 783 1542 784
rect 1484 785 1485 786
rect 1535 785 1536 786
rect 1486 787 1487 788
rect 1703 787 1704 788
rect 1489 789 1490 790
rect 1697 789 1698 790
rect 1505 791 1506 792
rect 1597 791 1598 792
rect 1507 793 1508 794
rect 1817 793 1818 794
rect 1510 795 1511 796
rect 1745 795 1746 796
rect 1511 797 1512 798
rect 1513 797 1514 798
rect 1516 797 1517 798
rect 1727 797 1728 798
rect 1477 799 1478 800
rect 1517 799 1518 800
rect 1519 799 1520 800
rect 1793 799 1794 800
rect 1523 801 1524 802
rect 1582 801 1583 802
rect 1525 803 1526 804
rect 1763 803 1764 804
rect 1543 805 1544 806
rect 1999 805 2000 806
rect 1546 807 1547 808
rect 1832 807 1833 808
rect 1547 809 1548 810
rect 1889 809 1890 810
rect 1552 811 1553 812
rect 1877 811 1878 812
rect 1555 813 1556 814
rect 1751 813 1752 814
rect 1558 815 1559 816
rect 1928 815 1929 816
rect 1561 817 1562 818
rect 1955 817 1956 818
rect 1564 819 1565 820
rect 1757 819 1758 820
rect 1567 821 1568 822
rect 1835 821 1836 822
rect 1549 823 1550 824
rect 1568 823 1569 824
rect 1550 825 1551 826
rect 1739 825 1740 826
rect 1571 827 1572 828
rect 1639 827 1640 828
rect 1579 829 1580 830
rect 1841 829 1842 830
rect 1594 831 1595 832
rect 1820 831 1821 832
rect 1458 833 1459 834
rect 1595 833 1596 834
rect 1600 833 1601 834
rect 1958 833 1959 834
rect 1601 835 1602 836
rect 1603 835 1604 836
rect 1606 835 1607 836
rect 1907 835 1908 836
rect 1609 837 1610 838
rect 1910 837 1911 838
rect 1612 839 1613 840
rect 1937 839 1938 840
rect 1615 841 1616 842
rect 1916 841 1917 842
rect 1449 843 1450 844
rect 1616 843 1617 844
rect 1450 845 1451 846
rect 1610 845 1611 846
rect 1618 845 1619 846
rect 1986 845 1987 846
rect 1452 847 1453 848
rect 1619 847 1620 848
rect 1453 849 1454 850
rect 1604 849 1605 850
rect 1622 849 1623 850
rect 2012 849 2013 850
rect 1625 851 1626 852
rect 1799 851 1800 852
rect 1492 853 1493 854
rect 1625 853 1626 854
rect 1493 855 1494 856
rect 1952 855 1953 856
rect 1629 857 1630 858
rect 1691 857 1692 858
rect 1632 859 1633 860
rect 1769 859 1770 860
rect 1495 861 1496 862
rect 1631 861 1632 862
rect 1496 863 1497 864
rect 1829 863 1830 864
rect 1636 865 1637 866
rect 1736 865 1737 866
rect 1498 867 1499 868
rect 1637 867 1638 868
rect 1642 867 1643 868
rect 2009 867 2010 868
rect 1461 869 1462 870
rect 1643 869 1644 870
rect 1462 871 1463 872
rect 1931 871 1932 872
rect 1655 873 1656 874
rect 2032 873 2033 874
rect 1673 875 1674 876
rect 1996 875 1997 876
rect 1775 877 1776 878
rect 1967 877 1968 878
rect 1787 879 1788 880
rect 1971 879 1972 880
rect 1811 881 1812 882
rect 2015 881 2016 882
rect 1847 883 1848 884
rect 1992 883 1993 884
rect 1853 885 1854 886
rect 1989 885 1990 886
rect 1859 887 1860 888
rect 2022 887 2023 888
rect 1913 889 1914 890
rect 1919 889 1920 890
rect 1925 889 1926 890
rect 2036 889 2037 890
rect 1934 891 1935 892
rect 2039 891 2040 892
rect 1940 893 1941 894
rect 2018 893 2019 894
rect 1943 895 1944 896
rect 2006 895 2007 896
rect 1974 897 1975 898
rect 2025 897 2026 898
rect 1977 899 1978 900
rect 2003 899 2004 900
rect 1417 908 1418 909
rect 1556 908 1557 909
rect 1430 910 1431 911
rect 1643 910 1644 911
rect 1443 912 1444 913
rect 1901 912 1902 913
rect 1448 914 1449 915
rect 2288 914 2289 915
rect 1450 916 1451 917
rect 2219 916 2220 917
rect 1455 918 1456 919
rect 1574 918 1575 919
rect 1459 920 1460 921
rect 1631 920 1632 921
rect 1474 922 1475 923
rect 1526 922 1527 923
rect 1477 924 1478 925
rect 1511 924 1512 925
rect 1481 926 1482 927
rect 2063 926 2064 927
rect 1484 928 1485 929
rect 2213 928 2214 929
rect 1483 930 1484 931
rect 1568 930 1569 931
rect 1486 932 1487 933
rect 1943 932 1944 933
rect 1490 934 1491 935
rect 1853 934 1854 935
rect 1493 936 1494 937
rect 2159 936 2160 937
rect 1474 938 1475 939
rect 1493 938 1494 939
rect 1502 938 1503 939
rect 2240 938 2241 939
rect 1505 940 1506 941
rect 1514 940 1515 941
rect 1505 942 1506 943
rect 2237 942 2238 943
rect 1517 944 1518 945
rect 1532 944 1533 945
rect 1520 946 1521 947
rect 1523 946 1524 947
rect 1535 946 1536 947
rect 2111 946 2112 947
rect 1541 948 1542 949
rect 2129 948 2130 949
rect 1547 950 1548 951
rect 1910 950 1911 951
rect 1550 952 1551 953
rect 2183 952 2184 953
rect 1420 954 1421 955
rect 1550 954 1551 955
rect 1586 954 1587 955
rect 1616 954 1617 955
rect 1592 956 1593 957
rect 2276 956 2277 957
rect 1601 958 1602 959
rect 1712 958 1713 959
rect 1589 960 1590 961
rect 1601 960 1602 961
rect 1496 962 1497 963
rect 1589 962 1590 963
rect 1607 962 1608 963
rect 1673 962 1674 963
rect 1613 964 1614 965
rect 1679 964 1680 965
rect 1595 966 1596 967
rect 1679 966 1680 967
rect 1595 968 1596 969
rect 2282 968 2283 969
rect 1619 970 1620 971
rect 1883 970 1884 971
rect 1619 972 1620 973
rect 1685 972 1686 973
rect 1439 974 1440 975
rect 1685 974 1686 975
rect 1438 976 1439 977
rect 1568 976 1569 977
rect 1625 976 1626 977
rect 2345 976 2346 977
rect 1625 978 1626 979
rect 1703 978 1704 979
rect 1423 980 1424 981
rect 1703 980 1704 981
rect 1424 982 1425 983
rect 1979 982 1980 983
rect 1631 984 1632 985
rect 1721 984 1722 985
rect 1637 986 1638 987
rect 2048 986 2049 987
rect 1471 988 1472 989
rect 1637 988 1638 989
rect 1643 988 1644 989
rect 1697 988 1698 989
rect 1649 990 1650 991
rect 1673 990 1674 991
rect 1649 992 1650 993
rect 1667 992 1668 993
rect 1667 994 1668 995
rect 2374 994 2375 995
rect 1676 996 1677 997
rect 1682 996 1683 997
rect 1691 996 1692 997
rect 1865 996 1866 997
rect 1697 998 1698 999
rect 1769 998 1770 999
rect 1709 1000 1710 1001
rect 1871 1000 1872 1001
rect 1436 1002 1437 1003
rect 1709 1002 1710 1003
rect 1721 1002 1722 1003
rect 1757 1002 1758 1003
rect 1724 1004 1725 1005
rect 2045 1004 2046 1005
rect 1739 1006 1740 1007
rect 2177 1006 2178 1007
rect 1727 1008 1728 1009
rect 1739 1008 1740 1009
rect 1727 1010 1728 1011
rect 2424 1010 2425 1011
rect 1745 1012 1746 1013
rect 2093 1012 2094 1013
rect 1431 1014 1432 1015
rect 1745 1014 1746 1015
rect 1751 1014 1752 1015
rect 1823 1014 1824 1015
rect 1733 1016 1734 1017
rect 1751 1016 1752 1017
rect 1688 1018 1689 1019
rect 1733 1018 1734 1019
rect 1757 1018 1758 1019
rect 1775 1018 1776 1019
rect 1465 1020 1466 1021
rect 1775 1020 1776 1021
rect 1769 1022 1770 1023
rect 2015 1022 2016 1023
rect 1426 1024 1427 1025
rect 2015 1024 2016 1025
rect 1427 1026 1428 1027
rect 1598 1026 1599 1027
rect 1781 1026 1782 1027
rect 1853 1026 1854 1027
rect 1793 1028 1794 1029
rect 2069 1028 2070 1029
rect 1793 1030 1794 1031
rect 2364 1030 2365 1031
rect 1817 1032 1818 1033
rect 2087 1032 2088 1033
rect 1462 1034 1463 1035
rect 1817 1034 1818 1035
rect 1462 1036 1463 1037
rect 2324 1036 2325 1037
rect 1820 1038 1821 1039
rect 2216 1038 2217 1039
rect 1829 1040 1830 1041
rect 2153 1040 2154 1041
rect 1763 1042 1764 1043
rect 1829 1042 1830 1043
rect 1763 1044 1764 1045
rect 2371 1044 2372 1045
rect 1832 1046 1833 1047
rect 2165 1046 2166 1047
rect 1835 1048 1836 1049
rect 2141 1048 2142 1049
rect 1787 1050 1788 1051
rect 1835 1050 1836 1051
rect 1787 1052 1788 1053
rect 1811 1052 1812 1053
rect 1661 1054 1662 1055
rect 1811 1054 1812 1055
rect 1859 1054 1860 1055
rect 2051 1054 2052 1055
rect 1859 1056 1860 1057
rect 2022 1056 2023 1057
rect 1706 1058 1707 1059
rect 2021 1058 2022 1059
rect 1877 1060 1878 1061
rect 2099 1060 2100 1061
rect 1805 1062 1806 1063
rect 1877 1062 1878 1063
rect 1715 1064 1716 1065
rect 1805 1064 1806 1065
rect 1715 1066 1716 1067
rect 2421 1066 2422 1067
rect 1889 1068 1890 1069
rect 2171 1068 2172 1069
rect 1799 1070 1800 1071
rect 1889 1070 1890 1071
rect 1799 1072 1800 1073
rect 2367 1072 2368 1073
rect 1895 1074 1896 1075
rect 2081 1074 2082 1075
rect 1895 1076 1896 1077
rect 1967 1076 1968 1077
rect 1907 1078 1908 1079
rect 2321 1078 2322 1079
rect 1571 1080 1572 1081
rect 1907 1080 1908 1081
rect 1913 1080 1914 1081
rect 2442 1080 2443 1081
rect 1913 1082 1914 1083
rect 1928 1082 1929 1083
rect 1916 1084 1917 1085
rect 2105 1084 2106 1085
rect 1919 1086 1920 1087
rect 2255 1086 2256 1087
rect 1655 1088 1656 1089
rect 1919 1088 1920 1089
rect 1433 1090 1434 1091
rect 1655 1090 1656 1091
rect 1434 1092 1435 1093
rect 2327 1092 2328 1093
rect 1922 1094 1923 1095
rect 2252 1094 2253 1095
rect 1736 1096 1737 1097
rect 1922 1096 1923 1097
rect 1441 1098 1442 1099
rect 1736 1098 1737 1099
rect 1925 1098 1926 1099
rect 2291 1098 2292 1099
rect 1925 1100 1926 1101
rect 2029 1100 2030 1101
rect 1931 1102 1932 1103
rect 2438 1102 2439 1103
rect 1841 1104 1842 1105
rect 1931 1104 1932 1105
rect 1841 1106 1842 1107
rect 2018 1106 2019 1107
rect 1934 1108 1935 1109
rect 1943 1108 1944 1109
rect 1937 1110 1938 1111
rect 2330 1110 2331 1111
rect 1937 1112 1938 1113
rect 2032 1112 2033 1113
rect 1446 1114 1447 1115
rect 2033 1114 2034 1115
rect 1445 1116 1446 1117
rect 1661 1116 1662 1117
rect 1940 1116 1941 1117
rect 2123 1116 2124 1117
rect 1952 1118 1953 1119
rect 2339 1118 2340 1119
rect 1955 1120 1956 1121
rect 2075 1120 2076 1121
rect 1610 1122 1611 1123
rect 1955 1122 1956 1123
rect 1958 1122 1959 1123
rect 2258 1122 2259 1123
rect 1961 1124 1962 1125
rect 2195 1124 2196 1125
rect 1961 1126 1962 1127
rect 2389 1126 2390 1127
rect 1964 1128 1965 1129
rect 2057 1128 2058 1129
rect 1974 1130 1975 1131
rect 2294 1130 2295 1131
rect 1604 1132 1605 1133
rect 1973 1132 1974 1133
rect 1977 1132 1978 1133
rect 2333 1132 2334 1133
rect 1986 1134 1987 1135
rect 2249 1134 2250 1135
rect 1847 1136 1848 1137
rect 1985 1136 1986 1137
rect 1847 1138 1848 1139
rect 1971 1138 1972 1139
rect 1992 1138 1993 1139
rect 2027 1138 2028 1139
rect 1991 1140 1992 1141
rect 1999 1140 2000 1141
rect 1996 1142 1997 1143
rect 2234 1142 2235 1143
rect 1997 1144 1998 1145
rect 2348 1144 2349 1145
rect 2003 1146 2004 1147
rect 2201 1146 2202 1147
rect 1989 1148 1990 1149
rect 2003 1148 2004 1149
rect 2006 1148 2007 1149
rect 2207 1148 2208 1149
rect 2009 1150 2010 1151
rect 2358 1150 2359 1151
rect 1453 1152 1454 1153
rect 2009 1152 2010 1153
rect 1452 1154 1453 1155
rect 1580 1154 1581 1155
rect 2012 1154 2013 1155
rect 2361 1154 2362 1155
rect 1634 1156 1635 1157
rect 2012 1156 2013 1157
rect 2025 1156 2026 1157
rect 2117 1156 2118 1157
rect 2039 1158 2040 1159
rect 2138 1158 2139 1159
rect 2036 1160 2037 1161
rect 2039 1160 2040 1161
rect 2036 1162 2037 1163
rect 2431 1162 2432 1163
rect 2135 1164 2136 1165
rect 2435 1164 2436 1165
rect 2189 1166 2190 1167
rect 2445 1166 2446 1167
rect 2231 1168 2232 1169
rect 2428 1168 2429 1169
rect 2297 1170 2298 1171
rect 2352 1170 2353 1171
rect 2336 1172 2337 1173
rect 2392 1172 2393 1173
rect 2342 1174 2343 1175
rect 2355 1174 2356 1175
rect 2383 1174 2384 1175
rect 2410 1174 2411 1175
rect 2386 1176 2387 1177
rect 2407 1176 2408 1177
rect 2401 1178 2402 1179
rect 2417 1178 2418 1179
rect 2404 1180 2405 1181
rect 2414 1180 2415 1181
rect 1417 1189 1418 1190
rect 1589 1189 1590 1190
rect 1417 1191 1418 1192
rect 1967 1191 1968 1192
rect 1420 1193 1421 1194
rect 2066 1193 2067 1194
rect 1427 1195 1428 1196
rect 2282 1195 2283 1196
rect 1427 1197 1428 1198
rect 2060 1197 2061 1198
rect 1434 1199 1435 1200
rect 1739 1199 1740 1200
rect 1438 1201 1439 1202
rect 2054 1201 2055 1202
rect 1438 1203 1439 1204
rect 1655 1203 1656 1204
rect 1448 1205 1449 1206
rect 2583 1205 2584 1206
rect 1448 1207 1449 1208
rect 1835 1207 1836 1208
rect 1455 1209 1456 1210
rect 2036 1209 2037 1210
rect 1455 1211 1456 1212
rect 1571 1211 1572 1212
rect 1462 1213 1463 1214
rect 2078 1213 2079 1214
rect 1466 1215 1467 1216
rect 1631 1215 1632 1216
rect 1474 1217 1475 1218
rect 2252 1217 2253 1218
rect 1473 1219 1474 1220
rect 2156 1219 2157 1220
rect 1476 1221 1477 1222
rect 2669 1221 2670 1222
rect 1480 1223 1481 1224
rect 1520 1223 1521 1224
rect 1483 1225 1484 1226
rect 1901 1225 1902 1226
rect 1483 1227 1484 1228
rect 1589 1227 1590 1228
rect 1490 1229 1491 1230
rect 1973 1229 1974 1230
rect 1471 1231 1472 1232
rect 1973 1231 1974 1232
rect 1493 1233 1494 1234
rect 1835 1233 1836 1234
rect 1502 1235 1503 1236
rect 1886 1235 1887 1236
rect 1505 1237 1506 1238
rect 1592 1237 1593 1238
rect 1514 1239 1515 1240
rect 1583 1239 1584 1240
rect 1523 1241 1524 1242
rect 1676 1241 1677 1242
rect 1529 1243 1530 1244
rect 2549 1243 2550 1244
rect 1547 1245 1548 1246
rect 1922 1245 1923 1246
rect 1550 1247 1551 1248
rect 1970 1247 1971 1248
rect 1559 1249 1560 1250
rect 2352 1249 2353 1250
rect 1577 1251 1578 1252
rect 2324 1251 2325 1252
rect 1631 1253 1632 1254
rect 2237 1253 2238 1254
rect 1643 1255 1644 1256
rect 2421 1255 2422 1256
rect 1712 1257 1713 1258
rect 2102 1257 2103 1258
rect 1781 1259 1782 1260
rect 2015 1259 2016 1260
rect 1486 1261 1487 1262
rect 2015 1261 2016 1262
rect 1487 1263 1488 1264
rect 2057 1263 2058 1264
rect 1598 1265 1599 1266
rect 2057 1265 2058 1266
rect 1793 1267 1794 1268
rect 2225 1267 2226 1268
rect 1793 1269 1794 1270
rect 2189 1269 2190 1270
rect 1757 1271 1758 1272
rect 2189 1271 2190 1272
rect 1757 1273 1758 1274
rect 2021 1273 2022 1274
rect 1829 1275 1830 1276
rect 2367 1275 2368 1276
rect 1829 1277 1830 1278
rect 2087 1277 2088 1278
rect 1685 1279 1686 1280
rect 2087 1279 2088 1280
rect 1685 1281 1686 1282
rect 2213 1281 2214 1282
rect 1841 1283 1842 1284
rect 2642 1283 2643 1284
rect 1841 1285 1842 1286
rect 1955 1285 1956 1286
rect 1847 1287 1848 1288
rect 2243 1287 2244 1288
rect 1459 1289 1460 1290
rect 1847 1289 1848 1290
rect 1459 1291 1460 1292
rect 2063 1291 2064 1292
rect 1673 1293 1674 1294
rect 2063 1293 2064 1294
rect 1574 1295 1575 1296
rect 1673 1295 1674 1296
rect 1859 1295 1860 1296
rect 2237 1295 2238 1296
rect 1859 1297 1860 1298
rect 2009 1297 2010 1298
rect 1424 1299 1425 1300
rect 2009 1299 2010 1300
rect 1424 1301 1425 1302
rect 1499 1301 1500 1302
rect 1889 1301 1890 1302
rect 2374 1301 2375 1302
rect 1595 1303 1596 1304
rect 2375 1303 2376 1304
rect 1595 1305 1596 1306
rect 2276 1305 2277 1306
rect 1889 1307 1890 1308
rect 2099 1307 2100 1308
rect 1703 1309 1704 1310
rect 2099 1309 2100 1310
rect 1703 1311 1704 1312
rect 2111 1311 2112 1312
rect 1895 1313 1896 1314
rect 2213 1313 2214 1314
rect 1895 1315 1896 1316
rect 2048 1315 2049 1316
rect 1901 1317 1902 1318
rect 1919 1317 1920 1318
rect 1420 1319 1421 1320
rect 1919 1319 1920 1320
rect 1925 1319 1926 1320
rect 2285 1319 2286 1320
rect 1865 1321 1866 1322
rect 1925 1321 1926 1322
rect 1865 1323 1866 1324
rect 2093 1323 2094 1324
rect 1637 1325 1638 1326
rect 2093 1325 2094 1326
rect 1452 1327 1453 1328
rect 1637 1327 1638 1328
rect 1452 1329 1453 1330
rect 1907 1329 1908 1330
rect 1871 1331 1872 1332
rect 1907 1331 1908 1332
rect 1727 1333 1728 1334
rect 1871 1333 1872 1334
rect 1727 1335 1728 1336
rect 2153 1335 2154 1336
rect 1751 1337 1752 1338
rect 2153 1337 2154 1338
rect 1751 1339 1752 1340
rect 2033 1339 2034 1340
rect 1613 1341 1614 1342
rect 2033 1341 2034 1342
rect 1613 1343 1614 1344
rect 2240 1343 2241 1344
rect 1931 1345 1932 1346
rect 2279 1345 2280 1346
rect 1931 1347 1932 1348
rect 2105 1347 2106 1348
rect 1943 1349 1944 1350
rect 2303 1349 2304 1350
rect 1943 1351 1944 1352
rect 2027 1351 2028 1352
rect 1949 1353 1950 1354
rect 2543 1353 2544 1354
rect 1985 1355 1986 1356
rect 2027 1355 2028 1356
rect 1763 1357 1764 1358
rect 1985 1357 1986 1358
rect 1763 1359 1764 1360
rect 2177 1359 2178 1360
rect 1715 1361 1716 1362
rect 2177 1361 2178 1362
rect 1715 1363 1716 1364
rect 2219 1363 2220 1364
rect 1787 1365 1788 1366
rect 2219 1365 2220 1366
rect 1431 1367 1432 1368
rect 1787 1367 1788 1368
rect 1431 1369 1432 1370
rect 1505 1369 1506 1370
rect 1991 1369 1992 1370
rect 2315 1369 2316 1370
rect 1991 1371 1992 1372
rect 2635 1371 2636 1372
rect 2003 1373 2004 1374
rect 2111 1373 2112 1374
rect 1775 1375 1776 1376
rect 2003 1375 2004 1376
rect 1775 1377 1776 1378
rect 2183 1377 2184 1378
rect 2012 1379 2013 1380
rect 2024 1379 2025 1380
rect 2045 1379 2046 1380
rect 2108 1379 2109 1380
rect 1607 1381 1608 1382
rect 2045 1381 2046 1382
rect 2105 1381 2106 1382
rect 2371 1381 2372 1382
rect 2117 1383 2118 1384
rect 2381 1383 2382 1384
rect 1805 1385 1806 1386
rect 2117 1385 2118 1386
rect 1805 1387 1806 1388
rect 2069 1387 2070 1388
rect 1709 1389 1710 1390
rect 2069 1389 2070 1390
rect 1709 1391 1710 1392
rect 2129 1391 2130 1392
rect 2051 1393 2052 1394
rect 2129 1393 2130 1394
rect 1619 1395 1620 1396
rect 2051 1395 2052 1396
rect 1526 1397 1527 1398
rect 1619 1397 1620 1398
rect 2123 1397 2124 1398
rect 2351 1397 2352 1398
rect 1661 1399 1662 1400
rect 2123 1399 2124 1400
rect 1556 1401 1557 1402
rect 1661 1401 1662 1402
rect 2135 1401 2136 1402
rect 2420 1401 2421 1402
rect 1667 1403 1668 1404
rect 2135 1403 2136 1404
rect 1568 1405 1569 1406
rect 1667 1405 1668 1406
rect 2138 1405 2139 1406
rect 2309 1405 2310 1406
rect 2141 1407 2142 1408
rect 2369 1407 2370 1408
rect 1913 1409 1914 1410
rect 2141 1409 2142 1410
rect 1586 1411 1587 1412
rect 1913 1411 1914 1412
rect 2183 1411 2184 1412
rect 2392 1411 2393 1412
rect 2195 1413 2196 1414
rect 2453 1413 2454 1414
rect 1769 1415 1770 1416
rect 2195 1415 2196 1416
rect 1462 1417 1463 1418
rect 1769 1417 1770 1418
rect 2198 1417 2199 1418
rect 2216 1417 2217 1418
rect 2204 1419 2205 1420
rect 2255 1419 2256 1420
rect 1961 1421 1962 1422
rect 2255 1421 2256 1422
rect 1961 1423 1962 1424
rect 2540 1423 2541 1424
rect 2207 1425 2208 1426
rect 2447 1425 2448 1426
rect 1877 1427 1878 1428
rect 2207 1427 2208 1428
rect 1877 1429 1878 1430
rect 1883 1429 1884 1430
rect 1490 1431 1491 1432
rect 1883 1431 1884 1432
rect 2231 1431 2232 1432
rect 2477 1431 2478 1432
rect 1799 1433 1800 1434
rect 2231 1433 2232 1434
rect 2249 1433 2250 1434
rect 2501 1433 2502 1434
rect 1853 1435 1854 1436
rect 2249 1435 2250 1436
rect 2258 1435 2259 1436
rect 2507 1435 2508 1436
rect 2261 1437 2262 1438
rect 2336 1437 2337 1438
rect 2267 1439 2268 1440
rect 2639 1439 2640 1440
rect 2273 1441 2274 1442
rect 2389 1441 2390 1442
rect 2288 1443 2289 1444
rect 2495 1443 2496 1444
rect 2291 1445 2292 1446
rect 2498 1445 2499 1446
rect 2291 1447 2292 1448
rect 2632 1447 2633 1448
rect 2294 1449 2295 1450
rect 2537 1449 2538 1450
rect 2297 1451 2298 1452
rect 2513 1451 2514 1452
rect 1937 1453 1938 1454
rect 2297 1453 2298 1454
rect 1817 1455 1818 1456
rect 1937 1455 1938 1456
rect 1679 1457 1680 1458
rect 1817 1457 1818 1458
rect 1580 1459 1581 1460
rect 1679 1459 1680 1460
rect 2321 1459 2322 1460
rect 2378 1459 2379 1460
rect 1997 1461 1998 1462
rect 2321 1461 2322 1462
rect 1979 1463 1980 1464
rect 1997 1463 1998 1464
rect 1811 1465 1812 1466
rect 1979 1465 1980 1466
rect 1601 1467 1602 1468
rect 1811 1467 1812 1468
rect 1441 1469 1442 1470
rect 1601 1469 1602 1470
rect 1441 1471 1442 1472
rect 1955 1471 1956 1472
rect 2327 1471 2328 1472
rect 2564 1471 2565 1472
rect 2327 1473 2328 1474
rect 2703 1473 2704 1474
rect 2330 1475 2331 1476
rect 2465 1475 2466 1476
rect 2333 1477 2334 1478
rect 2570 1477 2571 1478
rect 2075 1479 2076 1480
rect 2333 1479 2334 1480
rect 1625 1481 1626 1482
rect 2075 1481 2076 1482
rect 1532 1483 1533 1484
rect 1625 1483 1626 1484
rect 1532 1485 1533 1486
rect 2147 1485 2148 1486
rect 2339 1485 2340 1486
rect 2546 1485 2547 1486
rect 2039 1487 2040 1488
rect 2339 1487 2340 1488
rect 1649 1489 1650 1490
rect 2039 1489 2040 1490
rect 1649 1491 1650 1492
rect 1736 1491 1737 1492
rect 2342 1491 2343 1492
rect 2519 1491 2520 1492
rect 2345 1493 2346 1494
rect 2687 1493 2688 1494
rect 2345 1495 2346 1496
rect 2579 1495 2580 1496
rect 2348 1497 2349 1498
rect 2573 1497 2574 1498
rect 2355 1499 2356 1500
rect 2525 1499 2526 1500
rect 2358 1501 2359 1502
rect 2595 1501 2596 1502
rect 1469 1503 1470 1504
rect 2357 1503 2358 1504
rect 2361 1503 2362 1504
rect 2531 1503 2532 1504
rect 2364 1505 2365 1506
rect 2424 1505 2425 1506
rect 2081 1507 2082 1508
rect 2363 1507 2364 1508
rect 1445 1509 1446 1510
rect 2081 1509 2082 1510
rect 1445 1511 1446 1512
rect 2021 1511 2022 1512
rect 2234 1511 2235 1512
rect 2423 1511 2424 1512
rect 2383 1513 2384 1514
rect 2435 1513 2436 1514
rect 2386 1515 2387 1516
rect 2607 1515 2608 1516
rect 2393 1517 2394 1518
rect 2700 1517 2701 1518
rect 2399 1519 2400 1520
rect 2445 1519 2446 1520
rect 2401 1521 2402 1522
rect 2651 1521 2652 1522
rect 2404 1523 2405 1524
rect 2645 1523 2646 1524
rect 2405 1525 2406 1526
rect 2710 1525 2711 1526
rect 2407 1527 2408 1528
rect 2622 1527 2623 1528
rect 2410 1529 2411 1530
rect 2619 1529 2620 1530
rect 2414 1531 2415 1532
rect 2666 1531 2667 1532
rect 2417 1533 2418 1534
rect 2663 1533 2664 1534
rect 2417 1535 2418 1536
rect 2714 1535 2715 1536
rect 2428 1537 2429 1538
rect 2483 1537 2484 1538
rect 2431 1539 2432 1540
rect 2486 1539 2487 1540
rect 2438 1541 2439 1542
rect 2707 1541 2708 1542
rect 2442 1543 2443 1544
rect 2504 1543 2505 1544
rect 2201 1545 2202 1546
rect 2441 1545 2442 1546
rect 1823 1547 1824 1548
rect 2201 1547 2202 1548
rect 1733 1549 1734 1550
rect 1823 1549 1824 1550
rect 1733 1551 1734 1552
rect 2159 1551 2160 1552
rect 1697 1553 1698 1554
rect 2159 1553 2160 1554
rect 1434 1555 1435 1556
rect 1697 1555 1698 1556
rect 2459 1555 2460 1556
rect 2672 1555 2673 1556
rect 2489 1557 2490 1558
rect 2586 1557 2587 1558
rect 2558 1559 2559 1560
rect 2723 1559 2724 1560
rect 2561 1561 2562 1562
rect 2720 1561 2721 1562
rect 2576 1563 2577 1564
rect 2717 1563 2718 1564
rect 2601 1565 2602 1566
rect 2628 1565 2629 1566
rect 2604 1567 2605 1568
rect 2625 1567 2626 1568
rect 2675 1567 2676 1568
rect 2693 1567 2694 1568
rect 2690 1569 2691 1570
rect 2696 1569 2697 1570
rect 1424 1578 1425 1579
rect 1517 1578 1518 1579
rect 1417 1580 1418 1581
rect 1424 1580 1425 1581
rect 1427 1580 1428 1581
rect 2174 1580 2175 1581
rect 1431 1582 1432 1583
rect 2045 1582 2046 1583
rect 1445 1584 1446 1585
rect 1931 1584 1932 1585
rect 1448 1586 1449 1587
rect 1469 1586 1470 1587
rect 1448 1588 1449 1589
rect 1619 1588 1620 1589
rect 1452 1590 1453 1591
rect 1787 1590 1788 1591
rect 1452 1592 1453 1593
rect 1865 1592 1866 1593
rect 1455 1594 1456 1595
rect 1781 1594 1782 1595
rect 1466 1596 1467 1597
rect 2318 1596 2319 1597
rect 1476 1598 1477 1599
rect 2246 1598 2247 1599
rect 1469 1600 1470 1601
rect 1476 1600 1477 1601
rect 1483 1600 1484 1601
rect 1583 1600 1584 1601
rect 1485 1602 1486 1603
rect 2123 1602 2124 1603
rect 1487 1604 1488 1605
rect 1883 1604 1884 1605
rect 1502 1606 1503 1607
rect 2369 1606 2370 1607
rect 1505 1608 1506 1609
rect 1541 1608 1542 1609
rect 1532 1610 1533 1611
rect 2900 1610 2901 1611
rect 1565 1612 1566 1613
rect 2078 1612 2079 1613
rect 1577 1614 1578 1615
rect 1607 1614 1608 1615
rect 1547 1616 1548 1617
rect 1577 1616 1578 1617
rect 1473 1618 1474 1619
rect 1547 1618 1548 1619
rect 1473 1620 1474 1621
rect 2525 1620 2526 1621
rect 1625 1622 1626 1623
rect 1655 1622 1656 1623
rect 1480 1624 1481 1625
rect 1625 1624 1626 1625
rect 1643 1624 1644 1625
rect 1886 1624 1887 1625
rect 1661 1626 1662 1627
rect 1691 1626 1692 1627
rect 1631 1628 1632 1629
rect 1661 1628 1662 1629
rect 1589 1630 1590 1631
rect 1631 1630 1632 1631
rect 1679 1630 1680 1631
rect 2778 1630 2779 1631
rect 1667 1632 1668 1633
rect 1679 1632 1680 1633
rect 1709 1632 1710 1633
rect 1739 1632 1740 1633
rect 1685 1634 1686 1635
rect 1709 1634 1710 1635
rect 1745 1634 1746 1635
rect 1781 1634 1782 1635
rect 1715 1636 1716 1637
rect 1745 1636 1746 1637
rect 1751 1636 1752 1637
rect 1799 1636 1800 1637
rect 1721 1638 1722 1639
rect 1751 1638 1752 1639
rect 1703 1640 1704 1641
rect 1721 1640 1722 1641
rect 1673 1642 1674 1643
rect 1703 1642 1704 1643
rect 1649 1644 1650 1645
rect 1673 1644 1674 1645
rect 1613 1646 1614 1647
rect 1649 1646 1650 1647
rect 1571 1648 1572 1649
rect 1613 1648 1614 1649
rect 1571 1650 1572 1651
rect 2156 1650 2157 1651
rect 1763 1652 1764 1653
rect 1787 1652 1788 1653
rect 1727 1654 1728 1655
rect 1763 1654 1764 1655
rect 1697 1656 1698 1657
rect 1727 1656 1728 1657
rect 1637 1658 1638 1659
rect 1697 1658 1698 1659
rect 1595 1660 1596 1661
rect 1637 1660 1638 1661
rect 1559 1662 1560 1663
rect 1595 1662 1596 1663
rect 1523 1664 1524 1665
rect 1559 1664 1560 1665
rect 1523 1666 1524 1667
rect 2060 1666 2061 1667
rect 1805 1668 1806 1669
rect 1883 1668 1884 1669
rect 1434 1670 1435 1671
rect 1805 1670 1806 1671
rect 1817 1670 1818 1671
rect 1853 1670 1854 1671
rect 1775 1672 1776 1673
rect 1817 1672 1818 1673
rect 1601 1674 1602 1675
rect 1775 1674 1776 1675
rect 1835 1674 1836 1675
rect 1865 1674 1866 1675
rect 1835 1676 1836 1677
rect 2867 1676 2868 1677
rect 1889 1678 1890 1679
rect 2826 1678 2827 1679
rect 1841 1680 1842 1681
rect 1889 1680 1890 1681
rect 1841 1682 1842 1683
rect 2635 1682 2636 1683
rect 1931 1684 1932 1685
rect 2291 1684 2292 1685
rect 1943 1686 1944 1687
rect 2543 1686 2544 1687
rect 1895 1688 1896 1689
rect 1943 1688 1944 1689
rect 1970 1688 1971 1689
rect 2072 1688 2073 1689
rect 1973 1690 1974 1691
rect 2045 1690 2046 1691
rect 1793 1692 1794 1693
rect 1973 1692 1974 1693
rect 1455 1694 1456 1695
rect 1793 1694 1794 1695
rect 1991 1694 1992 1695
rect 2771 1694 2772 1695
rect 1937 1696 1938 1697
rect 1991 1696 1992 1697
rect 1490 1698 1491 1699
rect 1937 1698 1938 1699
rect 2021 1698 2022 1699
rect 2123 1698 2124 1699
rect 1979 1700 1980 1701
rect 2021 1700 2022 1701
rect 1417 1702 1418 1703
rect 1979 1702 1980 1703
rect 2054 1702 2055 1703
rect 2168 1702 2169 1703
rect 2066 1704 2067 1705
rect 2162 1704 2163 1705
rect 2108 1706 2109 1707
rect 2222 1706 2223 1707
rect 2177 1708 2178 1709
rect 2291 1708 2292 1709
rect 1441 1710 1442 1711
rect 2177 1710 2178 1711
rect 1441 1712 1442 1713
rect 1847 1712 1848 1713
rect 1811 1714 1812 1715
rect 1847 1714 1848 1715
rect 1757 1716 1758 1717
rect 1811 1716 1812 1717
rect 2198 1716 2199 1717
rect 2324 1716 2325 1717
rect 2102 1718 2103 1719
rect 2198 1718 2199 1719
rect 2204 1718 2205 1719
rect 2270 1718 2271 1719
rect 1529 1720 1530 1721
rect 2204 1720 2205 1721
rect 1499 1722 1500 1723
rect 1529 1722 1530 1723
rect 1499 1724 1500 1725
rect 2741 1724 2742 1725
rect 2243 1726 2244 1727
rect 2369 1726 2370 1727
rect 2153 1728 2154 1729
rect 2243 1728 2244 1729
rect 2033 1730 2034 1731
rect 2153 1730 2154 1731
rect 1955 1732 1956 1733
rect 2033 1732 2034 1733
rect 1907 1734 1908 1735
rect 1955 1734 1956 1735
rect 1859 1736 1860 1737
rect 1907 1736 1908 1737
rect 1823 1738 1824 1739
rect 1859 1738 1860 1739
rect 1459 1740 1460 1741
rect 1823 1740 1824 1741
rect 1459 1742 1460 1743
rect 2126 1742 2127 1743
rect 2261 1742 2262 1743
rect 2411 1742 2412 1743
rect 2147 1744 2148 1745
rect 2261 1744 2262 1745
rect 2063 1746 2064 1747
rect 2147 1746 2148 1747
rect 1420 1748 1421 1749
rect 2063 1748 2064 1749
rect 1420 1750 1421 1751
rect 1913 1750 1914 1751
rect 1829 1752 1830 1753
rect 1913 1752 1914 1753
rect 1769 1754 1770 1755
rect 1829 1754 1830 1755
rect 1733 1756 1734 1757
rect 1769 1756 1770 1757
rect 1427 1758 1428 1759
rect 1733 1758 1734 1759
rect 2285 1758 2286 1759
rect 2429 1758 2430 1759
rect 2165 1760 2166 1761
rect 2285 1760 2286 1761
rect 2051 1762 2052 1763
rect 2165 1762 2166 1763
rect 1488 1764 1489 1765
rect 2051 1764 2052 1765
rect 2321 1764 2322 1765
rect 2435 1764 2436 1765
rect 1492 1766 1493 1767
rect 2321 1766 2322 1767
rect 2327 1766 2328 1767
rect 2471 1766 2472 1767
rect 2207 1768 2208 1769
rect 2327 1768 2328 1769
rect 2093 1770 2094 1771
rect 2207 1770 2208 1771
rect 2093 1772 2094 1773
rect 2840 1772 2841 1773
rect 2333 1774 2334 1775
rect 2579 1774 2580 1775
rect 2219 1776 2220 1777
rect 2333 1776 2334 1777
rect 2105 1778 2106 1779
rect 2219 1778 2220 1779
rect 1466 1780 1467 1781
rect 2105 1780 2106 1781
rect 2378 1780 2379 1781
rect 2492 1780 2493 1781
rect 2381 1782 2382 1783
rect 2525 1782 2526 1783
rect 2255 1784 2256 1785
rect 2381 1784 2382 1785
rect 2171 1786 2172 1787
rect 2255 1786 2256 1787
rect 2057 1788 2058 1789
rect 2171 1788 2172 1789
rect 1985 1790 1986 1791
rect 2057 1790 2058 1791
rect 1462 1792 1463 1793
rect 1985 1792 1986 1793
rect 1462 1794 1463 1795
rect 2024 1794 2025 1795
rect 2387 1794 2388 1795
rect 2775 1794 2776 1795
rect 2423 1796 2424 1797
rect 2579 1796 2580 1797
rect 2279 1798 2280 1799
rect 2423 1798 2424 1799
rect 2279 1800 2280 1801
rect 2768 1800 2769 1801
rect 2441 1802 2442 1803
rect 2707 1802 2708 1803
rect 2303 1804 2304 1805
rect 2441 1804 2442 1805
rect 2189 1806 2190 1807
rect 2303 1806 2304 1807
rect 2141 1808 2142 1809
rect 2189 1808 2190 1809
rect 2099 1810 2100 1811
rect 2141 1810 2142 1811
rect 2003 1812 2004 1813
rect 2099 1812 2100 1813
rect 1961 1814 1962 1815
rect 2003 1814 2004 1815
rect 1925 1816 1926 1817
rect 1961 1816 1962 1817
rect 1877 1818 1878 1819
rect 1925 1818 1926 1819
rect 1431 1820 1432 1821
rect 1877 1820 1878 1821
rect 2447 1820 2448 1821
rect 2555 1820 2556 1821
rect 2309 1822 2310 1823
rect 2447 1822 2448 1823
rect 2309 1824 2310 1825
rect 2918 1824 2919 1825
rect 2459 1826 2460 1827
rect 2615 1826 2616 1827
rect 2315 1828 2316 1829
rect 2459 1828 2460 1829
rect 2486 1828 2487 1829
rect 2630 1828 2631 1829
rect 2498 1830 2499 1831
rect 2583 1830 2584 1831
rect 2501 1832 2502 1833
rect 2654 1832 2655 1833
rect 2357 1834 2358 1835
rect 2501 1834 2502 1835
rect 2213 1836 2214 1837
rect 2357 1836 2358 1837
rect 2117 1838 2118 1839
rect 2213 1838 2214 1839
rect 2117 1840 2118 1841
rect 2393 1840 2394 1841
rect 2393 1842 2394 1843
rect 2639 1842 2640 1843
rect 2489 1844 2490 1845
rect 2639 1844 2640 1845
rect 2375 1846 2376 1847
rect 2489 1846 2490 1847
rect 2249 1848 2250 1849
rect 2375 1848 2376 1849
rect 2135 1850 2136 1851
rect 2249 1850 2250 1851
rect 2069 1852 2070 1853
rect 2135 1852 2136 1853
rect 1967 1854 1968 1855
rect 2069 1854 2070 1855
rect 1919 1856 1920 1857
rect 1967 1856 1968 1857
rect 1871 1858 1872 1859
rect 1919 1858 1920 1859
rect 1434 1860 1435 1861
rect 1871 1860 1872 1861
rect 2507 1860 2508 1861
rect 2657 1860 2658 1861
rect 2363 1862 2364 1863
rect 2507 1862 2508 1863
rect 2237 1864 2238 1865
rect 2363 1864 2364 1865
rect 2237 1866 2238 1867
rect 2642 1866 2643 1867
rect 2540 1868 2541 1869
rect 2672 1868 2673 1869
rect 2543 1870 2544 1871
rect 2907 1870 2908 1871
rect 2546 1872 2547 1873
rect 2744 1872 2745 1873
rect 2549 1874 2550 1875
rect 2747 1874 2748 1875
rect 2399 1876 2400 1877
rect 2549 1876 2550 1877
rect 2267 1878 2268 1879
rect 2399 1878 2400 1879
rect 2201 1880 2202 1881
rect 2267 1880 2268 1881
rect 2075 1882 2076 1883
rect 2201 1882 2202 1883
rect 2027 1884 2028 1885
rect 2075 1884 2076 1885
rect 2027 1886 2028 1887
rect 2837 1886 2838 1887
rect 2564 1888 2565 1889
rect 2756 1888 2757 1889
rect 2570 1890 2571 1891
rect 2830 1890 2831 1891
rect 2573 1892 2574 1893
rect 2632 1892 2633 1893
rect 2417 1894 2418 1895
rect 2573 1894 2574 1895
rect 2273 1896 2274 1897
rect 2417 1896 2418 1897
rect 2159 1898 2160 1899
rect 2273 1898 2274 1899
rect 2039 1900 2040 1901
rect 2159 1900 2160 1901
rect 1495 1902 1496 1903
rect 2039 1902 2040 1903
rect 2465 1902 2466 1903
rect 2633 1902 2634 1903
rect 2465 1904 2466 1905
rect 2870 1904 2871 1905
rect 2576 1906 2577 1907
rect 2911 1906 2912 1907
rect 2591 1908 2592 1909
rect 2669 1908 2670 1909
rect 2513 1910 2514 1911
rect 2669 1910 2670 1911
rect 2595 1912 2596 1913
rect 2787 1912 2788 1913
rect 2597 1914 2598 1915
rect 2823 1914 2824 1915
rect 2601 1916 2602 1917
rect 2820 1916 2821 1917
rect 2604 1918 2605 1919
rect 2781 1918 2782 1919
rect 2453 1920 2454 1921
rect 2603 1920 2604 1921
rect 2297 1922 2298 1923
rect 2453 1922 2454 1923
rect 2195 1924 2196 1925
rect 2297 1924 2298 1925
rect 2081 1926 2082 1927
rect 2195 1926 2196 1927
rect 2081 1928 2082 1929
rect 2111 1928 2112 1929
rect 2009 1930 2010 1931
rect 2111 1930 2112 1931
rect 2009 1932 2010 1933
rect 2129 1932 2130 1933
rect 2129 1934 2130 1935
rect 2904 1934 2905 1935
rect 2607 1936 2608 1937
rect 2799 1936 2800 1937
rect 2609 1938 2610 1939
rect 2717 1938 2718 1939
rect 2619 1940 2620 1941
rect 2811 1940 2812 1941
rect 2622 1942 2623 1943
rect 2814 1942 2815 1943
rect 2477 1944 2478 1945
rect 2621 1944 2622 1945
rect 2345 1946 2346 1947
rect 2477 1946 2478 1947
rect 2225 1948 2226 1949
rect 2345 1948 2346 1949
rect 2183 1950 2184 1951
rect 2225 1950 2226 1951
rect 2087 1952 2088 1953
rect 2183 1952 2184 1953
rect 2015 1954 2016 1955
rect 2087 1954 2088 1955
rect 1997 1956 1998 1957
rect 2015 1956 2016 1957
rect 1949 1958 1950 1959
rect 1997 1958 1998 1959
rect 1901 1960 1902 1961
rect 1949 1960 1950 1961
rect 1445 1962 1446 1963
rect 1901 1962 1902 1963
rect 2625 1962 2626 1963
rect 2817 1962 2818 1963
rect 2628 1964 2629 1965
rect 2925 1964 2926 1965
rect 2483 1966 2484 1967
rect 2627 1966 2628 1967
rect 2339 1968 2340 1969
rect 2483 1968 2484 1969
rect 2339 1970 2340 1971
rect 2703 1970 2704 1971
rect 2645 1972 2646 1973
rect 2843 1972 2844 1973
rect 2651 1974 2652 1975
rect 2849 1974 2850 1975
rect 2651 1976 2652 1977
rect 2928 1976 2929 1977
rect 2663 1978 2664 1979
rect 2861 1978 2862 1979
rect 2495 1980 2496 1981
rect 2663 1980 2664 1981
rect 2351 1982 2352 1983
rect 2495 1982 2496 1983
rect 2231 1984 2232 1985
rect 2351 1984 2352 1985
rect 2231 1986 2232 1987
rect 2708 1986 2709 1987
rect 2666 1988 2667 1989
rect 2864 1988 2865 1989
rect 2586 1990 2587 1991
rect 2666 1990 2667 1991
rect 2405 1992 2406 1993
rect 2585 1992 2586 1993
rect 2405 1994 2406 1995
rect 2921 1994 2922 1995
rect 2675 1996 2676 1997
rect 2873 1996 2874 1997
rect 2519 1998 2520 1999
rect 2675 1998 2676 1999
rect 2519 2000 2520 2001
rect 2897 2000 2898 2001
rect 2687 2002 2688 2003
rect 2696 2002 2697 2003
rect 2531 2004 2532 2005
rect 2696 2004 2697 2005
rect 2504 2006 2505 2007
rect 2531 2006 2532 2007
rect 2690 2006 2691 2007
rect 2894 2006 2895 2007
rect 2693 2008 2694 2009
rect 2891 2008 2892 2009
rect 2537 2010 2538 2011
rect 2693 2010 2694 2011
rect 1438 2012 1439 2013
rect 2537 2012 2538 2013
rect 1438 2014 1439 2015
rect 2315 2014 2316 2015
rect 2700 2014 2701 2015
rect 2702 2014 2703 2015
rect 2710 2014 2711 2015
rect 2879 2014 2880 2015
rect 1583 2016 1584 2017
rect 2711 2016 2712 2017
rect 2714 2016 2715 2017
rect 2765 2016 2766 2017
rect 2561 2018 2562 2019
rect 2714 2018 2715 2019
rect 2420 2020 2421 2021
rect 2561 2020 2562 2021
rect 2720 2020 2721 2021
rect 2726 2020 2727 2021
rect 2558 2022 2559 2023
rect 2720 2022 2721 2023
rect 2723 2022 2724 2023
rect 2882 2022 2883 2023
rect 2738 2024 2739 2025
rect 2914 2024 2915 2025
rect 2762 2026 2763 2027
rect 2833 2026 2834 2027
rect 1417 2035 1418 2036
rect 2103 2035 2104 2036
rect 1420 2037 1421 2038
rect 1989 2037 1990 2038
rect 1424 2039 1425 2040
rect 3018 2039 3019 2040
rect 1427 2041 1428 2042
rect 1899 2041 1900 2042
rect 1431 2043 1432 2044
rect 1490 2043 1491 2044
rect 1432 2045 1433 2046
rect 2337 2045 2338 2046
rect 1434 2047 1435 2048
rect 1865 2047 1866 2048
rect 1436 2049 1437 2050
rect 1959 2049 1960 2050
rect 1438 2051 1439 2052
rect 2165 2051 2166 2052
rect 1443 2053 1444 2054
rect 1853 2053 1854 2054
rect 1445 2055 1446 2056
rect 1689 2055 1690 2056
rect 1448 2057 1449 2058
rect 2198 2057 2199 2058
rect 1450 2059 1451 2060
rect 1733 2059 1734 2060
rect 1452 2061 1453 2062
rect 2174 2061 2175 2062
rect 1453 2063 1454 2064
rect 1779 2063 1780 2064
rect 1455 2065 1456 2066
rect 2289 2065 2290 2066
rect 1457 2067 1458 2068
rect 1821 2067 1822 2068
rect 1462 2069 1463 2070
rect 2708 2069 2709 2070
rect 1464 2071 1465 2072
rect 2199 2071 2200 2072
rect 1466 2073 1467 2074
rect 2099 2073 2100 2074
rect 1467 2075 1468 2076
rect 2057 2075 2058 2076
rect 1469 2077 1470 2078
rect 2097 2077 2098 2078
rect 1471 2079 1472 2080
rect 2121 2079 2122 2080
rect 1473 2081 1474 2082
rect 2021 2081 2022 2082
rect 1474 2083 1475 2084
rect 1673 2083 1674 2084
rect 1476 2085 1477 2086
rect 2151 2085 2152 2086
rect 1483 2087 1484 2088
rect 1803 2087 1804 2088
rect 1485 2089 1486 2090
rect 1587 2089 1588 2090
rect 1488 2091 1489 2092
rect 2379 2091 2380 2092
rect 1492 2093 1493 2094
rect 1931 2093 1932 2094
rect 1497 2095 1498 2096
rect 1607 2095 1608 2096
rect 1499 2097 1500 2098
rect 2013 2097 2014 2098
rect 1500 2099 1501 2100
rect 1611 2099 1612 2100
rect 1502 2101 1503 2102
rect 1977 2101 1978 2102
rect 1515 2103 1516 2104
rect 2126 2103 2127 2104
rect 1486 2105 1487 2106
rect 2127 2105 2128 2106
rect 1521 2107 1522 2108
rect 1547 2107 1548 2108
rect 1523 2109 1524 2110
rect 2778 2109 2779 2110
rect 1529 2111 1530 2112
rect 1533 2111 1534 2112
rect 1541 2111 1542 2112
rect 1551 2111 1552 2112
rect 1545 2113 1546 2114
rect 1565 2113 1566 2114
rect 1557 2115 1558 2116
rect 1571 2115 1572 2116
rect 1559 2117 1560 2118
rect 1569 2117 1570 2118
rect 1563 2119 1564 2120
rect 2162 2119 2163 2120
rect 1575 2121 1576 2122
rect 1577 2121 1578 2122
rect 1583 2121 1584 2122
rect 1599 2121 1600 2122
rect 1593 2123 1594 2124
rect 1595 2123 1596 2124
rect 1613 2123 1614 2124
rect 1629 2123 1630 2124
rect 1623 2125 1624 2126
rect 2318 2125 2319 2126
rect 1429 2127 1430 2128
rect 2319 2127 2320 2128
rect 1625 2129 1626 2130
rect 1641 2129 1642 2130
rect 1631 2131 1632 2132
rect 1647 2131 1648 2132
rect 1637 2133 1638 2134
rect 1653 2133 1654 2134
rect 1643 2135 1644 2136
rect 1659 2135 1660 2136
rect 1649 2137 1650 2138
rect 1671 2137 1672 2138
rect 1655 2139 1656 2140
rect 1683 2139 1684 2140
rect 1661 2141 1662 2142
rect 1665 2141 1666 2142
rect 1677 2141 1678 2142
rect 1775 2141 1776 2142
rect 1691 2143 1692 2144
rect 1737 2143 1738 2144
rect 1692 2145 1693 2146
rect 2019 2145 2020 2146
rect 1695 2147 1696 2148
rect 1709 2147 1710 2148
rect 1697 2149 1698 2150
rect 1719 2149 1720 2150
rect 1701 2151 1702 2152
rect 1721 2151 1722 2152
rect 1703 2153 1704 2154
rect 1725 2153 1726 2154
rect 1707 2155 1708 2156
rect 1739 2155 1740 2156
rect 1727 2157 1728 2158
rect 1773 2157 1774 2158
rect 1743 2159 1744 2160
rect 1745 2159 1746 2160
rect 1749 2159 1750 2160
rect 2222 2159 2223 2160
rect 1751 2161 1752 2162
rect 1785 2161 1786 2162
rect 1761 2163 1762 2164
rect 2669 2163 2670 2164
rect 1763 2165 1764 2166
rect 1809 2165 1810 2166
rect 1769 2167 1770 2168
rect 1815 2167 1816 2168
rect 1781 2169 1782 2170
rect 1827 2169 1828 2170
rect 1787 2171 1788 2172
rect 1851 2171 1852 2172
rect 1791 2173 1792 2174
rect 2666 2173 2667 2174
rect 1793 2175 1794 2176
rect 1833 2175 1834 2176
rect 1797 2177 1798 2178
rect 2633 2177 2634 2178
rect 1799 2179 1800 2180
rect 1839 2179 1840 2180
rect 1805 2181 1806 2182
rect 1869 2181 1870 2182
rect 1811 2183 1812 2184
rect 1845 2183 1846 2184
rect 1817 2185 1818 2186
rect 1875 2185 1876 2186
rect 1823 2187 1824 2188
rect 1857 2187 1858 2188
rect 1829 2189 1830 2190
rect 1863 2189 1864 2190
rect 1835 2191 1836 2192
rect 1881 2191 1882 2192
rect 1841 2193 1842 2194
rect 1887 2193 1888 2194
rect 1847 2195 1848 2196
rect 1935 2195 1936 2196
rect 1859 2197 1860 2198
rect 1941 2197 1942 2198
rect 1871 2199 1872 2200
rect 1953 2199 1954 2200
rect 1877 2201 1878 2202
rect 1965 2201 1966 2202
rect 1883 2203 1884 2204
rect 1911 2203 1912 2204
rect 1889 2205 1890 2206
rect 1929 2205 1930 2206
rect 1893 2207 1894 2208
rect 1973 2207 1974 2208
rect 1901 2209 1902 2210
rect 1983 2209 1984 2210
rect 1905 2211 1906 2212
rect 1985 2211 1986 2212
rect 1907 2213 1908 2214
rect 1947 2213 1948 2214
rect 1913 2215 1914 2216
rect 1923 2215 1924 2216
rect 1919 2217 1920 2218
rect 2007 2217 2008 2218
rect 1925 2219 1926 2220
rect 2001 2219 2002 2220
rect 1937 2221 1938 2222
rect 1995 2221 1996 2222
rect 1943 2223 1944 2224
rect 2055 2223 2056 2224
rect 1949 2225 1950 2226
rect 2025 2225 2026 2226
rect 1955 2227 1956 2228
rect 2067 2227 2068 2228
rect 1961 2229 1962 2230
rect 2079 2229 2080 2230
rect 1971 2231 1972 2232
rect 2117 2231 2118 2232
rect 1979 2233 1980 2234
rect 2109 2233 2110 2234
rect 1991 2235 1992 2236
rect 2115 2235 2116 2236
rect 1997 2237 1998 2238
rect 2043 2237 2044 2238
rect 2003 2239 2004 2240
rect 2049 2239 2050 2240
rect 2009 2241 2010 2242
rect 2031 2241 2032 2242
rect 2015 2243 2016 2244
rect 2145 2243 2146 2244
rect 2027 2245 2028 2246
rect 2157 2245 2158 2246
rect 2033 2247 2034 2248
rect 2163 2247 2164 2248
rect 2037 2249 2038 2250
rect 2093 2249 2094 2250
rect 2045 2251 2046 2252
rect 2175 2251 2176 2252
rect 2051 2253 2052 2254
rect 2181 2253 2182 2254
rect 2061 2255 2062 2256
rect 2639 2255 2640 2256
rect 2063 2257 2064 2258
rect 2187 2257 2188 2258
rect 2069 2259 2070 2260
rect 2193 2259 2194 2260
rect 2075 2261 2076 2262
rect 2577 2261 2578 2262
rect 2081 2263 2082 2264
rect 2601 2263 2602 2264
rect 2085 2265 2086 2266
rect 2477 2265 2478 2266
rect 2087 2267 2088 2268
rect 2217 2267 2218 2268
rect 2091 2269 2092 2270
rect 2768 2269 2769 2270
rect 2105 2271 2106 2272
rect 2229 2271 2230 2272
rect 2111 2273 2112 2274
rect 2235 2273 2236 2274
rect 2129 2275 2130 2276
rect 2241 2275 2242 2276
rect 2133 2277 2134 2278
rect 3012 2277 3013 2278
rect 2139 2279 2140 2280
rect 2471 2279 2472 2280
rect 2141 2281 2142 2282
rect 2277 2281 2278 2282
rect 2147 2283 2148 2284
rect 2916 2283 2917 2284
rect 2153 2285 2154 2286
rect 2295 2285 2296 2286
rect 2159 2287 2160 2288
rect 2301 2287 2302 2288
rect 2171 2289 2172 2290
rect 2313 2289 2314 2290
rect 2177 2291 2178 2292
rect 2283 2291 2284 2292
rect 2183 2293 2184 2294
rect 2307 2293 2308 2294
rect 2189 2295 2190 2296
rect 2967 2295 2968 2296
rect 2195 2297 2196 2298
rect 2771 2297 2772 2298
rect 2072 2299 2073 2300
rect 2196 2299 2197 2300
rect 1967 2301 1968 2302
rect 2073 2301 2074 2302
rect 2201 2301 2202 2302
rect 2331 2301 2332 2302
rect 2207 2303 2208 2304
rect 2355 2303 2356 2304
rect 2211 2305 2212 2306
rect 3118 2305 3119 2306
rect 2213 2307 2214 2308
rect 2265 2307 2266 2308
rect 2219 2309 2220 2310
rect 2367 2309 2368 2310
rect 2225 2311 2226 2312
rect 2253 2311 2254 2312
rect 2231 2313 2232 2314
rect 2343 2313 2344 2314
rect 2237 2315 2238 2316
rect 2511 2315 2512 2316
rect 2243 2317 2244 2318
rect 2373 2317 2374 2318
rect 2249 2319 2250 2320
rect 2711 2319 2712 2320
rect 1459 2321 1460 2322
rect 2250 2321 2251 2322
rect 1460 2323 1461 2324
rect 2168 2323 2169 2324
rect 2039 2325 2040 2326
rect 2169 2325 2170 2326
rect 2255 2325 2256 2326
rect 2391 2325 2392 2326
rect 2259 2327 2260 2328
rect 2381 2327 2382 2328
rect 2261 2329 2262 2330
rect 2397 2329 2398 2330
rect 2267 2331 2268 2332
rect 2361 2331 2362 2332
rect 2273 2333 2274 2334
rect 2415 2333 2416 2334
rect 2279 2335 2280 2336
rect 2427 2335 2428 2336
rect 2285 2337 2286 2338
rect 2421 2337 2422 2338
rect 2291 2339 2292 2340
rect 2904 2339 2905 2340
rect 2297 2341 2298 2342
rect 2403 2341 2404 2342
rect 2303 2343 2304 2344
rect 2439 2343 2440 2344
rect 2309 2345 2310 2346
rect 2451 2345 2452 2346
rect 2310 2347 2311 2348
rect 2918 2347 2919 2348
rect 2315 2349 2316 2350
rect 2433 2349 2434 2350
rect 1517 2351 1518 2352
rect 2316 2351 2317 2352
rect 2321 2351 2322 2352
rect 2457 2351 2458 2352
rect 1679 2353 1680 2354
rect 2322 2353 2323 2354
rect 2327 2353 2328 2354
rect 2385 2353 2386 2354
rect 2333 2355 2334 2356
rect 2475 2355 2476 2356
rect 2204 2357 2205 2358
rect 2334 2357 2335 2358
rect 1495 2359 1496 2360
rect 2205 2359 2206 2360
rect 2339 2359 2340 2360
rect 2481 2359 2482 2360
rect 1446 2361 1447 2362
rect 2340 2361 2341 2362
rect 2345 2361 2346 2362
rect 2469 2361 2470 2362
rect 2349 2363 2350 2364
rect 2411 2363 2412 2364
rect 2351 2365 2352 2366
rect 2487 2365 2488 2366
rect 2357 2367 2358 2368
rect 2463 2367 2464 2368
rect 2369 2369 2370 2370
rect 2499 2369 2500 2370
rect 1441 2371 1442 2372
rect 2370 2371 2371 2372
rect 2375 2371 2376 2372
rect 2505 2371 2506 2372
rect 2246 2373 2247 2374
rect 2376 2373 2377 2374
rect 2123 2375 2124 2376
rect 2247 2375 2248 2376
rect 2387 2375 2388 2376
rect 2541 2375 2542 2376
rect 2393 2377 2394 2378
rect 2529 2377 2530 2378
rect 2399 2379 2400 2380
rect 2535 2379 2536 2380
rect 2400 2381 2401 2382
rect 2492 2381 2493 2382
rect 2363 2383 2364 2384
rect 2493 2383 2494 2384
rect 2270 2385 2271 2386
rect 2364 2385 2365 2386
rect 2135 2387 2136 2388
rect 2271 2387 2272 2388
rect 2405 2387 2406 2388
rect 2523 2387 2524 2388
rect 2409 2389 2410 2390
rect 2775 2389 2776 2390
rect 2417 2391 2418 2392
rect 2553 2391 2554 2392
rect 2423 2393 2424 2394
rect 2565 2393 2566 2394
rect 2429 2395 2430 2396
rect 2571 2395 2572 2396
rect 2435 2397 2436 2398
rect 2870 2397 2871 2398
rect 2436 2399 2437 2400
rect 3114 2399 3115 2400
rect 2441 2401 2442 2402
rect 2583 2401 2584 2402
rect 2445 2403 2446 2404
rect 2840 2403 2841 2404
rect 1493 2405 1494 2406
rect 2841 2405 2842 2406
rect 2447 2407 2448 2408
rect 2589 2407 2590 2408
rect 2453 2409 2454 2410
rect 2595 2409 2596 2410
rect 2459 2411 2460 2412
rect 2607 2411 2608 2412
rect 2324 2413 2325 2414
rect 2460 2413 2461 2414
rect 2325 2415 2326 2416
rect 2823 2415 2824 2416
rect 2465 2417 2466 2418
rect 2837 2417 2838 2418
rect 2483 2419 2484 2420
rect 2613 2419 2614 2420
rect 2489 2421 2490 2422
rect 2826 2421 2827 2422
rect 2495 2423 2496 2424
rect 3015 2423 3016 2424
rect 2507 2425 2508 2426
rect 2661 2425 2662 2426
rect 2508 2427 2509 2428
rect 2663 2427 2664 2428
rect 2517 2429 2518 2430
rect 3057 2429 3058 2430
rect 2519 2431 2520 2432
rect 2673 2431 2674 2432
rect 2525 2433 2526 2434
rect 2679 2433 2680 2434
rect 2531 2435 2532 2436
rect 2691 2435 2692 2436
rect 2547 2437 2548 2438
rect 3054 2437 3055 2438
rect 2549 2439 2550 2440
rect 2709 2439 2710 2440
rect 2555 2441 2556 2442
rect 3024 2441 3025 2442
rect 2559 2443 2560 2444
rect 3128 2443 3129 2444
rect 2585 2445 2586 2446
rect 2751 2445 2752 2446
rect 2591 2447 2592 2448
rect 2769 2447 2770 2448
rect 2603 2449 2604 2450
rect 2775 2449 2776 2450
rect 2619 2451 2620 2452
rect 3064 2451 3065 2452
rect 2625 2453 2626 2454
rect 3061 2453 3062 2454
rect 2627 2455 2628 2456
rect 2793 2455 2794 2456
rect 2630 2457 2631 2458
rect 2796 2457 2797 2458
rect 2631 2459 2632 2460
rect 2900 2459 2901 2460
rect 2637 2461 2638 2462
rect 3121 2461 3122 2462
rect 2643 2463 2644 2464
rect 3107 2463 3108 2464
rect 2649 2465 2650 2466
rect 3104 2465 3105 2466
rect 2651 2467 2652 2468
rect 2823 2467 2824 2468
rect 2654 2469 2655 2470
rect 2925 2469 2926 2470
rect 2501 2471 2502 2472
rect 2655 2471 2656 2472
rect 2667 2471 2668 2472
rect 2897 2471 2898 2472
rect 2675 2473 2676 2474
rect 2835 2473 2836 2474
rect 2685 2475 2686 2476
rect 3111 2475 3112 2476
rect 2696 2477 2697 2478
rect 2886 2477 2887 2478
rect 2537 2479 2538 2480
rect 2697 2479 2698 2480
rect 2720 2479 2721 2480
rect 2898 2479 2899 2480
rect 2561 2481 2562 2482
rect 2721 2481 2722 2482
rect 2726 2481 2727 2482
rect 2904 2481 2905 2482
rect 2727 2483 2728 2484
rect 3027 2483 3028 2484
rect 2733 2485 2734 2486
rect 2867 2485 2868 2486
rect 2741 2487 2742 2488
rect 2868 2487 2869 2488
rect 2756 2489 2757 2490
rect 2946 2489 2947 2490
rect 2757 2491 2758 2492
rect 2907 2491 2908 2492
rect 2762 2493 2763 2494
rect 2952 2493 2953 2494
rect 2597 2495 2598 2496
rect 2763 2495 2764 2496
rect 2781 2495 2782 2496
rect 2970 2495 2971 2496
rect 2609 2497 2610 2498
rect 2781 2497 2782 2498
rect 2787 2497 2788 2498
rect 2982 2497 2983 2498
rect 2615 2499 2616 2500
rect 2787 2499 2788 2500
rect 2799 2499 2800 2500
rect 2988 2499 2989 2500
rect 1439 2501 1440 2502
rect 2799 2501 2800 2502
rect 2805 2501 2806 2502
rect 3125 2501 3126 2502
rect 2811 2503 2812 2504
rect 3000 2503 3001 2504
rect 2811 2505 2812 2506
rect 2964 2505 2965 2506
rect 2814 2507 2815 2508
rect 3003 2507 3004 2508
rect 2817 2509 2818 2510
rect 3006 2509 3007 2510
rect 2820 2511 2821 2512
rect 3009 2511 3010 2512
rect 2826 2513 2827 2514
rect 2928 2513 2929 2514
rect 2738 2515 2739 2516
rect 2928 2515 2929 2516
rect 2573 2517 2574 2518
rect 2739 2517 2740 2518
rect 2830 2517 2831 2518
rect 2919 2517 2920 2518
rect 2657 2519 2658 2520
rect 2829 2519 2830 2520
rect 2833 2519 2834 2520
rect 3021 2519 3022 2520
rect 2843 2521 2844 2522
rect 3030 2521 3031 2522
rect 2847 2523 2848 2524
rect 3100 2523 3101 2524
rect 2849 2525 2850 2526
rect 3036 2525 3037 2526
rect 2853 2527 2854 2528
rect 3097 2527 3098 2528
rect 2861 2529 2862 2530
rect 3048 2529 3049 2530
rect 2864 2531 2865 2532
rect 3051 2531 3052 2532
rect 2693 2533 2694 2534
rect 2865 2533 2866 2534
rect 2873 2533 2874 2534
rect 3079 2533 3080 2534
rect 2702 2535 2703 2536
rect 2874 2535 2875 2536
rect 2543 2537 2544 2538
rect 2703 2537 2704 2538
rect 2879 2537 2880 2538
rect 3076 2537 3077 2538
rect 2744 2539 2745 2540
rect 2880 2539 2881 2540
rect 2579 2541 2580 2542
rect 2745 2541 2746 2542
rect 2891 2541 2892 2542
rect 3091 2541 3092 2542
rect 2714 2543 2715 2544
rect 2892 2543 2893 2544
rect 2621 2545 2622 2546
rect 2715 2545 2716 2546
rect 2894 2545 2895 2546
rect 3094 2545 3095 2546
rect 2911 2547 2912 2548
rect 2943 2547 2944 2548
rect 2882 2549 2883 2550
rect 2910 2549 2911 2550
rect 2747 2551 2748 2552
rect 2883 2551 2884 2552
rect 2914 2551 2915 2552
rect 2940 2551 2941 2552
rect 2921 2553 2922 2554
rect 3073 2553 3074 2554
rect 2765 2555 2766 2556
rect 2922 2555 2923 2556
rect 1420 2564 1421 2565
rect 2259 2564 2260 2565
rect 1434 2566 1435 2567
rect 1604 2566 1605 2567
rect 1436 2568 1437 2569
rect 2151 2568 2152 2569
rect 1439 2570 1440 2571
rect 2319 2570 2320 2571
rect 1441 2572 1442 2573
rect 2177 2572 2178 2573
rect 1443 2574 1444 2575
rect 2307 2574 2308 2575
rect 1450 2576 1451 2577
rect 1773 2576 1774 2577
rect 1438 2578 1439 2579
rect 1450 2578 1451 2579
rect 1457 2578 1458 2579
rect 1947 2578 1948 2579
rect 1456 2580 1457 2581
rect 1641 2580 1642 2581
rect 1464 2582 1465 2583
rect 2181 2582 2182 2583
rect 1463 2584 1464 2585
rect 2322 2584 2323 2585
rect 1474 2586 1475 2587
rect 2115 2586 2116 2587
rect 1473 2588 1474 2589
rect 1863 2588 1864 2589
rect 1486 2590 1487 2591
rect 2793 2590 2794 2591
rect 1488 2592 1489 2593
rect 1923 2592 1924 2593
rect 1427 2594 1428 2595
rect 1922 2594 1923 2595
rect 1490 2596 1491 2597
rect 1839 2596 1840 2597
rect 1491 2598 1492 2599
rect 2049 2598 2050 2599
rect 1493 2600 1494 2601
rect 2858 2600 2859 2601
rect 1497 2602 1498 2603
rect 1593 2602 1594 2603
rect 1498 2604 1499 2605
rect 2048 2604 2049 2605
rect 1500 2606 1501 2607
rect 2400 2606 2401 2607
rect 1521 2608 1522 2609
rect 3114 2608 3115 2609
rect 1526 2610 1527 2611
rect 1545 2610 1546 2611
rect 1533 2612 1534 2613
rect 1538 2612 1539 2613
rect 1569 2612 1570 2613
rect 1580 2612 1581 2613
rect 1568 2614 1569 2615
rect 1575 2614 1576 2615
rect 1563 2616 1564 2617
rect 1574 2616 1575 2617
rect 1551 2618 1552 2619
rect 1562 2618 1563 2619
rect 1550 2620 1551 2621
rect 1557 2620 1558 2621
rect 1417 2622 1418 2623
rect 1556 2622 1557 2623
rect 1587 2622 1588 2623
rect 1592 2622 1593 2623
rect 1601 2622 1602 2623
rect 2984 2622 2985 2623
rect 1611 2624 1612 2625
rect 2441 2624 2442 2625
rect 1616 2626 1617 2627
rect 3164 2626 3165 2627
rect 1629 2628 1630 2629
rect 1634 2628 1635 2629
rect 1677 2628 1678 2629
rect 1766 2628 1767 2629
rect 1676 2630 1677 2631
rect 1683 2630 1684 2631
rect 1665 2632 1666 2633
rect 1682 2632 1683 2633
rect 1653 2634 1654 2635
rect 1664 2634 1665 2635
rect 1623 2636 1624 2637
rect 1652 2636 1653 2637
rect 1689 2636 1690 2637
rect 3030 2636 3031 2637
rect 1688 2638 1689 2639
rect 1719 2638 1720 2639
rect 1695 2640 1696 2641
rect 1712 2640 1713 2641
rect 1694 2642 1695 2643
rect 1725 2642 1726 2643
rect 1701 2644 1702 2645
rect 1724 2644 1725 2645
rect 1707 2646 1708 2647
rect 1730 2646 1731 2647
rect 1706 2648 1707 2649
rect 1737 2648 1738 2649
rect 1718 2650 1719 2651
rect 1749 2650 1750 2651
rect 1736 2652 1737 2653
rect 1743 2652 1744 2653
rect 1453 2654 1454 2655
rect 1742 2654 1743 2655
rect 1748 2654 1749 2655
rect 1779 2654 1780 2655
rect 1754 2656 1755 2657
rect 1785 2656 1786 2657
rect 1761 2658 1762 2659
rect 2990 2658 2991 2659
rect 1671 2660 1672 2661
rect 1760 2660 1761 2661
rect 1659 2662 1660 2663
rect 1670 2662 1671 2663
rect 1647 2664 1648 2665
rect 1658 2664 1659 2665
rect 1772 2664 1773 2665
rect 1833 2664 1834 2665
rect 1784 2666 1785 2667
rect 1845 2666 1846 2667
rect 1797 2668 1798 2669
rect 2912 2668 2913 2669
rect 1796 2670 1797 2671
rect 1857 2670 1858 2671
rect 1832 2672 1833 2673
rect 1851 2672 1852 2673
rect 1838 2674 1839 2675
rect 1875 2674 1876 2675
rect 1844 2676 1845 2677
rect 1971 2676 1972 2677
rect 1850 2678 1851 2679
rect 1881 2678 1882 2679
rect 1856 2680 1857 2681
rect 1899 2680 1900 2681
rect 1862 2682 1863 2683
rect 1977 2682 1978 2683
rect 1880 2684 1881 2685
rect 1893 2684 1894 2685
rect 1887 2686 1888 2687
rect 3155 2686 3156 2687
rect 1886 2688 1887 2689
rect 1929 2688 1930 2689
rect 1424 2690 1425 2691
rect 1928 2690 1929 2691
rect 1892 2692 1893 2693
rect 1905 2692 1906 2693
rect 1898 2694 1899 2695
rect 1935 2694 1936 2695
rect 1904 2696 1905 2697
rect 1941 2696 1942 2697
rect 1911 2698 1912 2699
rect 2964 2698 2965 2699
rect 1910 2700 1911 2701
rect 1953 2700 1954 2701
rect 1916 2702 1917 2703
rect 1959 2702 1960 2703
rect 1934 2704 1935 2705
rect 1965 2704 1966 2705
rect 1940 2706 1941 2707
rect 3027 2706 3028 2707
rect 1946 2708 1947 2709
rect 1995 2708 1996 2709
rect 1952 2710 1953 2711
rect 1983 2710 1984 2711
rect 1958 2712 1959 2713
rect 1989 2712 1990 2713
rect 1964 2714 1965 2715
rect 3024 2714 3025 2715
rect 1970 2716 1971 2717
rect 3015 2716 3016 2717
rect 1976 2718 1977 2719
rect 2007 2718 2008 2719
rect 1982 2720 1983 2721
rect 2001 2720 2002 2721
rect 1988 2722 1989 2723
rect 3107 2722 3108 2723
rect 1994 2724 1995 2725
rect 2031 2724 2032 2725
rect 2000 2726 2001 2727
rect 2025 2726 2026 2727
rect 2006 2728 2007 2729
rect 2037 2728 2038 2729
rect 2019 2730 2020 2731
rect 2792 2730 2793 2731
rect 2018 2732 2019 2733
rect 2043 2732 2044 2733
rect 2024 2734 2025 2735
rect 2055 2734 2056 2735
rect 2030 2736 2031 2737
rect 2085 2736 2086 2737
rect 2036 2738 2037 2739
rect 2067 2738 2068 2739
rect 2042 2740 2043 2741
rect 2079 2740 2080 2741
rect 1483 2742 1484 2743
rect 2078 2742 2079 2743
rect 1446 2744 1447 2745
rect 1482 2744 1483 2745
rect 2054 2744 2055 2745
rect 3226 2744 3227 2745
rect 2061 2746 2062 2747
rect 2930 2746 2931 2747
rect 2060 2748 2061 2749
rect 2073 2748 2074 2749
rect 1432 2750 1433 2751
rect 2072 2750 2073 2751
rect 1431 2752 1432 2753
rect 1599 2752 1600 2753
rect 1598 2754 1599 2755
rect 2943 2754 2944 2755
rect 2084 2756 2085 2757
rect 2103 2756 2104 2757
rect 2097 2758 2098 2759
rect 2102 2758 2103 2759
rect 2091 2760 2092 2761
rect 2096 2760 2097 2761
rect 2090 2762 2091 2763
rect 2109 2762 2110 2763
rect 1471 2764 1472 2765
rect 2108 2764 2109 2765
rect 1470 2766 1471 2767
rect 2066 2766 2067 2767
rect 2114 2766 2115 2767
rect 2121 2766 2122 2767
rect 2120 2768 2121 2769
rect 2127 2768 2128 2769
rect 1495 2770 1496 2771
rect 2126 2770 2127 2771
rect 2150 2770 2151 2771
rect 2157 2770 2158 2771
rect 2156 2772 2157 2773
rect 2163 2772 2164 2773
rect 2162 2774 2163 2775
rect 2205 2774 2206 2775
rect 2180 2776 2181 2777
rect 2199 2776 2200 2777
rect 2187 2778 2188 2779
rect 2222 2778 2223 2779
rect 2186 2780 2187 2781
rect 3152 2780 3153 2781
rect 2196 2782 2197 2783
rect 2231 2782 2232 2783
rect 2198 2784 2199 2785
rect 2217 2784 2218 2785
rect 2204 2786 2205 2787
rect 2253 2786 2254 2787
rect 2216 2788 2217 2789
rect 3185 2788 3186 2789
rect 2229 2790 2230 2791
rect 2258 2790 2259 2791
rect 2193 2792 2194 2793
rect 2228 2792 2229 2793
rect 2192 2794 2193 2795
rect 3107 2794 3108 2795
rect 2241 2796 2242 2797
rect 2967 2796 2968 2797
rect 2240 2798 2241 2799
rect 2553 2798 2554 2799
rect 2250 2800 2251 2801
rect 2285 2800 2286 2801
rect 2252 2802 2253 2803
rect 2547 2802 2548 2803
rect 2271 2804 2272 2805
rect 2306 2804 2307 2805
rect 2270 2806 2271 2807
rect 2577 2806 2578 2807
rect 2295 2808 2296 2809
rect 2318 2808 2319 2809
rect 2294 2810 2295 2811
rect 2325 2810 2326 2811
rect 2301 2812 2302 2813
rect 2324 2812 2325 2813
rect 2316 2814 2317 2815
rect 2351 2814 2352 2815
rect 2364 2814 2365 2815
rect 2876 2814 2877 2815
rect 2334 2816 2335 2817
rect 2363 2816 2364 2817
rect 2310 2818 2311 2819
rect 2333 2818 2334 2819
rect 2370 2818 2371 2819
rect 2405 2818 2406 2819
rect 2376 2820 2377 2821
rect 2387 2820 2388 2821
rect 2340 2822 2341 2823
rect 2375 2822 2376 2823
rect 2436 2822 2437 2823
rect 2495 2822 2496 2823
rect 2451 2824 2452 2825
rect 2919 2824 2920 2825
rect 2409 2826 2410 2827
rect 2450 2826 2451 2827
rect 2403 2828 2404 2829
rect 2408 2828 2409 2829
rect 2367 2830 2368 2831
rect 2402 2830 2403 2831
rect 2460 2830 2461 2831
rect 2501 2830 2502 2831
rect 2493 2832 2494 2833
rect 2552 2832 2553 2833
rect 2433 2834 2434 2835
rect 2492 2834 2493 2835
rect 1429 2836 1430 2837
rect 2432 2836 2433 2837
rect 2499 2836 2500 2837
rect 2546 2836 2547 2837
rect 2457 2838 2458 2839
rect 2498 2838 2499 2839
rect 2415 2840 2416 2841
rect 2456 2840 2457 2841
rect 2379 2842 2380 2843
rect 2414 2842 2415 2843
rect 2378 2844 2379 2845
rect 2385 2844 2386 2845
rect 2373 2846 2374 2847
rect 2384 2846 2385 2847
rect 2337 2848 2338 2849
rect 2372 2848 2373 2849
rect 2289 2850 2290 2851
rect 2336 2850 2337 2851
rect 2529 2850 2530 2851
rect 2576 2850 2577 2851
rect 2481 2852 2482 2853
rect 2528 2852 2529 2853
rect 2439 2854 2440 2855
rect 2480 2854 2481 2855
rect 2397 2856 2398 2857
rect 2438 2856 2439 2857
rect 2361 2858 2362 2859
rect 2396 2858 2397 2859
rect 2331 2860 2332 2861
rect 2360 2860 2361 2861
rect 2283 2862 2284 2863
rect 2330 2862 2331 2863
rect 2247 2864 2248 2865
rect 2282 2864 2283 2865
rect 2246 2866 2247 2867
rect 2517 2866 2518 2867
rect 2475 2868 2476 2869
rect 2516 2868 2517 2869
rect 2474 2870 2475 2871
rect 2916 2870 2917 2871
rect 2613 2872 2614 2873
rect 3061 2872 3062 2873
rect 2601 2874 2602 2875
rect 2612 2874 2613 2875
rect 2571 2876 2572 2877
rect 2600 2876 2601 2877
rect 2523 2878 2524 2879
rect 2570 2878 2571 2879
rect 1586 2880 1587 2881
rect 2522 2880 2523 2881
rect 2655 2880 2656 2881
rect 3229 2880 3230 2881
rect 2595 2882 2596 2883
rect 2654 2882 2655 2883
rect 2594 2884 2595 2885
rect 3189 2884 3190 2885
rect 2745 2886 2746 2887
rect 2816 2886 2817 2887
rect 2691 2888 2692 2889
rect 2744 2888 2745 2889
rect 2631 2890 2632 2891
rect 2690 2890 2691 2891
rect 2787 2890 2788 2891
rect 3240 2890 3241 2891
rect 2721 2892 2722 2893
rect 2786 2892 2787 2893
rect 2667 2894 2668 2895
rect 2720 2894 2721 2895
rect 2666 2896 2667 2897
rect 3064 2896 3065 2897
rect 2796 2898 2797 2899
rect 2888 2898 2889 2899
rect 2805 2900 2806 2901
rect 2936 2900 2937 2901
rect 2739 2902 2740 2903
rect 2804 2902 2805 2903
rect 2685 2904 2686 2905
rect 2738 2904 2739 2905
rect 2211 2906 2212 2907
rect 2684 2906 2685 2907
rect 2210 2908 2211 2909
rect 2349 2908 2350 2909
rect 2313 2910 2314 2911
rect 2348 2910 2349 2911
rect 2277 2912 2278 2913
rect 2312 2912 2313 2913
rect 2276 2914 2277 2915
rect 2511 2914 2512 2915
rect 2487 2916 2488 2917
rect 2510 2916 2511 2917
rect 2445 2918 2446 2919
rect 2486 2918 2487 2919
rect 1692 2920 1693 2921
rect 2444 2920 2445 2921
rect 2811 2920 2812 2921
rect 2942 2920 2943 2921
rect 1505 2922 1506 2923
rect 2810 2922 2811 2923
rect 2826 2922 2827 2923
rect 2906 2922 2907 2923
rect 2829 2924 2830 2925
rect 2918 2924 2919 2925
rect 2763 2926 2764 2927
rect 2828 2926 2829 2927
rect 2762 2928 2763 2929
rect 3247 2928 3248 2929
rect 2835 2930 2836 2931
rect 3026 2930 3027 2931
rect 2757 2932 2758 2933
rect 2834 2932 2835 2933
rect 2697 2934 2698 2935
rect 2756 2934 2757 2935
rect 2643 2936 2644 2937
rect 2696 2936 2697 2937
rect 2642 2938 2643 2939
rect 3233 2938 3234 2939
rect 2841 2940 2842 2941
rect 3097 2940 3098 2941
rect 2775 2942 2776 2943
rect 2840 2942 2841 2943
rect 2709 2944 2710 2945
rect 2774 2944 2775 2945
rect 2637 2946 2638 2947
rect 2708 2946 2709 2947
rect 2636 2948 2637 2949
rect 2894 2948 2895 2949
rect 2847 2950 2848 2951
rect 2954 2950 2955 2951
rect 2781 2952 2782 2953
rect 2846 2952 2847 2953
rect 2727 2954 2728 2955
rect 2780 2954 2781 2955
rect 2673 2956 2674 2957
rect 2726 2956 2727 2957
rect 2619 2958 2620 2959
rect 2672 2958 2673 2959
rect 2618 2960 2619 2961
rect 3219 2960 3220 2961
rect 2853 2962 2854 2963
rect 2948 2962 2949 2963
rect 2769 2964 2770 2965
rect 2852 2964 2853 2965
rect 2703 2966 2704 2967
rect 2768 2966 2769 2967
rect 2649 2968 2650 2969
rect 2702 2968 2703 2969
rect 2589 2970 2590 2971
rect 2648 2970 2649 2971
rect 2588 2972 2589 2973
rect 3192 2972 3193 2973
rect 2865 2974 2866 2975
rect 2960 2974 2961 2975
rect 2799 2976 2800 2977
rect 2864 2976 2865 2977
rect 2733 2978 2734 2979
rect 2798 2978 2799 2979
rect 2133 2980 2134 2981
rect 2732 2980 2733 2981
rect 2132 2982 2133 2983
rect 2139 2982 2140 2983
rect 2138 2984 2139 2985
rect 2169 2984 2170 2985
rect 1467 2986 1468 2987
rect 2168 2986 2169 2987
rect 1466 2988 1467 2989
rect 1640 2988 1641 2989
rect 2868 2988 2869 2989
rect 2966 2988 2967 2989
rect 2870 2990 2871 2991
rect 3222 2990 3223 2991
rect 2883 2992 2884 2993
rect 3059 2992 3060 2993
rect 2886 2994 2887 2995
rect 3032 2994 3033 2995
rect 2898 2996 2899 2997
rect 3014 2996 3015 2997
rect 2910 2998 2911 2999
rect 3057 2998 3058 2999
rect 2823 3000 2824 3001
rect 2909 3000 2910 3001
rect 2751 3002 2752 3003
rect 2822 3002 2823 3003
rect 2679 3004 2680 3005
rect 2750 3004 2751 3005
rect 2625 3006 2626 3007
rect 2678 3006 2679 3007
rect 2583 3008 2584 3009
rect 2624 3008 2625 3009
rect 2535 3010 2536 3011
rect 2582 3010 2583 3011
rect 2534 3012 2535 3013
rect 2897 3012 2898 3013
rect 2880 3014 2881 3015
rect 3056 3014 3057 3015
rect 1803 3016 1804 3017
rect 2879 3016 2880 3017
rect 1802 3018 1803 3019
rect 1815 3018 1816 3019
rect 1502 3020 1503 3021
rect 1814 3020 1815 3021
rect 2924 3020 2925 3021
rect 3125 3020 3126 3021
rect 2928 3022 2929 3023
rect 3071 3022 3072 3023
rect 2940 3024 2941 3025
rect 3068 3024 3069 3025
rect 2946 3026 2947 3027
rect 3086 3026 3087 3027
rect 2963 3028 2964 3029
rect 3118 3028 3119 3029
rect 2972 3030 2973 3031
rect 3100 3030 3101 3031
rect 2996 3032 2997 3033
rect 3243 3032 3244 3033
rect 3000 3034 3001 3035
rect 3140 3034 3141 3035
rect 3003 3036 3004 3037
rect 3143 3036 3144 3037
rect 2508 3038 2509 3039
rect 3002 3038 3003 3039
rect 3006 3038 3007 3039
rect 3146 3038 3147 3039
rect 1791 3040 1792 3041
rect 3005 3040 3006 3041
rect 1790 3042 1791 3043
rect 1809 3042 1810 3043
rect 1808 3044 1809 3045
rect 1821 3044 1822 3045
rect 1820 3046 1821 3047
rect 1827 3046 1828 3047
rect 1826 3048 1827 3049
rect 1869 3048 1870 3049
rect 1868 3050 1869 3051
rect 2013 3050 2014 3051
rect 2012 3052 2013 3053
rect 3012 3052 3013 3053
rect 3009 3054 3010 3055
rect 3149 3054 3150 3055
rect 2892 3056 2893 3057
rect 3008 3056 3009 3057
rect 2715 3058 2716 3059
rect 2891 3058 2892 3059
rect 2661 3060 2662 3061
rect 2714 3060 2715 3061
rect 2607 3062 2608 3063
rect 2660 3062 2661 3063
rect 2559 3064 2560 3065
rect 2606 3064 2607 3065
rect 2558 3066 2559 3067
rect 2565 3066 2566 3067
rect 2541 3068 2542 3069
rect 2564 3068 2565 3069
rect 2463 3070 2464 3071
rect 2540 3070 2541 3071
rect 2421 3072 2422 3073
rect 2462 3072 2463 3073
rect 1589 3074 1590 3075
rect 2420 3074 2421 3075
rect 3018 3074 3019 3075
rect 3158 3074 3159 3075
rect 3021 3076 3022 3077
rect 3161 3076 3162 3077
rect 2904 3078 2905 3079
rect 3020 3078 3021 3079
rect 3036 3078 3037 3079
rect 3179 3078 3180 3079
rect 3044 3080 3045 3081
rect 3167 3080 3168 3081
rect 3048 3082 3049 3083
rect 3054 3082 3055 3083
rect 3051 3084 3052 3085
rect 3176 3084 3177 3085
rect 2874 3086 2875 3087
rect 3050 3086 3051 3087
rect 3073 3086 3074 3087
rect 3213 3086 3214 3087
rect 2366 3088 2367 3089
rect 3074 3088 3075 3089
rect 3076 3088 3077 3089
rect 3216 3088 3217 3089
rect 2300 3090 2301 3091
rect 3077 3090 3078 3091
rect 3079 3090 3080 3091
rect 3111 3090 3112 3091
rect 2922 3092 2923 3093
rect 3080 3092 3081 3093
rect 2970 3094 2971 3095
rect 3110 3094 3111 3095
rect 3091 3096 3092 3097
rect 3201 3096 3202 3097
rect 2952 3098 2953 3099
rect 3092 3098 3093 3099
rect 3094 3098 3095 3099
rect 3204 3098 3205 3099
rect 3104 3100 3105 3101
rect 3182 3100 3183 3101
rect 2505 3102 2506 3103
rect 3104 3102 3105 3103
rect 2469 3104 2470 3105
rect 2504 3104 2505 3105
rect 2427 3106 2428 3107
rect 2468 3106 2469 3107
rect 2391 3108 2392 3109
rect 2426 3108 2427 3109
rect 2355 3110 2356 3111
rect 2390 3110 2391 3111
rect 2343 3112 2344 3113
rect 2354 3112 2355 3113
rect 2265 3114 2266 3115
rect 2342 3114 2343 3115
rect 2235 3116 2236 3117
rect 2264 3116 2265 3117
rect 1460 3118 1461 3119
rect 2234 3118 2235 3119
rect 1459 3120 1460 3121
rect 2288 3120 2289 3121
rect 3121 3120 3122 3121
rect 3236 3120 3237 3121
rect 2982 3122 2983 3123
rect 3122 3122 3123 3123
rect 3128 3122 3129 3123
rect 3250 3122 3251 3123
rect 2988 3124 2989 3125
rect 3128 3124 3129 3125
rect 1417 3133 1418 3134
rect 1922 3133 1923 3134
rect 1420 3135 1421 3136
rect 2048 3135 2049 3136
rect 1427 3137 1428 3138
rect 1916 3137 1917 3138
rect 1431 3139 1432 3140
rect 2387 3139 2388 3140
rect 1431 3141 1432 3142
rect 2156 3141 2157 3142
rect 1441 3143 1442 3144
rect 2302 3143 2303 3144
rect 1459 3145 1460 3146
rect 1946 3145 1947 3146
rect 1463 3147 1464 3148
rect 1688 3147 1689 3148
rect 1427 3149 1428 3150
rect 1687 3149 1688 3150
rect 1450 3151 1451 3152
rect 1462 3151 1463 3152
rect 1438 3153 1439 3154
rect 1450 3153 1451 3154
rect 1438 3155 1439 3156
rect 2612 3155 2613 3156
rect 1466 3157 1467 3158
rect 1904 3157 1905 3158
rect 1468 3159 1469 3160
rect 3037 3159 3038 3160
rect 1473 3161 1474 3162
rect 2060 3161 2061 3162
rect 1485 3163 1486 3164
rect 2282 3163 2283 3164
rect 1488 3165 1489 3166
rect 2222 3165 2223 3166
rect 1491 3167 1492 3168
rect 2114 3167 2115 3168
rect 1495 3169 1496 3170
rect 2042 3169 2043 3170
rect 1482 3171 1483 3172
rect 1494 3171 1495 3172
rect 1498 3171 1499 3172
rect 2036 3171 2037 3172
rect 1502 3173 1503 3174
rect 2072 3173 2073 3174
rect 1505 3175 1506 3176
rect 2012 3175 2013 3176
rect 1507 3177 1508 3178
rect 1568 3177 1569 3178
rect 1514 3179 1515 3180
rect 1519 3179 1520 3180
rect 1526 3179 1527 3180
rect 1531 3179 1532 3180
rect 1525 3181 1526 3182
rect 1616 3181 1617 3182
rect 1528 3183 1529 3184
rect 2501 3183 2502 3184
rect 1538 3185 1539 3186
rect 1543 3185 1544 3186
rect 1562 3185 1563 3186
rect 1567 3185 1568 3186
rect 1556 3187 1557 3188
rect 1561 3187 1562 3188
rect 1478 3189 1479 3190
rect 1555 3189 1556 3190
rect 1586 3189 1587 3190
rect 2024 3189 2025 3190
rect 1580 3191 1581 3192
rect 1585 3191 1586 3192
rect 1574 3193 1575 3194
rect 1579 3193 1580 3194
rect 1475 3195 1476 3196
rect 1573 3195 1574 3196
rect 1592 3195 1593 3196
rect 1615 3195 1616 3196
rect 1601 3197 1602 3198
rect 1604 3197 1605 3198
rect 1434 3199 1435 3200
rect 1603 3199 1604 3200
rect 1434 3201 1435 3202
rect 1612 3201 1613 3202
rect 1609 3203 1610 3204
rect 3044 3203 3045 3204
rect 1658 3205 1659 3206
rect 3074 3205 3075 3206
rect 1652 3207 1653 3208
rect 1657 3207 1658 3208
rect 1694 3207 1695 3208
rect 1699 3207 1700 3208
rect 1712 3207 1713 3208
rect 3243 3207 3244 3208
rect 1706 3209 1707 3210
rect 1711 3209 1712 3210
rect 1724 3209 1725 3210
rect 2422 3209 2423 3210
rect 1723 3211 1724 3212
rect 3247 3211 3248 3212
rect 1748 3213 1749 3214
rect 1777 3213 1778 3214
rect 1736 3215 1737 3216
rect 1747 3215 1748 3216
rect 1844 3215 1845 3216
rect 1921 3215 1922 3216
rect 1802 3217 1803 3218
rect 1843 3217 1844 3218
rect 1772 3219 1773 3220
rect 1801 3219 1802 3220
rect 1742 3221 1743 3222
rect 1771 3221 1772 3222
rect 1730 3223 1731 3224
rect 1741 3223 1742 3224
rect 1424 3225 1425 3226
rect 1729 3225 1730 3226
rect 1424 3227 1425 3228
rect 1693 3227 1694 3228
rect 1862 3227 1863 3228
rect 3152 3227 3153 3228
rect 1820 3229 1821 3230
rect 1861 3229 1862 3230
rect 1819 3231 1820 3232
rect 1826 3231 1827 3232
rect 1825 3233 1826 3234
rect 1832 3233 1833 3234
rect 1796 3235 1797 3236
rect 1831 3235 1832 3236
rect 1795 3237 1796 3238
rect 1850 3237 1851 3238
rect 1790 3239 1791 3240
rect 1849 3239 1850 3240
rect 1789 3241 1790 3242
rect 1808 3241 1809 3242
rect 1807 3243 1808 3244
rect 1838 3243 1839 3244
rect 1837 3245 1838 3246
rect 1856 3245 1857 3246
rect 1873 3245 1874 3246
rect 1880 3245 1881 3246
rect 1879 3247 1880 3248
rect 1892 3247 1893 3248
rect 1868 3249 1869 3250
rect 1891 3249 1892 3250
rect 1814 3251 1815 3252
rect 1867 3251 1868 3252
rect 1784 3253 1785 3254
rect 1813 3253 1814 3254
rect 1903 3253 1904 3254
rect 1928 3253 1929 3254
rect 1915 3255 1916 3256
rect 2792 3255 2793 3256
rect 1927 3257 1928 3258
rect 1952 3257 1953 3258
rect 1621 3259 1622 3260
rect 1951 3259 1952 3260
rect 1945 3261 1946 3262
rect 1976 3261 1977 3262
rect 1975 3263 1976 3264
rect 2000 3263 2001 3264
rect 1999 3265 2000 3266
rect 2030 3265 2031 3266
rect 1482 3267 1483 3268
rect 2029 3267 2030 3268
rect 2011 3269 2012 3270
rect 2066 3269 2067 3270
rect 2023 3271 2024 3272
rect 2090 3271 2091 3272
rect 2035 3273 2036 3274
rect 2096 3273 2097 3274
rect 2041 3275 2042 3276
rect 2102 3275 2103 3276
rect 2047 3277 2048 3278
rect 2078 3277 2079 3278
rect 2054 3279 2055 3280
rect 2065 3279 2066 3280
rect 2053 3281 2054 3282
rect 2108 3281 2109 3282
rect 2059 3283 2060 3284
rect 2120 3283 2121 3284
rect 2071 3285 2072 3286
rect 2138 3285 2139 3286
rect 2080 3287 2081 3288
rect 2879 3287 2880 3288
rect 2089 3289 2090 3290
rect 2150 3289 2151 3290
rect 2095 3291 2096 3292
rect 2180 3291 2181 3292
rect 2101 3293 2102 3294
rect 2186 3293 2187 3294
rect 2107 3295 2108 3296
rect 2174 3295 2175 3296
rect 2113 3297 2114 3298
rect 2162 3297 2163 3298
rect 1598 3299 1599 3300
rect 2161 3299 2162 3300
rect 1510 3301 1511 3302
rect 1597 3301 1598 3302
rect 2119 3301 2120 3302
rect 2666 3301 2667 3302
rect 2132 3303 2133 3304
rect 3155 3303 3156 3304
rect 2131 3305 2132 3306
rect 2210 3305 2211 3306
rect 2137 3307 2138 3308
rect 2270 3307 2271 3308
rect 2149 3309 2150 3310
rect 2216 3309 2217 3310
rect 2155 3311 2156 3312
rect 2252 3311 2253 3312
rect 2173 3313 2174 3314
rect 2228 3313 2229 3314
rect 1456 3315 1457 3316
rect 2227 3315 2228 3316
rect 1456 3317 1457 3318
rect 2177 3317 2178 3318
rect 2176 3319 2177 3320
rect 2231 3319 2232 3320
rect 2179 3321 2180 3322
rect 2234 3321 2235 3322
rect 2185 3323 2186 3324
rect 2588 3323 2589 3324
rect 2194 3325 2195 3326
rect 2285 3325 2286 3326
rect 2204 3327 2205 3328
rect 3136 3327 3137 3328
rect 2203 3329 2204 3330
rect 2264 3329 2265 3330
rect 2206 3331 2207 3332
rect 2351 3331 2352 3332
rect 2209 3333 2210 3334
rect 2258 3333 2259 3334
rect 2215 3335 2216 3336
rect 2600 3335 2601 3336
rect 2221 3337 2222 3338
rect 2564 3337 2565 3338
rect 2233 3339 2234 3340
rect 2288 3339 2289 3340
rect 2240 3341 2241 3342
rect 3189 3341 3190 3342
rect 2239 3343 2240 3344
rect 2660 3343 2661 3344
rect 2198 3345 2199 3346
rect 2659 3345 2660 3346
rect 2197 3347 2198 3348
rect 2594 3347 2595 3348
rect 2251 3349 2252 3350
rect 2342 3349 2343 3350
rect 2257 3351 2258 3352
rect 2300 3351 2301 3352
rect 1441 3353 1442 3354
rect 2299 3353 2300 3354
rect 2263 3355 2264 3356
rect 2366 3355 2367 3356
rect 2269 3357 2270 3358
rect 2306 3357 2307 3358
rect 2276 3359 2277 3360
rect 3077 3359 3078 3360
rect 1886 3361 1887 3362
rect 3076 3361 3077 3362
rect 1885 3363 1886 3364
rect 1898 3363 1899 3364
rect 1897 3365 1898 3366
rect 1910 3365 1911 3366
rect 1909 3367 1910 3368
rect 1934 3367 1935 3368
rect 1933 3369 1934 3370
rect 1958 3369 1959 3370
rect 1957 3371 1958 3372
rect 1982 3371 1983 3372
rect 1589 3373 1590 3374
rect 1981 3373 1982 3374
rect 2275 3373 2276 3374
rect 2312 3373 2313 3374
rect 2281 3375 2282 3376
rect 2330 3375 2331 3376
rect 2284 3377 2285 3378
rect 2333 3377 2334 3378
rect 2287 3379 2288 3380
rect 2336 3379 2337 3380
rect 2305 3381 2306 3382
rect 2534 3381 2535 3382
rect 2311 3383 2312 3384
rect 2897 3383 2898 3384
rect 2324 3385 2325 3386
rect 2329 3385 2330 3386
rect 2192 3387 2193 3388
rect 2323 3387 2324 3388
rect 1417 3389 1418 3390
rect 2191 3389 2192 3390
rect 2335 3389 2336 3390
rect 2546 3389 2547 3390
rect 2341 3391 2342 3392
rect 2384 3391 2385 3392
rect 2354 3393 2355 3394
rect 2662 3393 2663 3394
rect 2353 3395 2354 3396
rect 2474 3395 2475 3396
rect 2365 3397 2366 3398
rect 2498 3397 2499 3398
rect 2375 3399 2376 3400
rect 2410 3399 2411 3400
rect 2363 3401 2364 3402
rect 2374 3401 2375 3402
rect 2383 3401 2384 3402
rect 2690 3401 2691 3402
rect 2396 3403 2397 3404
rect 2894 3403 2895 3404
rect 2395 3405 2396 3406
rect 2480 3405 2481 3406
rect 2434 3407 2435 3408
rect 2495 3407 2496 3408
rect 2441 3409 2442 3410
rect 2446 3409 2447 3410
rect 2405 3411 2406 3412
rect 2440 3411 2441 3412
rect 1550 3413 1551 3414
rect 2404 3413 2405 3414
rect 2468 3413 2469 3414
rect 2497 3413 2498 3414
rect 2432 3415 2433 3416
rect 2467 3415 2468 3416
rect 2420 3417 2421 3418
rect 2431 3417 2432 3418
rect 2414 3419 2415 3420
rect 2419 3419 2420 3420
rect 2413 3421 2414 3422
rect 2510 3421 2511 3422
rect 2470 3423 2471 3424
rect 2876 3423 2877 3424
rect 2473 3425 2474 3426
rect 2570 3425 2571 3426
rect 2479 3427 2480 3428
rect 2696 3427 2697 3428
rect 2126 3429 2127 3430
rect 2695 3429 2696 3430
rect 2125 3431 2126 3432
rect 2672 3431 2673 3432
rect 2504 3433 2505 3434
rect 3185 3433 3186 3434
rect 2486 3435 2487 3436
rect 2503 3435 2504 3436
rect 2450 3437 2451 3438
rect 2485 3437 2486 3438
rect 2444 3439 2445 3440
rect 2449 3439 2450 3440
rect 2438 3441 2439 3442
rect 2443 3441 2444 3442
rect 2402 3443 2403 3444
rect 2437 3443 2438 3444
rect 1500 3445 1501 3446
rect 2401 3445 2402 3446
rect 2509 3445 2510 3446
rect 3182 3445 3183 3446
rect 2528 3447 2529 3448
rect 2545 3447 2546 3448
rect 2527 3449 2528 3450
rect 2654 3449 2655 3450
rect 2533 3451 2534 3452
rect 2576 3451 2577 3452
rect 2552 3453 2553 3454
rect 3104 3453 3105 3454
rect 2551 3455 2552 3456
rect 2582 3455 2583 3456
rect 2558 3457 2559 3458
rect 3192 3457 3193 3458
rect 2557 3459 2558 3460
rect 3107 3459 3108 3460
rect 2563 3461 2564 3462
rect 2606 3461 2607 3462
rect 2569 3463 2570 3464
rect 3198 3463 3199 3464
rect 2575 3465 2576 3466
rect 3195 3465 3196 3466
rect 2581 3467 2582 3468
rect 2648 3467 2649 3468
rect 2587 3469 2588 3470
rect 2624 3469 2625 3470
rect 2599 3471 2600 3472
rect 2963 3471 2964 3472
rect 2605 3473 2606 3474
rect 2636 3473 2637 3474
rect 2611 3475 2612 3476
rect 2642 3475 2643 3476
rect 2623 3477 2624 3478
rect 3236 3477 3237 3478
rect 2629 3479 2630 3480
rect 3240 3479 3241 3480
rect 2635 3481 2636 3482
rect 2714 3481 2715 3482
rect 2647 3483 2648 3484
rect 2720 3483 2721 3484
rect 2653 3485 2654 3486
rect 2726 3485 2727 3486
rect 2665 3487 2666 3488
rect 3118 3487 3119 3488
rect 2671 3489 2672 3490
rect 2738 3489 2739 3490
rect 1970 3491 1971 3492
rect 2737 3491 2738 3492
rect 1420 3493 1421 3494
rect 1969 3493 1970 3494
rect 2684 3493 2685 3494
rect 3115 3493 3116 3494
rect 1503 3495 1504 3496
rect 2683 3495 2684 3496
rect 2689 3495 2690 3496
rect 2744 3495 2745 3496
rect 2708 3497 2709 3498
rect 3226 3497 3227 3498
rect 2707 3499 2708 3500
rect 3250 3499 3251 3500
rect 2713 3501 2714 3502
rect 2756 3501 2757 3502
rect 2719 3503 2720 3504
rect 2750 3503 2751 3504
rect 2725 3505 2726 3506
rect 2768 3505 2769 3506
rect 2743 3507 2744 3508
rect 2798 3507 2799 3508
rect 2749 3509 2750 3510
rect 2804 3509 2805 3510
rect 2755 3511 2756 3512
rect 3188 3511 3189 3512
rect 2767 3513 2768 3514
rect 3229 3513 3230 3514
rect 2774 3515 2775 3516
rect 3170 3515 3171 3516
rect 2773 3517 2774 3518
rect 2828 3517 2829 3518
rect 1940 3519 1941 3520
rect 2827 3519 2828 3520
rect 1624 3521 1625 3522
rect 1939 3521 1940 3522
rect 2791 3521 2792 3522
rect 2822 3521 2823 3522
rect 2797 3523 2798 3524
rect 2834 3523 2835 3524
rect 2803 3525 2804 3526
rect 3219 3525 3220 3526
rect 2641 3527 2642 3528
rect 3219 3527 3220 3528
rect 2821 3529 2822 3530
rect 2846 3529 2847 3530
rect 2833 3531 2834 3532
rect 2912 3531 2913 3532
rect 2845 3533 2846 3534
rect 2864 3533 2865 3534
rect 2852 3535 2853 3536
rect 2863 3535 2864 3536
rect 2870 3535 2871 3536
rect 2884 3535 2885 3536
rect 2869 3537 2870 3538
rect 3152 3537 3153 3538
rect 2875 3539 2876 3540
rect 2924 3539 2925 3540
rect 2881 3541 2882 3542
rect 2891 3541 2892 3542
rect 2888 3543 2889 3544
rect 3073 3543 3074 3544
rect 2887 3545 2888 3546
rect 2930 3545 2931 3546
rect 2893 3547 2894 3548
rect 2936 3547 2937 3548
rect 2911 3549 2912 3550
rect 2942 3549 2943 3550
rect 2918 3551 2919 3552
rect 3155 3551 3156 3552
rect 2917 3553 2918 3554
rect 2972 3553 2973 3554
rect 2923 3555 2924 3556
rect 3005 3555 3006 3556
rect 2935 3557 2936 3558
rect 2966 3557 2967 3558
rect 1470 3559 1471 3560
rect 2965 3559 2966 3560
rect 1471 3561 1472 3562
rect 2348 3561 2349 3562
rect 2347 3563 2348 3564
rect 2408 3563 2409 3564
rect 2372 3565 2373 3566
rect 2407 3565 2408 3566
rect 2360 3567 2361 3568
rect 2371 3567 2372 3568
rect 2359 3569 2360 3570
rect 2492 3569 2493 3570
rect 2491 3571 2492 3572
rect 2618 3571 2619 3572
rect 2617 3573 2618 3574
rect 2702 3573 2703 3574
rect 2701 3575 2702 3576
rect 2762 3575 2763 3576
rect 2761 3577 2762 3578
rect 3191 3577 3192 3578
rect 2944 3579 2945 3580
rect 2960 3579 2961 3580
rect 2948 3581 2949 3582
rect 3052 3581 3053 3582
rect 2947 3583 2948 3584
rect 2984 3583 2985 3584
rect 2971 3585 2972 3586
rect 3008 3585 3009 3586
rect 2977 3587 2978 3588
rect 3014 3587 3015 3588
rect 2983 3589 2984 3590
rect 3020 3589 3021 3590
rect 3002 3591 3003 3592
rect 3040 3591 3041 3592
rect 3001 3593 3002 3594
rect 3026 3593 3027 3594
rect 3013 3595 3014 3596
rect 3164 3595 3165 3596
rect 3019 3597 3020 3598
rect 3056 3597 3057 3598
rect 3022 3599 3023 3600
rect 3059 3599 3060 3600
rect 3034 3601 3035 3602
rect 3071 3601 3072 3602
rect 3043 3603 3044 3604
rect 3080 3603 3081 3604
rect 3050 3605 3051 3606
rect 3167 3605 3168 3606
rect 2144 3607 2145 3608
rect 3049 3607 3050 3608
rect 2143 3609 2144 3610
rect 2246 3609 2247 3610
rect 2245 3611 2246 3612
rect 2294 3611 2295 3612
rect 2293 3613 2294 3614
rect 2378 3613 2379 3614
rect 2377 3615 2378 3616
rect 2426 3615 2427 3616
rect 2390 3617 2391 3618
rect 2425 3617 2426 3618
rect 2389 3619 2390 3620
rect 3133 3619 3134 3620
rect 3055 3621 3056 3622
rect 3086 3621 3087 3622
rect 3061 3623 3062 3624
rect 3092 3623 3093 3624
rect 3079 3625 3080 3626
rect 3110 3625 3111 3626
rect 3091 3627 3092 3628
rect 3122 3627 3123 3628
rect 3097 3629 3098 3630
rect 3143 3629 3144 3630
rect 2996 3631 2997 3632
rect 3142 3631 3143 3632
rect 2995 3633 2996 3634
rect 3032 3633 3033 3634
rect 3031 3635 3032 3636
rect 3068 3635 3069 3636
rect 3109 3635 3110 3636
rect 3146 3635 3147 3636
rect 2786 3637 2787 3638
rect 3145 3637 3146 3638
rect 2785 3639 2786 3640
rect 2816 3639 2817 3640
rect 1964 3641 1965 3642
rect 2815 3641 2816 3642
rect 1963 3643 1964 3644
rect 1988 3643 1989 3644
rect 1987 3645 1988 3646
rect 1994 3645 1995 3646
rect 1993 3647 1994 3648
rect 2006 3647 2007 3648
rect 2005 3649 2006 3650
rect 2018 3649 2019 3650
rect 2017 3651 2018 3652
rect 2084 3651 2085 3652
rect 2083 3653 2084 3654
rect 2168 3653 2169 3654
rect 2167 3655 2168 3656
rect 2678 3655 2679 3656
rect 2677 3657 2678 3658
rect 3209 3657 3210 3658
rect 3112 3659 3113 3660
rect 3149 3659 3150 3660
rect 3121 3661 3122 3662
rect 3158 3661 3159 3662
rect 3124 3663 3125 3664
rect 3161 3663 3162 3664
rect 3128 3665 3129 3666
rect 3222 3665 3223 3666
rect 3127 3667 3128 3668
rect 3173 3667 3174 3668
rect 3130 3669 3131 3670
rect 3140 3669 3141 3670
rect 3139 3671 3140 3672
rect 3179 3671 3180 3672
rect 3164 3673 3165 3674
rect 3201 3673 3202 3674
rect 2318 3675 2319 3676
rect 3202 3675 3203 3676
rect 2317 3677 2318 3678
rect 2540 3677 2541 3678
rect 2522 3679 2523 3680
rect 2539 3679 2540 3680
rect 2516 3681 2517 3682
rect 2521 3681 2522 3682
rect 2515 3683 2516 3684
rect 3148 3683 3149 3684
rect 3167 3683 3168 3684
rect 3204 3683 3205 3684
rect 2593 3685 2594 3686
rect 3205 3685 3206 3686
rect 3176 3687 3177 3688
rect 3233 3687 3234 3688
rect 3182 3689 3183 3690
rect 3213 3689 3214 3690
rect 2941 3691 2942 3692
rect 3212 3691 3213 3692
rect 3185 3693 3186 3694
rect 3216 3693 3217 3694
rect 2954 3695 2955 3696
rect 3216 3695 3217 3696
rect 2953 3697 2954 3698
rect 2990 3697 2991 3698
rect 1417 3706 1418 3707
rect 1927 3706 1928 3707
rect 1434 3708 1435 3709
rect 2089 3708 2090 3709
rect 1434 3710 1435 3711
rect 1585 3710 1586 3711
rect 1438 3712 1439 3713
rect 1519 3712 1520 3713
rect 1438 3714 1439 3715
rect 1573 3714 1574 3715
rect 1468 3716 1469 3717
rect 2209 3716 2210 3717
rect 1475 3718 1476 3719
rect 2194 3718 2195 3719
rect 1478 3720 1479 3721
rect 1531 3720 1532 3721
rect 1485 3722 1486 3723
rect 1813 3722 1814 3723
rect 1468 3724 1469 3725
rect 1814 3724 1815 3725
rect 1485 3726 1486 3727
rect 2737 3726 2738 3727
rect 1503 3728 1504 3729
rect 1909 3728 1910 3729
rect 1503 3730 1504 3731
rect 1843 3730 1844 3731
rect 1507 3732 1508 3733
rect 1574 3732 1575 3733
rect 1507 3734 1508 3735
rect 1615 3734 1616 3735
rect 1510 3736 1511 3737
rect 3227 3736 3228 3737
rect 1514 3738 1515 3739
rect 3221 3738 3222 3739
rect 1517 3740 1518 3741
rect 2173 3740 2174 3741
rect 1528 3742 1529 3743
rect 3112 3742 3113 3743
rect 1592 3744 1593 3745
rect 1597 3744 1598 3745
rect 1598 3746 1599 3747
rect 1765 3746 1766 3747
rect 1612 3748 1613 3749
rect 2149 3748 2150 3749
rect 1624 3750 1625 3751
rect 2665 3750 2666 3751
rect 1628 3752 1629 3753
rect 1663 3752 1664 3753
rect 1424 3754 1425 3755
rect 1664 3754 1665 3755
rect 1417 3756 1418 3757
rect 1424 3756 1425 3757
rect 1633 3756 1634 3757
rect 2003 3756 2004 3757
rect 1652 3758 1653 3759
rect 2434 3758 2435 3759
rect 1675 3760 1676 3761
rect 3198 3760 3199 3761
rect 1706 3762 1707 3763
rect 1879 3762 1880 3763
rect 1717 3764 1718 3765
rect 1784 3764 1785 3765
rect 1669 3766 1670 3767
rect 1718 3766 1719 3767
rect 1670 3768 1671 3769
rect 1687 3768 1688 3769
rect 1688 3770 1689 3771
rect 1693 3770 1694 3771
rect 1529 3772 1530 3773
rect 1694 3772 1695 3773
rect 1736 3772 1737 3773
rect 1771 3772 1772 3773
rect 1482 3774 1483 3775
rect 1772 3774 1773 3775
rect 1482 3776 1483 3777
rect 2143 3776 2144 3777
rect 1844 3778 1845 3779
rect 1969 3778 1970 3779
rect 1856 3780 1857 3781
rect 1939 3780 1940 3781
rect 1871 3782 1872 3783
rect 2176 3782 2177 3783
rect 1880 3784 1881 3785
rect 1981 3784 1982 3785
rect 1910 3786 1911 3787
rect 2041 3786 2042 3787
rect 1928 3788 1929 3789
rect 2107 3788 2108 3789
rect 1940 3790 1941 3791
rect 2083 3790 2084 3791
rect 1961 3792 1962 3793
rect 2206 3792 2207 3793
rect 1970 3794 1971 3795
rect 2047 3794 2048 3795
rect 1982 3796 1983 3797
rect 2227 3796 2228 3797
rect 1609 3798 1610 3799
rect 2228 3798 2229 3799
rect 1510 3800 1511 3801
rect 1610 3800 1611 3801
rect 2027 3800 2028 3801
rect 2302 3800 2303 3801
rect 2042 3802 2043 3803
rect 2269 3802 2270 3803
rect 2051 3804 2052 3805
rect 2284 3804 2285 3805
rect 2063 3806 2064 3807
rect 2410 3806 2411 3807
rect 2078 3808 2079 3809
rect 2287 3808 2288 3809
rect 2084 3810 2085 3811
rect 2341 3810 2342 3811
rect 2090 3812 2091 3813
rect 2437 3812 2438 3813
rect 2099 3814 2100 3815
rect 2440 3814 2441 3815
rect 2105 3816 2106 3817
rect 2404 3816 2405 3817
rect 2108 3818 2109 3819
rect 2251 3818 2252 3819
rect 2059 3820 2060 3821
rect 2252 3820 2253 3821
rect 2060 3822 2061 3823
rect 2407 3822 2408 3823
rect 2137 3824 2138 3825
rect 3216 3824 3217 3825
rect 2138 3826 2139 3827
rect 2353 3826 2354 3827
rect 2144 3828 2145 3829
rect 2461 3828 2462 3829
rect 2150 3830 2151 3831
rect 2443 3830 2444 3831
rect 2174 3832 2175 3833
rect 2503 3832 2504 3833
rect 2197 3834 2198 3835
rect 2408 3834 2409 3835
rect 1500 3836 1501 3837
rect 2198 3836 2199 3837
rect 2210 3836 2211 3837
rect 2365 3836 2366 3837
rect 2131 3838 2132 3839
rect 2366 3838 2367 3839
rect 2132 3840 2133 3841
rect 2347 3840 2348 3841
rect 2215 3842 2216 3843
rect 3252 3842 3253 3843
rect 2216 3844 2217 3845
rect 2521 3844 2522 3845
rect 2101 3846 2102 3847
rect 2522 3846 2523 3847
rect 2102 3848 2103 3849
rect 2401 3848 2402 3849
rect 2185 3850 2186 3851
rect 2402 3850 2403 3851
rect 2186 3852 2187 3853
rect 2359 3852 2360 3853
rect 2257 3854 2258 3855
rect 2342 3854 2343 3855
rect 2258 3856 2259 3857
rect 2515 3856 2516 3857
rect 2167 3858 2168 3859
rect 2516 3858 2517 3859
rect 2168 3860 2169 3861
rect 2455 3860 2456 3861
rect 2263 3862 2264 3863
rect 3291 3862 3292 3863
rect 2161 3864 2162 3865
rect 2264 3864 2265 3865
rect 2162 3866 2163 3867
rect 2497 3866 2498 3867
rect 2239 3868 2240 3869
rect 2498 3868 2499 3869
rect 2240 3870 2241 3871
rect 2539 3870 2540 3871
rect 2270 3872 2271 3873
rect 2662 3872 2663 3873
rect 2288 3874 2289 3875
rect 2293 3874 2294 3875
rect 2294 3876 2295 3877
rect 2533 3876 2534 3877
rect 2317 3878 2318 3879
rect 2360 3878 2361 3879
rect 2318 3880 2319 3881
rect 2389 3880 2390 3881
rect 2348 3882 2349 3883
rect 2569 3882 2570 3883
rect 2354 3884 2355 3885
rect 2575 3884 2576 3885
rect 2390 3886 2391 3887
rect 2605 3886 2606 3887
rect 2323 3888 2324 3889
rect 2606 3888 2607 3889
rect 2324 3890 2325 3891
rect 2473 3890 2474 3891
rect 1999 3892 2000 3893
rect 2474 3892 2475 3893
rect 2000 3894 2001 3895
rect 2191 3894 2192 3895
rect 2192 3896 2193 3897
rect 2395 3896 2396 3897
rect 2396 3898 2397 3899
rect 2611 3898 2612 3899
rect 2422 3900 2423 3901
rect 2612 3900 2613 3901
rect 2438 3902 2439 3903
rect 2623 3902 2624 3903
rect 2444 3904 2445 3905
rect 2557 3904 2558 3905
rect 1993 3906 1994 3907
rect 2558 3906 2559 3907
rect 2446 3908 2447 3909
rect 2927 3908 2928 3909
rect 2456 3910 2457 3911
rect 3288 3910 3289 3911
rect 2462 3912 2463 3913
rect 3202 3912 3203 3913
rect 2479 3914 2480 3915
rect 2534 3914 2535 3915
rect 2119 3916 2120 3917
rect 2480 3916 2481 3917
rect 2120 3918 2121 3919
rect 2431 3918 2432 3919
rect 2432 3920 2433 3921
rect 2581 3920 2582 3921
rect 2485 3922 2486 3923
rect 3231 3922 3232 3923
rect 2125 3924 2126 3925
rect 2486 3924 2487 3925
rect 2126 3926 2127 3927
rect 2467 3926 2468 3927
rect 2468 3928 2469 3929
rect 2527 3928 2528 3929
rect 2504 3930 2505 3931
rect 2641 3930 2642 3931
rect 2509 3932 2510 3933
rect 3205 3932 3206 3933
rect 2510 3934 2511 3935
rect 3267 3934 3268 3935
rect 2528 3936 2529 3937
rect 3073 3936 3074 3937
rect 2540 3938 2541 3939
rect 2617 3938 2618 3939
rect 1849 3940 1850 3941
rect 2618 3940 2619 3941
rect 1621 3942 1622 3943
rect 1850 3942 1851 3943
rect 2563 3942 2564 3943
rect 3195 3942 3196 3943
rect 2383 3944 2384 3945
rect 2564 3944 2565 3945
rect 2155 3946 2156 3947
rect 2384 3946 2385 3947
rect 2156 3948 2157 3949
rect 2377 3948 2378 3949
rect 2005 3950 2006 3951
rect 2378 3950 2379 3951
rect 2006 3952 2007 3953
rect 2281 3952 2282 3953
rect 2282 3954 2283 3955
rect 2335 3954 2336 3955
rect 2336 3956 2337 3957
rect 2593 3956 2594 3957
rect 2570 3958 2571 3959
rect 2635 3958 2636 3959
rect 1753 3960 1754 3961
rect 2636 3960 2637 3961
rect 1478 3962 1479 3963
rect 1754 3962 1755 3963
rect 2576 3962 2577 3963
rect 2647 3962 2648 3963
rect 2582 3964 2583 3965
rect 2671 3964 2672 3965
rect 2594 3966 2595 3967
rect 3305 3966 3306 3967
rect 2624 3968 2625 3969
rect 2701 3968 2702 3969
rect 2642 3970 2643 3971
rect 2713 3970 2714 3971
rect 2659 3972 2660 3973
rect 2897 3972 2898 3973
rect 2660 3974 2661 3975
rect 3170 3974 3171 3975
rect 2666 3976 2667 3977
rect 3118 3976 3119 3977
rect 2672 3978 2673 3979
rect 2731 3978 2732 3979
rect 2683 3980 2684 3981
rect 3302 3980 3303 3981
rect 2684 3982 2685 3983
rect 2749 3982 2750 3983
rect 2689 3984 2690 3985
rect 3212 3984 3213 3985
rect 2690 3986 2691 3987
rect 2755 3986 2756 3987
rect 2695 3988 2696 3989
rect 3115 3988 3116 3989
rect 2696 3990 2697 3991
rect 2761 3990 2762 3991
rect 2702 3992 2703 3993
rect 2767 3992 2768 3993
rect 2714 3994 2715 3995
rect 3188 3994 3189 3995
rect 2725 3996 2726 3997
rect 3173 3996 3174 3997
rect 1861 3998 1862 3999
rect 2726 3998 2727 3999
rect 1862 4000 1863 4001
rect 2017 4000 2018 4001
rect 2018 4002 2019 4003
rect 2329 4002 2330 4003
rect 1987 4004 1988 4005
rect 2330 4004 2331 4005
rect 1988 4006 1989 4007
rect 2233 4006 2234 4007
rect 2234 4008 2235 4009
rect 3234 4008 3235 4009
rect 2732 4010 2733 4011
rect 2803 4010 2804 4011
rect 2743 4012 2744 4013
rect 3284 4012 3285 4013
rect 2744 4014 2745 4015
rect 2791 4014 2792 4015
rect 2750 4016 2751 4017
rect 2797 4016 2798 4017
rect 2756 4018 2757 4019
rect 2809 4018 2810 4019
rect 2762 4020 2763 4021
rect 2815 4020 2816 4021
rect 1807 4022 1808 4023
rect 2816 4022 2817 4023
rect 1808 4024 1809 4025
rect 1867 4024 1868 4025
rect 1868 4026 1869 4027
rect 2023 4026 2024 4027
rect 2024 4028 2025 4029
rect 2299 4028 2300 4029
rect 2300 4030 2301 4031
rect 2551 4030 2552 4031
rect 2065 4032 2066 4033
rect 2552 4032 2553 4033
rect 1475 4034 1476 4035
rect 2066 4034 2067 4035
rect 2768 4034 2769 4035
rect 2821 4034 2822 4035
rect 1795 4036 1796 4037
rect 2822 4036 2823 4037
rect 1796 4038 1797 4039
rect 1903 4038 1904 4039
rect 1500 4040 1501 4041
rect 1904 4040 1905 4041
rect 2779 4040 2780 4041
rect 3191 4040 3192 4041
rect 1825 4042 1826 4043
rect 2780 4042 2781 4043
rect 1826 4044 1827 4045
rect 1945 4044 1946 4045
rect 1946 4046 1947 4047
rect 2095 4046 2096 4047
rect 2096 4048 2097 4049
rect 2425 4048 2426 4049
rect 2426 4050 2427 4051
rect 2599 4050 2600 4051
rect 2600 4052 2601 4053
rect 2677 4052 2678 4053
rect 2678 4054 2679 4055
rect 3281 4054 3282 4055
rect 2792 4056 2793 4057
rect 2845 4056 2846 4057
rect 1709 4058 1710 4059
rect 2846 4058 2847 4059
rect 2798 4060 2799 4061
rect 3249 4060 3250 4061
rect 2804 4062 2805 4063
rect 2857 4062 2858 4063
rect 2080 4064 2081 4065
rect 2858 4064 2859 4065
rect 2081 4066 2082 4067
rect 2374 4066 2375 4067
rect 2810 4066 2811 4067
rect 2863 4066 2864 4067
rect 1747 4068 1748 4069
rect 2864 4068 2865 4069
rect 1748 4070 1749 4071
rect 1837 4070 1838 4071
rect 1838 4072 1839 4073
rect 1957 4072 1958 4073
rect 1958 4074 1959 4075
rect 2203 4074 2204 4075
rect 2204 4076 2205 4077
rect 2413 4076 2414 4077
rect 2113 4078 2114 4079
rect 2414 4078 2415 4079
rect 2114 4080 2115 4081
rect 2419 4080 2420 4081
rect 2420 4082 2421 4083
rect 2587 4082 2588 4083
rect 2588 4084 2589 4085
rect 2653 4084 2654 4085
rect 2654 4086 2655 4087
rect 2719 4086 2720 4087
rect 2720 4088 2721 4089
rect 2785 4088 2786 4089
rect 1921 4090 1922 4091
rect 2786 4090 2787 4091
rect 1922 4092 1923 4093
rect 2071 4092 2072 4093
rect 2053 4094 2054 4095
rect 2072 4094 2073 4095
rect 2054 4096 2055 4097
rect 2371 4096 2372 4097
rect 2221 4098 2222 4099
rect 2372 4098 2373 4099
rect 2222 4100 2223 4101
rect 3298 4100 3299 4101
rect 2839 4102 2840 4103
rect 3274 4102 3275 4103
rect 1741 4104 1742 4105
rect 2840 4104 2841 4105
rect 1742 4106 1743 4107
rect 1777 4106 1778 4107
rect 1723 4108 1724 4109
rect 1778 4108 1779 4109
rect 1724 4110 1725 4111
rect 1801 4110 1802 4111
rect 1802 4112 1803 4113
rect 1897 4112 1898 4113
rect 1891 4114 1892 4115
rect 1898 4114 1899 4115
rect 1892 4116 1893 4117
rect 2011 4116 2012 4117
rect 2012 4118 2013 4119
rect 2275 4118 2276 4119
rect 2276 4120 2277 4121
rect 2311 4120 2312 4121
rect 2245 4122 2246 4123
rect 2312 4122 2313 4123
rect 2246 4124 2247 4125
rect 2545 4124 2546 4125
rect 2029 4126 2030 4127
rect 2546 4126 2547 4127
rect 2852 4126 2853 4127
rect 2881 4126 2882 4127
rect 2855 4128 2856 4129
rect 3133 4128 3134 4129
rect 2869 4130 2870 4131
rect 2882 4130 2883 4131
rect 2875 4132 2876 4133
rect 3155 4132 3156 4133
rect 2876 4134 2877 4135
rect 2905 4134 2906 4135
rect 2879 4136 2880 4137
rect 2908 4136 2909 4137
rect 2884 4138 2885 4139
rect 3277 4138 3278 4139
rect 2900 4140 2901 4141
rect 3270 4140 3271 4141
rect 2906 4142 2907 4143
rect 3215 4142 3216 4143
rect 2917 4144 2918 4145
rect 2990 4144 2991 4145
rect 2918 4146 2919 4147
rect 3052 4146 3053 4147
rect 2923 4148 2924 4149
rect 3076 4148 3077 4149
rect 1601 4150 1602 4151
rect 2924 4150 2925 4151
rect 2941 4150 2942 4151
rect 2969 4150 2970 4151
rect 1525 4152 1526 4153
rect 2942 4152 2943 4153
rect 1526 4154 1527 4155
rect 1657 4154 1658 4155
rect 1427 4156 1428 4157
rect 1658 4156 1659 4157
rect 1427 4158 1428 4159
rect 2843 4158 2844 4159
rect 2971 4158 2972 4159
rect 3026 4158 3027 4159
rect 2893 4160 2894 4161
rect 2972 4160 2973 4161
rect 1759 4162 1760 4163
rect 2894 4162 2895 4163
rect 1760 4164 1761 4165
rect 1831 4164 1832 4165
rect 1681 4166 1682 4167
rect 1832 4166 1833 4167
rect 1682 4168 1683 4169
rect 1711 4168 1712 4169
rect 1699 4170 1700 4171
rect 1712 4170 1713 4171
rect 1700 4172 1701 4173
rect 1729 4172 1730 4173
rect 1730 4174 1731 4175
rect 1819 4174 1820 4175
rect 1820 4176 1821 4177
rect 1933 4176 1934 4177
rect 1934 4178 1935 4179
rect 3158 4178 3159 4179
rect 3001 4180 3002 4181
rect 3068 4180 3069 4181
rect 2947 4182 2948 4183
rect 3002 4182 3003 4183
rect 2944 4184 2945 4185
rect 2948 4184 2949 4185
rect 2470 4186 2471 4187
rect 2945 4186 2946 4187
rect 3008 4186 3009 4187
rect 3219 4186 3220 4187
rect 3019 4188 3020 4189
rect 3104 4188 3105 4189
rect 3020 4190 3021 4191
rect 3295 4190 3296 4191
rect 3022 4192 3023 4193
rect 3107 4192 3108 4193
rect 3031 4194 3032 4195
rect 3101 4194 3102 4195
rect 2977 4196 2978 4197
rect 3032 4196 3033 4197
rect 2911 4198 2912 4199
rect 2978 4198 2979 4199
rect 2912 4200 2913 4201
rect 3136 4200 3137 4201
rect 3034 4202 3035 4203
rect 3086 4202 3087 4203
rect 3040 4204 3041 4205
rect 3113 4204 3114 4205
rect 3043 4206 3044 4207
rect 3134 4206 3135 4207
rect 3044 4208 3045 4209
rect 3142 4208 3143 4209
rect 2648 4210 2649 4211
rect 3143 4210 3144 4211
rect 3049 4212 3050 4213
rect 3145 4212 3146 4213
rect 2965 4214 2966 4215
rect 3050 4214 3051 4215
rect 2966 4216 2967 4217
rect 3209 4216 3210 4217
rect 3055 4218 3056 4219
rect 3146 4218 3147 4219
rect 3061 4220 3062 4221
rect 3203 4220 3204 4221
rect 2995 4222 2996 4223
rect 3062 4222 3063 4223
rect 2887 4224 2888 4225
rect 2996 4224 2997 4225
rect 1915 4226 1916 4227
rect 2888 4226 2889 4227
rect 1431 4228 1432 4229
rect 1916 4228 1917 4229
rect 1431 4230 1432 4231
rect 1586 4230 1587 4231
rect 3091 4230 3092 4231
rect 3176 4230 3177 4231
rect 3109 4232 3110 4233
rect 3197 4232 3198 4233
rect 3037 4234 3038 4235
rect 3110 4234 3111 4235
rect 2983 4236 2984 4237
rect 3038 4236 3039 4237
rect 2935 4238 2936 4239
rect 2984 4238 2985 4239
rect 2936 4240 2937 4241
rect 3148 4240 3149 4241
rect 3121 4242 3122 4243
rect 3200 4242 3201 4243
rect 3122 4244 3123 4245
rect 3224 4244 3225 4245
rect 3124 4246 3125 4247
rect 3161 4246 3162 4247
rect 3127 4248 3128 4249
rect 3206 4248 3207 4249
rect 1420 4250 1421 4251
rect 3128 4250 3129 4251
rect 1420 4252 1421 4253
rect 1994 4252 1995 4253
rect 3130 4252 3131 4253
rect 3209 4252 3210 4253
rect 3139 4254 3140 4255
rect 3218 4254 3219 4255
rect 2305 4256 2306 4257
rect 3140 4256 3141 4257
rect 1963 4258 1964 4259
rect 2306 4258 2307 4259
rect 1964 4260 1965 4261
rect 2035 4260 2036 4261
rect 1471 4262 1472 4263
rect 2036 4262 2037 4263
rect 1471 4264 1472 4265
rect 2030 4264 2031 4265
rect 3152 4264 3153 4265
rect 3194 4264 3195 4265
rect 3164 4266 3165 4267
rect 3243 4266 3244 4267
rect 3079 4268 3080 4269
rect 3164 4268 3165 4269
rect 3013 4270 3014 4271
rect 3080 4270 3081 4271
rect 2953 4272 2954 4273
rect 3014 4272 3015 4273
rect 2833 4274 2834 4275
rect 2954 4274 2955 4275
rect 1789 4276 1790 4277
rect 2834 4276 2835 4277
rect 1790 4278 1791 4279
rect 1885 4278 1886 4279
rect 1886 4280 1887 4281
rect 1951 4280 1952 4281
rect 1441 4282 1442 4283
rect 1952 4282 1953 4283
rect 1441 4284 1442 4285
rect 2048 4284 2049 4285
rect 3167 4284 3168 4285
rect 3246 4284 3247 4285
rect 3182 4286 3183 4287
rect 3261 4286 3262 4287
rect 3097 4288 3098 4289
rect 3182 4288 3183 4289
rect 3098 4290 3099 4291
rect 3212 4290 3213 4291
rect 3185 4292 3186 4293
rect 3264 4292 3265 4293
rect 1431 4301 1432 4302
rect 1580 4301 1581 4302
rect 1441 4303 1442 4304
rect 1550 4303 1551 4304
rect 1441 4305 1442 4306
rect 2024 4305 2025 4306
rect 1468 4307 1469 4308
rect 2042 4307 2043 4308
rect 1468 4309 1469 4310
rect 2006 4309 2007 4310
rect 1503 4311 1504 4312
rect 1910 4311 1911 4312
rect 1510 4313 1511 4314
rect 1622 4313 1623 4314
rect 1510 4315 1511 4316
rect 1922 4315 1923 4316
rect 1517 4317 1518 4318
rect 3311 4317 3312 4318
rect 1517 4319 1518 4320
rect 1940 4319 1941 4320
rect 1526 4321 1527 4322
rect 1652 4321 1653 4322
rect 1485 4323 1486 4324
rect 1526 4323 1527 4324
rect 1485 4325 1486 4326
rect 2000 4325 2001 4326
rect 1541 4327 1542 4328
rect 2828 4327 2829 4328
rect 1586 4329 1587 4330
rect 1616 4329 1617 4330
rect 1601 4331 1602 4332
rect 3243 4331 3244 4332
rect 1610 4333 1611 4334
rect 1634 4333 1635 4334
rect 1434 4335 1435 4336
rect 1610 4335 1611 4336
rect 1628 4335 1629 4336
rect 1652 4335 1653 4336
rect 1507 4337 1508 4338
rect 1628 4337 1629 4338
rect 1507 4339 1508 4340
rect 1838 4339 1839 4340
rect 1500 4341 1501 4342
rect 1838 4341 1839 4342
rect 1500 4343 1501 4344
rect 1778 4343 1779 4344
rect 1640 4345 1641 4346
rect 1676 4345 1677 4346
rect 1604 4347 1605 4348
rect 1640 4347 1641 4348
rect 1661 4347 1662 4348
rect 3032 4347 3033 4348
rect 1709 4349 1710 4350
rect 2858 4349 2859 4350
rect 1514 4351 1515 4352
rect 2858 4351 2859 4352
rect 1478 4353 1479 4354
rect 1514 4353 1515 4354
rect 1778 4353 1779 4354
rect 2864 4353 2865 4354
rect 1856 4355 1857 4356
rect 2000 4355 2001 4356
rect 1434 4357 1435 4358
rect 1856 4357 1857 4358
rect 1868 4357 1869 4358
rect 2042 4357 2043 4358
rect 1754 4359 1755 4360
rect 1868 4359 1869 4360
rect 1424 4361 1425 4362
rect 1754 4361 1755 4362
rect 1424 4363 1425 4364
rect 1742 4363 1743 4364
rect 1712 4365 1713 4366
rect 1742 4365 1743 4366
rect 1712 4367 1713 4368
rect 1832 4367 1833 4368
rect 1832 4369 1833 4370
rect 2846 4369 2847 4370
rect 1871 4371 1872 4372
rect 2045 4371 2046 4372
rect 1880 4373 1881 4374
rect 2024 4373 2025 4374
rect 1772 4375 1773 4376
rect 1880 4375 1881 4376
rect 1682 4377 1683 4378
rect 1772 4377 1773 4378
rect 1886 4377 1887 4378
rect 2006 4377 2007 4378
rect 1886 4379 1887 4380
rect 2834 4379 2835 4380
rect 1898 4381 1899 4382
rect 1922 4381 1923 4382
rect 1898 4383 1899 4384
rect 2822 4383 2823 4384
rect 1940 4385 1941 4386
rect 3300 4385 3301 4386
rect 1961 4387 1962 4388
rect 2147 4387 2148 4388
rect 2003 4389 2004 4390
rect 2159 4389 2160 4390
rect 2027 4391 2028 4392
rect 2231 4391 2232 4392
rect 2051 4393 2052 4394
rect 2273 4393 2274 4394
rect 2063 4395 2064 4396
rect 2291 4395 2292 4396
rect 2081 4397 2082 4398
rect 2279 4397 2280 4398
rect 2099 4399 2100 4400
rect 2321 4399 2322 4400
rect 2105 4401 2106 4402
rect 2327 4401 2328 4402
rect 2216 4403 2217 4404
rect 3234 4403 3235 4404
rect 2216 4405 2217 4406
rect 2474 4405 2475 4406
rect 2246 4407 2247 4408
rect 2474 4407 2475 4408
rect 2288 4409 2289 4410
rect 3143 4409 3144 4410
rect 2060 4411 2061 4412
rect 2288 4411 2289 4412
rect 1892 4413 1893 4414
rect 2060 4413 2061 4414
rect 1748 4415 1749 4416
rect 1892 4415 1893 4416
rect 1748 4417 1749 4418
rect 1784 4417 1785 4418
rect 1784 4419 1785 4420
rect 2612 4419 2613 4420
rect 2357 4421 2358 4422
rect 2897 4421 2898 4422
rect 2402 4423 2403 4424
rect 3370 4423 3371 4424
rect 2192 4425 2193 4426
rect 2402 4425 2403 4426
rect 2108 4427 2109 4428
rect 2192 4427 2193 4428
rect 2429 4427 2430 4428
rect 2843 4427 2844 4428
rect 2438 4429 2439 4430
rect 2612 4429 2613 4430
rect 2438 4431 2439 4432
rect 2546 4431 2547 4432
rect 2354 4433 2355 4434
rect 2546 4433 2547 4434
rect 2186 4435 2187 4436
rect 2354 4435 2355 4436
rect 2186 4437 2187 4438
rect 2558 4437 2559 4438
rect 2384 4439 2385 4440
rect 2558 4439 2559 4440
rect 2162 4441 2163 4442
rect 2384 4441 2385 4442
rect 2162 4443 2163 4444
rect 2252 4443 2253 4444
rect 2252 4445 2253 4446
rect 2270 4445 2271 4446
rect 2048 4447 2049 4448
rect 2270 4447 2271 4448
rect 2048 4449 2049 4450
rect 2306 4449 2307 4450
rect 2138 4451 2139 4452
rect 2306 4451 2307 4452
rect 1976 4453 1977 4454
rect 2138 4453 2139 4454
rect 1478 4455 1479 4456
rect 1976 4455 1977 4456
rect 2450 4455 2451 4456
rect 3395 4455 3396 4456
rect 2222 4457 2223 4458
rect 2450 4457 2451 4458
rect 2018 4459 2019 4460
rect 2222 4459 2223 4460
rect 1874 4461 1875 4462
rect 2018 4461 2019 4462
rect 1760 4463 1761 4464
rect 1874 4463 1875 4464
rect 1503 4465 1504 4466
rect 1760 4465 1761 4466
rect 2504 4465 2505 4466
rect 3367 4465 3368 4466
rect 2294 4467 2295 4468
rect 2504 4467 2505 4468
rect 1427 4469 1428 4470
rect 2294 4469 2295 4470
rect 1427 4471 1428 4472
rect 2108 4471 2109 4472
rect 2594 4471 2595 4472
rect 2738 4471 2739 4472
rect 2426 4473 2427 4474
rect 2594 4473 2595 4474
rect 2210 4475 2211 4476
rect 2426 4475 2427 4476
rect 2078 4477 2079 4478
rect 2210 4477 2211 4478
rect 1904 4479 1905 4480
rect 2078 4479 2079 4480
rect 1808 4481 1809 4482
rect 1904 4481 1905 4482
rect 1420 4483 1421 4484
rect 1808 4483 1809 4484
rect 1420 4485 1421 4486
rect 2246 4485 2247 4486
rect 2684 4485 2685 4486
rect 3281 4485 3282 4486
rect 2534 4487 2535 4488
rect 2684 4487 2685 4488
rect 2414 4489 2415 4490
rect 2534 4489 2535 4490
rect 2414 4491 2415 4492
rect 3326 4491 3327 4492
rect 2690 4493 2691 4494
rect 2828 4493 2829 4494
rect 2540 4495 2541 4496
rect 2690 4495 2691 4496
rect 2348 4497 2349 4498
rect 2540 4497 2541 4498
rect 2126 4499 2127 4500
rect 2348 4499 2349 4500
rect 1970 4501 1971 4502
rect 2126 4501 2127 4502
rect 1820 4503 1821 4504
rect 1970 4503 1971 4504
rect 1820 4505 1821 4506
rect 2924 4505 2925 4506
rect 2696 4507 2697 4508
rect 2834 4507 2835 4508
rect 2696 4509 2697 4510
rect 2726 4509 2727 4510
rect 2582 4511 2583 4512
rect 2726 4511 2727 4512
rect 2390 4513 2391 4514
rect 2582 4513 2583 4514
rect 1417 4515 1418 4516
rect 2390 4515 2391 4516
rect 1417 4517 1418 4518
rect 1482 4517 1483 4518
rect 1482 4519 1483 4520
rect 1994 4519 1995 4520
rect 1850 4521 1851 4522
rect 1994 4521 1995 4522
rect 1475 4523 1476 4524
rect 1850 4523 1851 4524
rect 2708 4523 2709 4524
rect 3023 4523 3024 4524
rect 2570 4525 2571 4526
rect 2708 4525 2709 4526
rect 2408 4527 2409 4528
rect 2570 4527 2571 4528
rect 2198 4529 2199 4530
rect 2408 4529 2409 4530
rect 2030 4531 2031 4532
rect 2198 4531 2199 4532
rect 2030 4533 2031 4534
rect 2456 4533 2457 4534
rect 2456 4535 2457 4536
rect 3398 4535 3399 4536
rect 2714 4537 2715 4538
rect 3333 4537 3334 4538
rect 2576 4539 2577 4540
rect 2714 4539 2715 4540
rect 2480 4541 2481 4542
rect 2576 4541 2577 4542
rect 2282 4543 2283 4544
rect 2480 4543 2481 4544
rect 1438 4545 1439 4546
rect 2282 4545 2283 4546
rect 2786 4545 2787 4546
rect 2924 4545 2925 4546
rect 2648 4547 2649 4548
rect 2786 4547 2787 4548
rect 2516 4549 2517 4550
rect 2648 4549 2649 4550
rect 2324 4551 2325 4552
rect 2516 4551 2517 4552
rect 2102 4553 2103 4554
rect 2324 4553 2325 4554
rect 1964 4555 1965 4556
rect 2102 4555 2103 4556
rect 1538 4557 1539 4558
rect 1964 4557 1965 4558
rect 2792 4557 2793 4558
rect 2930 4557 2931 4558
rect 2654 4559 2655 4560
rect 2792 4559 2793 4560
rect 2492 4561 2493 4562
rect 2654 4561 2655 4562
rect 2342 4563 2343 4564
rect 2492 4563 2493 4564
rect 2120 4565 2121 4566
rect 2342 4565 2343 4566
rect 1946 4567 1947 4568
rect 2120 4567 2121 4568
rect 1946 4569 1947 4570
rect 3252 4569 3253 4570
rect 2822 4571 2823 4572
rect 3284 4571 3285 4572
rect 2840 4573 2841 4574
rect 3374 4573 3375 4574
rect 2702 4575 2703 4576
rect 2840 4575 2841 4576
rect 2564 4577 2565 4578
rect 2702 4577 2703 4578
rect 2522 4579 2523 4580
rect 2564 4579 2565 4580
rect 2372 4581 2373 4582
rect 2522 4581 2523 4582
rect 2180 4583 2181 4584
rect 2372 4583 2373 4584
rect 2180 4585 2181 4586
rect 2264 4585 2265 4586
rect 2084 4587 2085 4588
rect 2264 4587 2265 4588
rect 1928 4589 1929 4590
rect 2084 4589 2085 4590
rect 1814 4591 1815 4592
rect 1928 4591 1929 4592
rect 1814 4593 1815 4594
rect 2636 4593 2637 4594
rect 2486 4595 2487 4596
rect 2636 4595 2637 4596
rect 2360 4597 2361 4598
rect 2486 4597 2487 4598
rect 2150 4599 2151 4600
rect 2360 4599 2361 4600
rect 2150 4601 2151 4602
rect 2228 4601 2229 4602
rect 1438 4603 1439 4604
rect 2228 4603 2229 4604
rect 2855 4603 2856 4604
rect 2870 4603 2871 4604
rect 2864 4605 2865 4606
rect 3323 4605 3324 4606
rect 2876 4607 2877 4608
rect 3270 4607 3271 4608
rect 2744 4609 2745 4610
rect 2876 4609 2877 4610
rect 2600 4611 2601 4612
rect 2744 4611 2745 4612
rect 2420 4613 2421 4614
rect 2600 4613 2601 4614
rect 2204 4615 2205 4616
rect 2420 4615 2421 4616
rect 1471 4617 1472 4618
rect 2204 4617 2205 4618
rect 1471 4619 1472 4620
rect 2012 4619 2013 4620
rect 1844 4621 1845 4622
rect 2012 4621 2013 4622
rect 1724 4623 1725 4624
rect 1844 4623 1845 4624
rect 1664 4625 1665 4626
rect 1724 4625 1725 4626
rect 1529 4627 1530 4628
rect 1664 4627 1665 4628
rect 1529 4629 1530 4630
rect 1604 4629 1605 4630
rect 2906 4629 2907 4630
rect 3158 4629 3159 4630
rect 2906 4631 2907 4632
rect 3291 4631 3292 4632
rect 2918 4633 2919 4634
rect 3215 4633 3216 4634
rect 2816 4635 2817 4636
rect 2918 4635 2919 4636
rect 2678 4637 2679 4638
rect 2816 4637 2817 4638
rect 2552 4639 2553 4640
rect 2678 4639 2679 4640
rect 2336 4641 2337 4642
rect 2552 4641 2553 4642
rect 2114 4643 2115 4644
rect 2336 4643 2337 4644
rect 1952 4645 1953 4646
rect 2114 4645 2115 4646
rect 1796 4647 1797 4648
rect 1952 4647 1953 4648
rect 1796 4649 1797 4650
rect 2894 4649 2895 4650
rect 2762 4651 2763 4652
rect 2894 4651 2895 4652
rect 2624 4653 2625 4654
rect 2762 4653 2763 4654
rect 2462 4655 2463 4656
rect 2624 4655 2625 4656
rect 2240 4657 2241 4658
rect 2462 4657 2463 4658
rect 2036 4659 2037 4660
rect 2240 4659 2241 4660
rect 1862 4661 1863 4662
rect 2036 4661 2037 4662
rect 1730 4663 1731 4664
rect 1862 4663 1863 4664
rect 1670 4665 1671 4666
rect 1730 4665 1731 4666
rect 2921 4665 2922 4666
rect 2927 4665 2928 4666
rect 2945 4665 2946 4666
rect 2999 4665 3000 4666
rect 2966 4667 2967 4668
rect 3092 4667 3093 4668
rect 2966 4669 2967 4670
rect 3237 4669 3238 4670
rect 2969 4671 2970 4672
rect 3095 4671 3096 4672
rect 3002 4673 3003 4674
rect 3116 4673 3117 4674
rect 2852 4675 2853 4676
rect 3002 4675 3003 4676
rect 2720 4677 2721 4678
rect 2852 4677 2853 4678
rect 2588 4679 2589 4680
rect 2720 4679 2721 4680
rect 2396 4681 2397 4682
rect 2588 4681 2589 4682
rect 2174 4683 2175 4684
rect 2396 4683 2397 4684
rect 1988 4685 1989 4686
rect 2174 4685 2175 4686
rect 1431 4687 1432 4688
rect 1988 4687 1989 4688
rect 3005 4687 3006 4688
rect 3288 4687 3289 4688
rect 3014 4689 3015 4690
rect 3032 4689 3033 4690
rect 3014 4691 3015 4692
rect 3212 4691 3213 4692
rect 3038 4693 3039 4694
rect 3295 4693 3296 4694
rect 2972 4695 2973 4696
rect 3038 4695 3039 4696
rect 1706 4697 1707 4698
rect 2972 4697 2973 4698
rect 1706 4699 1707 4700
rect 1718 4699 1719 4700
rect 1658 4701 1659 4702
rect 1718 4701 1719 4702
rect 1658 4703 1659 4704
rect 3305 4703 3306 4704
rect 2996 4705 2997 4706
rect 3304 4705 3305 4706
rect 2942 4707 2943 4708
rect 2996 4707 2997 4708
rect 2942 4709 2943 4710
rect 3274 4709 3275 4710
rect 3056 4711 3057 4712
rect 3377 4711 3378 4712
rect 3062 4713 3063 4714
rect 3158 4713 3159 4714
rect 2936 4715 2937 4716
rect 3062 4715 3063 4716
rect 2798 4717 2799 4718
rect 2936 4717 2937 4718
rect 2660 4719 2661 4720
rect 2798 4719 2799 4720
rect 2498 4721 2499 4722
rect 2660 4721 2661 4722
rect 2318 4723 2319 4724
rect 2498 4723 2499 4724
rect 2090 4725 2091 4726
rect 2318 4725 2319 4726
rect 2090 4727 2091 4728
rect 3298 4727 3299 4728
rect 3068 4729 3069 4730
rect 3152 4729 3153 4730
rect 2948 4731 2949 4732
rect 3068 4731 3069 4732
rect 2804 4733 2805 4734
rect 2948 4733 2949 4734
rect 2672 4735 2673 4736
rect 2804 4735 2805 4736
rect 2528 4737 2529 4738
rect 2672 4737 2673 4738
rect 2366 4739 2367 4740
rect 2528 4739 2529 4740
rect 2144 4741 2145 4742
rect 2366 4741 2367 4742
rect 1958 4743 1959 4744
rect 2144 4743 2145 4744
rect 1802 4745 1803 4746
rect 1958 4745 1959 4746
rect 1802 4747 1803 4748
rect 2900 4747 2901 4748
rect 2768 4749 2769 4750
rect 2900 4749 2901 4750
rect 2630 4751 2631 4752
rect 2768 4751 2769 4752
rect 2468 4753 2469 4754
rect 2630 4753 2631 4754
rect 2234 4755 2235 4756
rect 2468 4755 2469 4756
rect 2234 4757 2235 4758
rect 2312 4757 2313 4758
rect 2096 4759 2097 4760
rect 2312 4759 2313 4760
rect 1934 4761 1935 4762
rect 2096 4761 2097 4762
rect 1790 4763 1791 4764
rect 1934 4763 1935 4764
rect 1700 4765 1701 4766
rect 1790 4765 1791 4766
rect 1598 4767 1599 4768
rect 1700 4767 1701 4768
rect 1568 4769 1569 4770
rect 1598 4769 1599 4770
rect 3074 4769 3075 4770
rect 3277 4769 3278 4770
rect 3080 4771 3081 4772
rect 3249 4771 3250 4772
rect 2990 4773 2991 4774
rect 3080 4773 3081 4774
rect 2990 4775 2991 4776
rect 3384 4775 3385 4776
rect 3098 4777 3099 4778
rect 3188 4777 3189 4778
rect 2978 4779 2979 4780
rect 3098 4779 3099 4780
rect 2888 4781 2889 4782
rect 2978 4781 2979 4782
rect 2756 4783 2757 4784
rect 2888 4783 2889 4784
rect 2666 4785 2667 4786
rect 2756 4785 2757 4786
rect 2510 4787 2511 4788
rect 2666 4787 2667 4788
rect 2300 4789 2301 4790
rect 2510 4789 2511 4790
rect 2132 4791 2133 4792
rect 2300 4791 2301 4792
rect 2072 4793 2073 4794
rect 2132 4793 2133 4794
rect 1916 4795 1917 4796
rect 2072 4795 2073 4796
rect 1916 4797 1917 4798
rect 2618 4797 2619 4798
rect 2444 4799 2445 4800
rect 2618 4799 2619 4800
rect 2258 4801 2259 4802
rect 2444 4801 2445 4802
rect 2066 4803 2067 4804
rect 2258 4803 2259 4804
rect 2066 4805 2067 4806
rect 2378 4805 2379 4806
rect 2168 4807 2169 4808
rect 2378 4807 2379 4808
rect 1982 4809 1983 4810
rect 2168 4809 2169 4810
rect 1826 4811 1827 4812
rect 1982 4811 1983 4812
rect 1736 4813 1737 4814
rect 1826 4813 1827 4814
rect 1688 4815 1689 4816
rect 1736 4815 1737 4816
rect 1688 4817 1689 4818
rect 1694 4817 1695 4818
rect 3101 4817 3102 4818
rect 3191 4817 3192 4818
rect 3104 4819 3105 4820
rect 3215 4819 3216 4820
rect 2984 4821 2985 4822
rect 3104 4821 3105 4822
rect 3128 4821 3129 4822
rect 3224 4821 3225 4822
rect 3050 4823 3051 4824
rect 3128 4823 3129 4824
rect 2912 4825 2913 4826
rect 3050 4825 3051 4826
rect 2774 4827 2775 4828
rect 2912 4827 2913 4828
rect 2774 4829 2775 4830
rect 3302 4829 3303 4830
rect 3134 4831 3135 4832
rect 3227 4831 3228 4832
rect 3026 4833 3027 4834
rect 3134 4833 3135 4834
rect 2882 4835 2883 4836
rect 3026 4835 3027 4836
rect 2750 4837 2751 4838
rect 2882 4837 2883 4838
rect 2750 4839 2751 4840
rect 2780 4839 2781 4840
rect 2642 4841 2643 4842
rect 2780 4841 2781 4842
rect 2642 4843 2643 4844
rect 3360 4843 3361 4844
rect 3140 4845 3141 4846
rect 3161 4845 3162 4846
rect 3164 4845 3165 4846
rect 3243 4845 3244 4846
rect 3107 4847 3108 4848
rect 3164 4847 3165 4848
rect 3176 4847 3177 4848
rect 3320 4847 3321 4848
rect 3086 4849 3087 4850
rect 3176 4849 3177 4850
rect 3194 4849 3195 4850
rect 3273 4849 3274 4850
rect 3110 4851 3111 4852
rect 3194 4851 3195 4852
rect 3008 4853 3009 4854
rect 3110 4853 3111 4854
rect 2954 4855 2955 4856
rect 3008 4855 3009 4856
rect 2810 4857 2811 4858
rect 2954 4857 2955 4858
rect 2732 4859 2733 4860
rect 2810 4859 2811 4860
rect 2606 4861 2607 4862
rect 2732 4861 2733 4862
rect 2432 4863 2433 4864
rect 2606 4863 2607 4864
rect 2276 4865 2277 4866
rect 2432 4865 2433 4866
rect 2054 4867 2055 4868
rect 2276 4867 2277 4868
rect 2054 4869 2055 4870
rect 2330 4869 2331 4870
rect 2156 4871 2157 4872
rect 2330 4871 2331 4872
rect 2156 4873 2157 4874
rect 3231 4873 3232 4874
rect 3170 4875 3171 4876
rect 3230 4875 3231 4876
rect 3197 4877 3198 4878
rect 3276 4877 3277 4878
rect 3113 4879 3114 4880
rect 3197 4879 3198 4880
rect 3200 4879 3201 4880
rect 3294 4879 3295 4880
rect 3200 4881 3201 4882
rect 3221 4881 3222 4882
rect 3203 4883 3204 4884
rect 3224 4883 3225 4884
rect 3044 4885 3045 4886
rect 3203 4885 3204 4886
rect 1475 4887 1476 4888
rect 3044 4887 3045 4888
rect 3206 4887 3207 4888
rect 3285 4887 3286 4888
rect 3122 4889 3123 4890
rect 3206 4889 3207 4890
rect 3020 4891 3021 4892
rect 3122 4891 3123 4892
rect 2879 4893 2880 4894
rect 3020 4893 3021 4894
rect 3209 4893 3210 4894
rect 3288 4893 3289 4894
rect 3212 4895 3213 4896
rect 3307 4895 3308 4896
rect 3218 4897 3219 4898
rect 3233 4897 3234 4898
rect 3146 4899 3147 4900
rect 3218 4899 3219 4900
rect 3240 4899 3241 4900
rect 3314 4899 3315 4900
rect 3246 4901 3247 4902
rect 3317 4901 3318 4902
rect 3261 4903 3262 4904
rect 3354 4903 3355 4904
rect 3182 4905 3183 4906
rect 3261 4905 3262 4906
rect 3264 4905 3265 4906
rect 3357 4905 3358 4906
rect 3267 4907 3268 4908
rect 3297 4907 3298 4908
rect 3291 4909 3292 4910
rect 3363 4909 3364 4910
rect 3330 4911 3331 4912
rect 3381 4911 3382 4912
rect 3336 4913 3337 4914
rect 3388 4913 3389 4914
rect 3342 4915 3343 4916
rect 3391 4915 3392 4916
rect 1434 4924 1435 4925
rect 1952 4924 1953 4925
rect 1438 4926 1439 4927
rect 2138 4926 2139 4927
rect 1447 4928 1448 4929
rect 2060 4928 2061 4929
rect 1471 4930 1472 4931
rect 2006 4930 2007 4931
rect 1478 4932 1479 4933
rect 1970 4932 1971 4933
rect 1477 4934 1478 4935
rect 1988 4934 1989 4935
rect 1482 4936 1483 4937
rect 2156 4936 2157 4937
rect 1488 4938 1489 4939
rect 2327 4938 2328 4939
rect 1491 4940 1492 4941
rect 2282 4940 2283 4941
rect 1503 4942 1504 4943
rect 1748 4942 1749 4943
rect 1514 4944 1515 4945
rect 2312 4944 2313 4945
rect 1510 4946 1511 4947
rect 2312 4946 2313 4947
rect 1517 4948 1518 4949
rect 2879 4948 2880 4949
rect 1519 4950 1520 4951
rect 2192 4950 2193 4951
rect 1526 4952 1527 4953
rect 1904 4952 1905 4953
rect 1526 4954 1527 4955
rect 2504 4954 2505 4955
rect 1529 4956 1530 4957
rect 3014 4956 3015 4957
rect 1538 4958 1539 4959
rect 1886 4958 1887 4959
rect 1541 4960 1542 4961
rect 1838 4960 1839 4961
rect 1468 4962 1469 4963
rect 1838 4962 1839 4963
rect 1462 4964 1463 4965
rect 1468 4964 1469 4965
rect 1456 4966 1457 4967
rect 1462 4966 1463 4967
rect 1450 4968 1451 4969
rect 1456 4968 1457 4969
rect 1556 4968 1557 4969
rect 2825 4968 2826 4969
rect 1574 4970 1575 4971
rect 1586 4970 1587 4971
rect 1580 4972 1581 4973
rect 2147 4972 2148 4973
rect 1634 4974 1635 4975
rect 1646 4974 1647 4975
rect 1622 4976 1623 4977
rect 1634 4976 1635 4977
rect 1610 4978 1611 4979
rect 1622 4978 1623 4979
rect 1598 4980 1599 4981
rect 1610 4980 1611 4981
rect 1562 4982 1563 4983
rect 1598 4982 1599 4983
rect 1550 4984 1551 4985
rect 1562 4984 1563 4985
rect 1652 4984 1653 4985
rect 1670 4984 1671 4985
rect 1640 4986 1641 4987
rect 1652 4986 1653 4987
rect 1628 4988 1629 4989
rect 1640 4988 1641 4989
rect 1616 4990 1617 4991
rect 1628 4990 1629 4991
rect 1694 4990 1695 4991
rect 1718 4990 1719 4991
rect 1742 4990 1743 4991
rect 1766 4990 1767 4991
rect 1742 4992 1743 4993
rect 1790 4992 1791 4993
rect 1748 4994 1749 4995
rect 1754 4994 1755 4995
rect 1688 4996 1689 4997
rect 1754 4996 1755 4997
rect 1481 4998 1482 4999
rect 1688 4998 1689 4999
rect 1790 4998 1791 4999
rect 1844 4998 1845 4999
rect 1829 5000 1830 5001
rect 2045 5000 2046 5001
rect 1844 5002 1845 5003
rect 2072 5002 2073 5003
rect 1904 5004 1905 5005
rect 2288 5004 2289 5005
rect 1661 5006 1662 5007
rect 2288 5006 2289 5007
rect 1907 5008 1908 5009
rect 2291 5008 2292 5009
rect 1910 5010 1911 5011
rect 2228 5010 2229 5011
rect 1937 5012 1938 5013
rect 2231 5012 2232 5013
rect 1952 5014 1953 5015
rect 2240 5014 2241 5015
rect 1970 5016 1971 5017
rect 2348 5016 2349 5017
rect 1976 5018 1977 5019
rect 2192 5018 2193 5019
rect 1976 5020 1977 5021
rect 2342 5020 2343 5021
rect 1982 5022 1983 5023
rect 2156 5022 2157 5023
rect 1982 5024 1983 5025
rect 2204 5024 2205 5025
rect 1988 5026 1989 5027
rect 2366 5026 2367 5027
rect 2006 5028 2007 5029
rect 2360 5028 2361 5029
rect 2060 5030 2061 5031
rect 2264 5030 2265 5031
rect 2069 5032 2070 5033
rect 2273 5032 2274 5033
rect 2072 5034 2073 5035
rect 2300 5034 2301 5035
rect 2102 5036 2103 5037
rect 2348 5036 2349 5037
rect 2102 5038 2103 5039
rect 2402 5038 2403 5039
rect 2132 5040 2133 5041
rect 2360 5040 2361 5041
rect 2132 5042 2133 5043
rect 2408 5042 2409 5043
rect 2126 5044 2127 5045
rect 2408 5044 2409 5045
rect 2126 5046 2127 5047
rect 2462 5046 2463 5047
rect 2138 5048 2139 5049
rect 2420 5048 2421 5049
rect 2150 5050 2151 5051
rect 2228 5050 2229 5051
rect 2150 5052 2151 5053
rect 2426 5052 2427 5053
rect 2159 5054 2160 5055
rect 2573 5054 2574 5055
rect 2180 5056 2181 5057
rect 2300 5056 2301 5057
rect 2090 5058 2091 5059
rect 2180 5058 2181 5059
rect 2090 5060 2091 5061
rect 2450 5060 2451 5061
rect 2204 5062 2205 5063
rect 2510 5062 2511 5063
rect 2234 5064 2235 5065
rect 2240 5064 2241 5065
rect 2234 5066 2235 5067
rect 3326 5066 3327 5067
rect 2264 5068 2265 5069
rect 2540 5068 2541 5069
rect 2282 5070 2283 5071
rect 2294 5070 2295 5071
rect 2294 5072 2295 5073
rect 2492 5072 2493 5073
rect 1868 5074 1869 5075
rect 2492 5074 2493 5075
rect 2342 5076 2343 5077
rect 2594 5076 2595 5077
rect 1760 5078 1761 5079
rect 2594 5078 2595 5079
rect 1760 5080 1761 5081
rect 1862 5080 1863 5081
rect 1862 5082 1863 5083
rect 2144 5082 2145 5083
rect 2144 5084 2145 5085
rect 2474 5084 2475 5085
rect 1874 5086 1875 5087
rect 2474 5086 2475 5087
rect 1658 5088 1659 5089
rect 1874 5088 1875 5089
rect 1604 5090 1605 5091
rect 1658 5090 1659 5091
rect 1592 5092 1593 5093
rect 1604 5092 1605 5093
rect 1433 5094 1434 5095
rect 1592 5094 1593 5095
rect 2357 5094 2358 5095
rect 3035 5094 3036 5095
rect 2279 5096 2280 5097
rect 2357 5096 2358 5097
rect 2366 5096 2367 5097
rect 2600 5096 2601 5097
rect 2216 5098 2217 5099
rect 2600 5098 2601 5099
rect 2216 5100 2217 5101
rect 2480 5100 2481 5101
rect 1856 5102 1857 5103
rect 2480 5102 2481 5103
rect 1856 5104 1857 5105
rect 2108 5104 2109 5105
rect 2108 5106 2109 5107
rect 2354 5106 2355 5107
rect 1475 5108 1476 5109
rect 2354 5108 2355 5109
rect 1474 5110 1475 5111
rect 2114 5110 2115 5111
rect 2114 5112 2115 5113
rect 3451 5112 3452 5113
rect 2402 5114 2403 5115
rect 3468 5114 3469 5115
rect 2420 5116 2421 5117
rect 2630 5116 2631 5117
rect 2426 5118 2427 5119
rect 2624 5118 2625 5119
rect 2444 5120 2445 5121
rect 3304 5120 3305 5121
rect 2444 5122 2445 5123
rect 2528 5122 2529 5123
rect 1994 5124 1995 5125
rect 2528 5124 2529 5125
rect 1994 5126 1995 5127
rect 2174 5126 2175 5127
rect 1889 5128 1890 5129
rect 2174 5128 2175 5129
rect 2450 5128 2451 5129
rect 2654 5128 2655 5129
rect 2462 5130 2463 5131
rect 2642 5130 2643 5131
rect 2468 5132 2469 5133
rect 3454 5132 3455 5133
rect 2024 5134 2025 5135
rect 2468 5134 2469 5135
rect 2024 5136 2025 5137
rect 2210 5136 2211 5137
rect 2210 5138 2211 5139
rect 2432 5138 2433 5139
rect 2432 5140 2433 5141
rect 2570 5140 2571 5141
rect 1880 5142 1881 5143
rect 2570 5142 2571 5143
rect 1880 5144 1881 5145
rect 2084 5144 2085 5145
rect 2084 5146 2085 5147
rect 2306 5146 2307 5147
rect 1507 5148 1508 5149
rect 2306 5148 2307 5149
rect 2504 5148 2505 5149
rect 2660 5148 2661 5149
rect 2186 5150 2187 5151
rect 2660 5150 2661 5151
rect 2120 5152 2121 5153
rect 2186 5152 2187 5153
rect 2120 5154 2121 5155
rect 3323 5154 3324 5155
rect 2510 5156 2511 5157
rect 2666 5156 2667 5157
rect 1541 5158 1542 5159
rect 2666 5158 2667 5159
rect 2540 5160 2541 5161
rect 3333 5160 3334 5161
rect 2552 5162 2553 5163
rect 3381 5162 3382 5163
rect 2552 5164 2553 5165
rect 2684 5164 2685 5165
rect 2576 5166 2577 5167
rect 3458 5166 3459 5167
rect 2576 5168 2577 5169
rect 2672 5168 2673 5169
rect 1940 5170 1941 5171
rect 2672 5170 2673 5171
rect 1940 5172 1941 5173
rect 2318 5172 2319 5173
rect 2318 5174 2319 5175
rect 2582 5174 2583 5175
rect 2048 5176 2049 5177
rect 2582 5176 2583 5177
rect 2048 5178 2049 5179
rect 2414 5178 2415 5179
rect 2414 5180 2415 5181
rect 3367 5180 3368 5181
rect 2618 5182 2619 5183
rect 3370 5182 3371 5183
rect 2030 5184 2031 5185
rect 2618 5184 2619 5185
rect 2030 5186 2031 5187
rect 2378 5186 2379 5187
rect 2378 5188 2379 5189
rect 2606 5188 2607 5189
rect 2606 5190 2607 5191
rect 2708 5190 2709 5191
rect 2624 5192 2625 5193
rect 2738 5192 2739 5193
rect 2630 5194 2631 5195
rect 2714 5194 2715 5195
rect 2642 5196 2643 5197
rect 2678 5196 2679 5197
rect 2654 5198 2655 5199
rect 2732 5198 2733 5199
rect 1850 5200 1851 5201
rect 2732 5200 2733 5201
rect 1424 5202 1425 5203
rect 1850 5202 1851 5203
rect 1423 5204 1424 5205
rect 1556 5204 1557 5205
rect 2678 5204 2679 5205
rect 2780 5204 2781 5205
rect 1512 5206 1513 5207
rect 2780 5206 2781 5207
rect 2684 5208 2685 5209
rect 3307 5208 3308 5209
rect 2708 5210 2709 5211
rect 2798 5210 2799 5211
rect 2714 5212 2715 5213
rect 2792 5212 2793 5213
rect 2738 5214 2739 5215
rect 2828 5214 2829 5215
rect 2744 5216 2745 5217
rect 3407 5216 3408 5217
rect 2744 5218 2745 5219
rect 2834 5218 2835 5219
rect 2762 5220 2763 5221
rect 3429 5220 3430 5221
rect 2762 5222 2763 5223
rect 2852 5222 2853 5223
rect 2768 5224 2769 5225
rect 3363 5224 3364 5225
rect 2756 5226 2757 5227
rect 2768 5226 2769 5227
rect 2792 5226 2793 5227
rect 2864 5226 2865 5227
rect 2798 5228 2799 5229
rect 2876 5228 2877 5229
rect 1500 5230 1501 5231
rect 2876 5230 2877 5231
rect 1494 5232 1495 5233
rect 1500 5232 1501 5233
rect 2816 5232 2817 5233
rect 3461 5232 3462 5233
rect 1946 5234 1947 5235
rect 2816 5234 2817 5235
rect 1946 5236 1947 5237
rect 2324 5236 2325 5237
rect 2324 5238 2325 5239
rect 2588 5238 2589 5239
rect 2054 5240 2055 5241
rect 2588 5240 2589 5241
rect 2054 5242 2055 5243
rect 3465 5242 3466 5243
rect 2828 5244 2829 5245
rect 2900 5244 2901 5245
rect 2834 5246 2835 5247
rect 2906 5246 2907 5247
rect 2846 5248 2847 5249
rect 2888 5248 2889 5249
rect 2750 5250 2751 5251
rect 2888 5250 2889 5251
rect 2750 5252 2751 5253
rect 2840 5252 2841 5253
rect 1916 5254 1917 5255
rect 2840 5254 2841 5255
rect 1916 5256 1917 5257
rect 2270 5256 2271 5257
rect 2270 5258 2271 5259
rect 2516 5258 2517 5259
rect 2000 5260 2001 5261
rect 2516 5260 2517 5261
rect 2000 5262 2001 5263
rect 2384 5262 2385 5263
rect 1427 5264 1428 5265
rect 2384 5264 2385 5265
rect 1426 5266 1427 5267
rect 1877 5266 1878 5267
rect 2852 5266 2853 5267
rect 2894 5266 2895 5267
rect 2858 5268 2859 5269
rect 3400 5268 3401 5269
rect 2858 5270 2859 5271
rect 2930 5270 2931 5271
rect 1898 5272 1899 5273
rect 2930 5272 2931 5273
rect 1898 5274 1899 5275
rect 2222 5274 2223 5275
rect 2222 5276 2223 5277
rect 2252 5276 2253 5277
rect 2252 5278 2253 5279
rect 3327 5278 3328 5279
rect 2864 5280 2865 5281
rect 2936 5280 2937 5281
rect 2870 5282 2871 5283
rect 3444 5282 3445 5283
rect 2870 5284 2871 5285
rect 2912 5284 2913 5285
rect 2894 5286 2895 5287
rect 2948 5286 2949 5287
rect 1706 5288 1707 5289
rect 2948 5288 2949 5289
rect 1706 5290 1707 5291
rect 1730 5290 1731 5291
rect 1730 5292 1731 5293
rect 2321 5292 2322 5293
rect 2900 5292 2901 5293
rect 2954 5292 2955 5293
rect 1832 5294 1833 5295
rect 2954 5294 2955 5295
rect 1431 5296 1432 5297
rect 1832 5296 1833 5297
rect 1430 5298 1431 5299
rect 1538 5298 1539 5299
rect 2912 5298 2913 5299
rect 2966 5298 2967 5299
rect 2921 5300 2922 5301
rect 3107 5300 3108 5301
rect 2924 5302 2925 5303
rect 3240 5302 3241 5303
rect 2918 5304 2919 5305
rect 2924 5304 2925 5305
rect 2918 5306 2919 5307
rect 3237 5306 3238 5307
rect 2942 5308 2943 5309
rect 3384 5308 3385 5309
rect 1964 5310 1965 5311
rect 2942 5310 2943 5311
rect 1964 5312 1965 5313
rect 2198 5312 2199 5313
rect 2078 5314 2079 5315
rect 2198 5314 2199 5315
rect 2078 5316 2079 5317
rect 2330 5316 2331 5317
rect 2096 5318 2097 5319
rect 2330 5318 2331 5319
rect 2096 5320 2097 5321
rect 2456 5320 2457 5321
rect 2456 5322 2457 5323
rect 2558 5322 2559 5323
rect 2558 5324 2559 5325
rect 2636 5324 2637 5325
rect 2636 5326 2637 5327
rect 2702 5326 2703 5327
rect 2702 5328 2703 5329
rect 2774 5328 2775 5329
rect 2774 5330 2775 5331
rect 2804 5330 2805 5331
rect 2804 5332 2805 5333
rect 2882 5332 2883 5333
rect 2696 5334 2697 5335
rect 2882 5334 2883 5335
rect 2696 5336 2697 5337
rect 3323 5336 3324 5337
rect 2960 5338 2961 5339
rect 3002 5338 3003 5339
rect 1712 5340 1713 5341
rect 3002 5340 3003 5341
rect 1712 5342 1713 5343
rect 1736 5342 1737 5343
rect 1664 5344 1665 5345
rect 1736 5344 1737 5345
rect 2963 5344 2964 5345
rect 3005 5344 3006 5345
rect 2966 5346 2967 5347
rect 2972 5346 2973 5347
rect 1808 5348 1809 5349
rect 2972 5348 2973 5349
rect 1808 5350 1809 5351
rect 1958 5350 1959 5351
rect 1958 5352 1959 5353
rect 2336 5352 2337 5353
rect 2336 5354 2337 5355
rect 2522 5354 2523 5355
rect 2066 5356 2067 5357
rect 2522 5356 2523 5357
rect 2066 5358 2067 5359
rect 2168 5358 2169 5359
rect 2168 5360 2169 5361
rect 2246 5360 2247 5361
rect 2246 5362 2247 5363
rect 2498 5362 2499 5363
rect 1928 5364 1929 5365
rect 2498 5364 2499 5365
rect 1928 5366 1929 5367
rect 2258 5366 2259 5367
rect 2258 5368 2259 5369
rect 2546 5368 2547 5369
rect 2546 5370 2547 5371
rect 2690 5370 2691 5371
rect 2690 5372 2691 5373
rect 2786 5372 2787 5373
rect 2786 5374 2787 5375
rect 3447 5374 3448 5375
rect 2981 5376 2982 5377
rect 3023 5376 3024 5377
rect 2429 5378 2430 5379
rect 3023 5378 3024 5379
rect 2984 5380 2985 5381
rect 3026 5380 3027 5381
rect 1778 5382 1779 5383
rect 3026 5382 3027 5383
rect 1444 5384 1445 5385
rect 1778 5384 1779 5385
rect 2999 5384 3000 5385
rect 3221 5384 3222 5385
rect 3014 5386 3015 5387
rect 3056 5386 3057 5387
rect 3032 5388 3033 5389
rect 3146 5388 3147 5389
rect 1796 5390 1797 5391
rect 3032 5390 3033 5391
rect 1796 5392 1797 5393
rect 1826 5392 1827 5393
rect 1826 5394 1827 5395
rect 2042 5394 2043 5395
rect 2042 5396 2043 5397
rect 2372 5396 2373 5397
rect 2372 5398 2373 5399
rect 2612 5398 2613 5399
rect 2612 5400 2613 5401
rect 2726 5400 2727 5401
rect 2726 5402 2727 5403
rect 2822 5402 2823 5403
rect 1515 5404 1516 5405
rect 2822 5404 2823 5405
rect 3050 5404 3051 5405
rect 3374 5404 3375 5405
rect 1820 5406 1821 5407
rect 3050 5406 3051 5407
rect 1820 5408 1821 5409
rect 2036 5408 2037 5409
rect 2036 5410 2037 5411
rect 2390 5410 2391 5411
rect 2162 5412 2163 5413
rect 2390 5412 2391 5413
rect 1485 5414 1486 5415
rect 2162 5414 2163 5415
rect 1484 5416 1485 5417
rect 1676 5416 1677 5417
rect 1676 5418 1677 5419
rect 3422 5418 3423 5419
rect 3056 5420 3057 5421
rect 3068 5420 3069 5421
rect 3068 5422 3069 5423
rect 3297 5422 3298 5423
rect 3098 5424 3099 5425
rect 3140 5424 3141 5425
rect 3116 5426 3117 5427
rect 3419 5426 3420 5427
rect 3104 5428 3105 5429
rect 3116 5428 3117 5429
rect 1700 5430 1701 5431
rect 3104 5430 3105 5431
rect 1700 5432 1701 5433
rect 1724 5432 1725 5433
rect 1724 5434 1725 5435
rect 1772 5434 1773 5435
rect 1417 5436 1418 5437
rect 1772 5436 1773 5437
rect 3170 5436 3171 5437
rect 3278 5436 3279 5437
rect 3170 5438 3171 5439
rect 3311 5438 3312 5439
rect 3182 5440 3183 5441
rect 3314 5440 3315 5441
rect 3188 5442 3189 5443
rect 3248 5442 3249 5443
rect 3128 5444 3129 5445
rect 3188 5444 3189 5445
rect 3038 5446 3039 5447
rect 3128 5446 3129 5447
rect 1437 5448 1438 5449
rect 3038 5448 3039 5449
rect 3203 5448 3204 5449
rect 3263 5448 3264 5449
rect 3206 5450 3207 5451
rect 3266 5450 3267 5451
rect 3158 5452 3159 5453
rect 3206 5452 3207 5453
rect 3134 5454 3135 5455
rect 3158 5454 3159 5455
rect 3044 5456 3045 5457
rect 3134 5456 3135 5457
rect 1802 5458 1803 5459
rect 3044 5458 3045 5459
rect 1802 5460 1803 5461
rect 1934 5460 1935 5461
rect 1441 5462 1442 5463
rect 1934 5462 1935 5463
rect 1440 5464 1441 5465
rect 2012 5464 2013 5465
rect 2012 5466 2013 5467
rect 2396 5466 2397 5467
rect 2396 5468 2397 5469
rect 3426 5468 3427 5469
rect 3212 5470 3213 5471
rect 3308 5470 3309 5471
rect 3164 5472 3165 5473
rect 3212 5472 3213 5473
rect 3122 5474 3123 5475
rect 3164 5474 3165 5475
rect 3080 5476 3081 5477
rect 3122 5476 3123 5477
rect 3074 5478 3075 5479
rect 3080 5478 3081 5479
rect 3062 5480 3063 5481
rect 3074 5480 3075 5481
rect 1522 5482 1523 5483
rect 3062 5482 3063 5483
rect 3215 5482 3216 5483
rect 3311 5482 3312 5483
rect 3218 5484 3219 5485
rect 3314 5484 3315 5485
rect 2996 5486 2997 5487
rect 3218 5486 3219 5487
rect 1814 5488 1815 5489
rect 2996 5488 2997 5489
rect 1529 5490 1530 5491
rect 1814 5490 1815 5491
rect 3224 5490 3225 5491
rect 3296 5490 3297 5491
rect 3176 5492 3177 5493
rect 3224 5492 3225 5493
rect 3236 5492 3237 5493
rect 3377 5492 3378 5493
rect 3243 5494 3244 5495
rect 3333 5494 3334 5495
rect 3251 5496 3252 5497
rect 3395 5496 3396 5497
rect 2990 5498 2991 5499
rect 3396 5498 3397 5499
rect 2990 5500 2991 5501
rect 3393 5500 3394 5501
rect 3273 5502 3274 5503
rect 3369 5502 3370 5503
rect 3272 5504 3273 5505
rect 3300 5504 3301 5505
rect 3276 5506 3277 5507
rect 3372 5506 3373 5507
rect 3194 5508 3195 5509
rect 3275 5508 3276 5509
rect 3194 5510 3195 5511
rect 3197 5510 3198 5511
rect 3285 5510 3286 5511
rect 3381 5510 3382 5511
rect 3230 5512 3231 5513
rect 3284 5512 3285 5513
rect 3191 5514 3192 5515
rect 3230 5514 3231 5515
rect 3288 5514 3289 5515
rect 3384 5514 3385 5515
rect 3317 5516 3318 5517
rect 3413 5516 3414 5517
rect 3320 5518 3321 5519
rect 3339 5518 3340 5519
rect 2720 5520 2721 5521
rect 3320 5520 3321 5521
rect 1922 5522 1923 5523
rect 2720 5522 2721 5523
rect 1922 5524 1923 5525
rect 2276 5524 2277 5525
rect 2276 5526 2277 5527
rect 2486 5526 2487 5527
rect 2486 5528 2487 5529
rect 2534 5528 2535 5529
rect 2534 5530 2535 5531
rect 2648 5530 2649 5531
rect 2438 5532 2439 5533
rect 2648 5532 2649 5533
rect 2018 5534 2019 5535
rect 2438 5534 2439 5535
rect 1886 5536 1887 5537
rect 2018 5536 2019 5537
rect 3330 5536 3331 5537
rect 3398 5536 3399 5537
rect 2936 5538 2937 5539
rect 3330 5538 3331 5539
rect 3336 5538 3337 5539
rect 3441 5538 3442 5539
rect 3342 5540 3343 5541
rect 3438 5540 3439 5541
rect 3354 5542 3355 5543
rect 3391 5542 3392 5543
rect 3294 5544 3295 5545
rect 3390 5544 3391 5545
rect 3357 5546 3358 5547
rect 3388 5546 3389 5547
rect 3261 5548 3262 5549
rect 3357 5548 3358 5549
rect 3200 5550 3201 5551
rect 3260 5550 3261 5551
rect 3152 5552 3153 5553
rect 3200 5552 3201 5553
rect 3110 5554 3111 5555
rect 3152 5554 3153 5555
rect 3008 5556 3009 5557
rect 3110 5556 3111 5557
rect 2978 5558 2979 5559
rect 3008 5558 3009 5559
rect 2978 5560 2979 5561
rect 3020 5560 3021 5561
rect 1784 5562 1785 5563
rect 3020 5562 3021 5563
rect 1784 5564 1785 5565
rect 1892 5564 1893 5565
rect 1420 5566 1421 5567
rect 1892 5566 1893 5567
rect 3291 5566 3292 5567
rect 3387 5566 3388 5567
rect 3233 5568 3234 5569
rect 3290 5568 3291 5569
rect 3360 5568 3361 5569
rect 3416 5568 3417 5569
rect 3403 5570 3404 5571
rect 3410 5570 3411 5571
rect 1420 5579 1421 5580
rect 1832 5579 1833 5580
rect 1423 5581 1424 5582
rect 1919 5581 1920 5582
rect 1433 5583 1434 5584
rect 1907 5583 1908 5584
rect 1434 5585 1435 5586
rect 1694 5585 1695 5586
rect 1437 5587 1438 5588
rect 1967 5587 1968 5588
rect 1438 5589 1439 5590
rect 2780 5589 2781 5590
rect 1440 5591 1441 5592
rect 2594 5591 2595 5592
rect 1441 5593 1442 5594
rect 1592 5593 1593 5594
rect 1444 5595 1445 5596
rect 1652 5595 1653 5596
rect 1445 5597 1446 5598
rect 1580 5597 1581 5598
rect 1481 5599 1482 5600
rect 2573 5599 2574 5600
rect 1482 5601 1483 5602
rect 2180 5601 2181 5602
rect 1477 5603 1478 5604
rect 2180 5603 2181 5604
rect 1484 5605 1485 5606
rect 2567 5605 2568 5606
rect 1488 5607 1489 5608
rect 2246 5607 2247 5608
rect 1515 5609 1516 5610
rect 2996 5609 2997 5610
rect 1519 5611 1520 5612
rect 1556 5611 1557 5612
rect 1522 5613 1523 5614
rect 3020 5613 3021 5614
rect 1532 5615 1533 5616
rect 1658 5615 1659 5616
rect 1535 5617 1536 5618
rect 1652 5617 1653 5618
rect 1541 5619 1542 5620
rect 2672 5619 2673 5620
rect 1544 5621 1545 5622
rect 1550 5621 1551 5622
rect 1544 5623 1545 5624
rect 2768 5623 2769 5624
rect 1547 5625 1548 5626
rect 2234 5625 2235 5626
rect 1556 5627 1557 5628
rect 1562 5627 1563 5628
rect 1568 5627 1569 5628
rect 1877 5627 1878 5628
rect 1580 5629 1581 5630
rect 1586 5629 1587 5630
rect 1592 5629 1593 5630
rect 1604 5629 1605 5630
rect 1604 5631 1605 5632
rect 1889 5631 1890 5632
rect 1426 5633 1427 5634
rect 1889 5633 1890 5634
rect 1427 5635 1428 5636
rect 1874 5635 1875 5636
rect 1616 5637 1617 5638
rect 1622 5637 1623 5638
rect 1622 5639 1623 5640
rect 1628 5639 1629 5640
rect 1598 5641 1599 5642
rect 1628 5641 1629 5642
rect 1598 5643 1599 5644
rect 1610 5643 1611 5644
rect 1430 5645 1431 5646
rect 1610 5645 1611 5646
rect 1664 5645 1665 5646
rect 1676 5645 1677 5646
rect 1676 5647 1677 5648
rect 1688 5647 1689 5648
rect 1682 5649 1683 5650
rect 1700 5649 1701 5650
rect 1688 5651 1689 5652
rect 1706 5651 1707 5652
rect 1694 5653 1695 5654
rect 1712 5653 1713 5654
rect 1700 5655 1701 5656
rect 1730 5655 1731 5656
rect 1712 5657 1713 5658
rect 1724 5657 1725 5658
rect 1526 5659 1527 5660
rect 1724 5659 1725 5660
rect 1525 5661 1526 5662
rect 2072 5661 2073 5662
rect 1718 5663 1719 5664
rect 1766 5663 1767 5664
rect 1730 5665 1731 5666
rect 1742 5665 1743 5666
rect 1742 5667 1743 5668
rect 1748 5667 1749 5668
rect 1670 5669 1671 5670
rect 1748 5669 1749 5670
rect 1754 5669 1755 5670
rect 3396 5669 3397 5670
rect 1754 5671 1755 5672
rect 2876 5671 2877 5672
rect 1766 5673 1767 5674
rect 1796 5673 1797 5674
rect 1736 5675 1737 5676
rect 1796 5675 1797 5676
rect 1431 5677 1432 5678
rect 1736 5677 1737 5678
rect 1808 5677 1809 5678
rect 1832 5677 1833 5678
rect 1485 5679 1486 5680
rect 1808 5679 1809 5680
rect 1868 5679 1869 5680
rect 2069 5679 2070 5680
rect 1874 5681 1875 5682
rect 1880 5681 1881 5682
rect 1880 5683 1881 5684
rect 2066 5683 2067 5684
rect 1886 5685 1887 5686
rect 2957 5685 2958 5686
rect 1424 5687 1425 5688
rect 1886 5687 1887 5688
rect 1925 5687 1926 5688
rect 1937 5687 1938 5688
rect 1988 5687 1989 5688
rect 3461 5687 3462 5688
rect 1940 5689 1941 5690
rect 1988 5689 1989 5690
rect 1928 5691 1929 5692
rect 1940 5691 1941 5692
rect 1928 5693 1929 5694
rect 1994 5693 1995 5694
rect 1946 5695 1947 5696
rect 1994 5695 1995 5696
rect 1922 5697 1923 5698
rect 1946 5697 1947 5698
rect 1910 5699 1911 5700
rect 1922 5699 1923 5700
rect 1898 5701 1899 5702
rect 1910 5701 1911 5702
rect 1417 5703 1418 5704
rect 1898 5703 1899 5704
rect 2033 5703 2034 5704
rect 2240 5703 2241 5704
rect 2042 5705 2043 5706
rect 2072 5705 2073 5706
rect 2030 5707 2031 5708
rect 2042 5707 2043 5708
rect 2120 5707 2121 5708
rect 3454 5707 3455 5708
rect 2090 5709 2091 5710
rect 2120 5709 2121 5710
rect 2054 5711 2055 5712
rect 2090 5711 2091 5712
rect 2036 5713 2037 5714
rect 2054 5713 2055 5714
rect 2036 5715 2037 5716
rect 2060 5715 2061 5716
rect 2012 5717 2013 5718
rect 2060 5717 2061 5718
rect 2012 5719 2013 5720
rect 2018 5719 2019 5720
rect 1970 5721 1971 5722
rect 2018 5721 2019 5722
rect 1489 5723 1490 5724
rect 1970 5723 1971 5724
rect 2234 5723 2235 5724
rect 2282 5723 2283 5724
rect 2228 5725 2229 5726
rect 2282 5725 2283 5726
rect 2186 5727 2187 5728
rect 2228 5727 2229 5728
rect 2240 5727 2241 5728
rect 2252 5727 2253 5728
rect 2246 5729 2247 5730
rect 2270 5729 2271 5730
rect 2252 5731 2253 5732
rect 2258 5731 2259 5732
rect 2258 5733 2259 5734
rect 2264 5733 2265 5734
rect 2264 5735 2265 5736
rect 3361 5735 3362 5736
rect 2270 5737 2271 5738
rect 2294 5737 2295 5738
rect 2276 5739 2277 5740
rect 3327 5739 3328 5740
rect 2276 5741 2277 5742
rect 2288 5741 2289 5742
rect 2198 5743 2199 5744
rect 2288 5743 2289 5744
rect 2198 5745 2199 5746
rect 2210 5745 2211 5746
rect 2210 5747 2211 5748
rect 2216 5747 2217 5748
rect 2156 5749 2157 5750
rect 2216 5749 2217 5750
rect 2144 5751 2145 5752
rect 2156 5751 2157 5752
rect 2114 5753 2115 5754
rect 2144 5753 2145 5754
rect 2084 5755 2085 5756
rect 2114 5755 2115 5756
rect 1474 5757 1475 5758
rect 2084 5757 2085 5758
rect 1475 5759 1476 5760
rect 2186 5759 2187 5760
rect 2294 5759 2295 5760
rect 2306 5759 2307 5760
rect 2300 5761 2301 5762
rect 3465 5761 3466 5762
rect 2300 5763 2301 5764
rect 2312 5763 2313 5764
rect 2306 5765 2307 5766
rect 2318 5765 2319 5766
rect 2312 5767 2313 5768
rect 2324 5767 2325 5768
rect 2318 5769 2319 5770
rect 2330 5769 2331 5770
rect 2324 5771 2325 5772
rect 2348 5771 2349 5772
rect 2330 5773 2331 5774
rect 2354 5773 2355 5774
rect 2333 5775 2334 5776
rect 2357 5775 2358 5776
rect 2336 5777 2337 5778
rect 3354 5777 3355 5778
rect 2336 5779 2337 5780
rect 2366 5779 2367 5780
rect 2348 5781 2349 5782
rect 2378 5781 2379 5782
rect 2354 5783 2355 5784
rect 2360 5783 2361 5784
rect 2360 5785 2361 5786
rect 2384 5785 2385 5786
rect 2366 5787 2367 5788
rect 2396 5787 2397 5788
rect 2378 5789 2379 5790
rect 2402 5789 2403 5790
rect 2384 5791 2385 5792
rect 3330 5791 3331 5792
rect 2396 5793 2397 5794
rect 2414 5793 2415 5794
rect 2402 5795 2403 5796
rect 2426 5795 2427 5796
rect 2408 5797 2409 5798
rect 2414 5797 2415 5798
rect 2408 5799 2409 5800
rect 3405 5799 3406 5800
rect 2420 5801 2421 5802
rect 3451 5801 3452 5802
rect 2222 5803 2223 5804
rect 3451 5803 3452 5804
rect 2192 5805 2193 5806
rect 2222 5805 2223 5806
rect 1478 5807 1479 5808
rect 2192 5807 2193 5808
rect 2420 5807 2421 5808
rect 2438 5807 2439 5808
rect 2426 5809 2427 5810
rect 2450 5809 2451 5810
rect 2438 5811 2439 5812
rect 2456 5811 2457 5812
rect 2450 5813 2451 5814
rect 2468 5813 2469 5814
rect 2456 5815 2457 5816
rect 2474 5815 2475 5816
rect 2468 5817 2469 5818
rect 3323 5817 3324 5818
rect 2474 5819 2475 5820
rect 2492 5819 2493 5820
rect 2486 5821 2487 5822
rect 3320 5821 3321 5822
rect 2486 5823 2487 5824
rect 3395 5823 3396 5824
rect 2492 5825 2493 5826
rect 2504 5825 2505 5826
rect 2504 5827 2505 5828
rect 2516 5827 2517 5828
rect 2516 5829 2517 5830
rect 2528 5829 2529 5830
rect 2528 5831 2529 5832
rect 2540 5831 2541 5832
rect 2540 5833 2541 5834
rect 2552 5833 2553 5834
rect 2591 5833 2592 5834
rect 2879 5833 2880 5834
rect 2594 5835 2595 5836
rect 2618 5835 2619 5836
rect 2606 5837 2607 5838
rect 2618 5837 2619 5838
rect 2606 5839 2607 5840
rect 2648 5839 2649 5840
rect 2648 5841 2649 5842
rect 2666 5841 2667 5842
rect 2672 5841 2673 5842
rect 2678 5841 2679 5842
rect 2678 5843 2679 5844
rect 2684 5843 2685 5844
rect 2684 5845 2685 5846
rect 2690 5845 2691 5846
rect 2690 5847 2691 5848
rect 2702 5847 2703 5848
rect 2696 5849 2697 5850
rect 3365 5849 3366 5850
rect 2696 5851 2697 5852
rect 2708 5851 2709 5852
rect 2702 5853 2703 5854
rect 2714 5853 2715 5854
rect 2708 5855 2709 5856
rect 2720 5855 2721 5856
rect 2714 5857 2715 5858
rect 3468 5857 3469 5858
rect 2720 5859 2721 5860
rect 2726 5859 2727 5860
rect 2726 5861 2727 5862
rect 3407 5861 3408 5862
rect 2756 5863 2757 5864
rect 2762 5863 2763 5864
rect 2762 5865 2763 5866
rect 2774 5865 2775 5866
rect 2768 5867 2769 5868
rect 2822 5867 2823 5868
rect 2774 5869 2775 5870
rect 3403 5869 3404 5870
rect 2780 5871 2781 5872
rect 3447 5871 3448 5872
rect 2432 5873 2433 5874
rect 3448 5873 3449 5874
rect 2432 5875 2433 5876
rect 2444 5875 2445 5876
rect 2444 5877 2445 5878
rect 2462 5877 2463 5878
rect 2462 5879 2463 5880
rect 2480 5879 2481 5880
rect 2480 5881 2481 5882
rect 2498 5881 2499 5882
rect 2498 5883 2499 5884
rect 2510 5883 2511 5884
rect 2510 5885 2511 5886
rect 2522 5885 2523 5886
rect 2522 5887 2523 5888
rect 2534 5887 2535 5888
rect 2534 5889 2535 5890
rect 2546 5889 2547 5890
rect 2546 5891 2547 5892
rect 2558 5891 2559 5892
rect 2558 5893 2559 5894
rect 2564 5893 2565 5894
rect 2564 5895 2565 5896
rect 2570 5895 2571 5896
rect 2570 5897 2571 5898
rect 2576 5897 2577 5898
rect 1516 5899 1517 5900
rect 2576 5899 2577 5900
rect 2786 5899 2787 5900
rect 3429 5899 3430 5900
rect 2786 5901 2787 5902
rect 2798 5901 2799 5902
rect 2792 5903 2793 5904
rect 3444 5903 3445 5904
rect 2792 5905 2793 5906
rect 2804 5905 2805 5906
rect 1512 5907 1513 5908
rect 2804 5907 2805 5908
rect 1513 5909 1514 5910
rect 1904 5909 1905 5910
rect 1904 5911 1905 5912
rect 1934 5911 1935 5912
rect 1916 5913 1917 5914
rect 1934 5913 1935 5914
rect 1892 5915 1893 5916
rect 1916 5915 1917 5916
rect 1491 5917 1492 5918
rect 1892 5917 1893 5918
rect 1492 5919 1493 5920
rect 2600 5919 2601 5920
rect 2600 5921 2601 5922
rect 2612 5921 2613 5922
rect 2612 5923 2613 5924
rect 2624 5923 2625 5924
rect 2624 5925 2625 5926
rect 2660 5925 2661 5926
rect 1538 5927 1539 5928
rect 2660 5927 2661 5928
rect 2798 5927 2799 5928
rect 2816 5927 2817 5928
rect 2801 5929 2802 5930
rect 3023 5929 3024 5930
rect 2807 5931 2808 5932
rect 2825 5931 2826 5932
rect 2810 5933 2811 5934
rect 3400 5933 3401 5934
rect 2810 5935 2811 5936
rect 2828 5935 2829 5936
rect 2816 5937 2817 5938
rect 2834 5937 2835 5938
rect 2822 5939 2823 5940
rect 2840 5939 2841 5940
rect 2828 5941 2829 5942
rect 2846 5941 2847 5942
rect 2834 5943 2835 5944
rect 2852 5943 2853 5944
rect 2840 5945 2841 5946
rect 2858 5945 2859 5946
rect 2846 5947 2847 5948
rect 2864 5947 2865 5948
rect 2852 5949 2853 5950
rect 2870 5949 2871 5950
rect 2858 5951 2859 5952
rect 3026 5951 3027 5952
rect 2864 5953 2865 5954
rect 2882 5953 2883 5954
rect 2870 5955 2871 5956
rect 2888 5955 2889 5956
rect 2876 5957 2877 5958
rect 2894 5957 2895 5958
rect 2882 5959 2883 5960
rect 2900 5959 2901 5960
rect 2888 5961 2889 5962
rect 2963 5961 2964 5962
rect 2900 5963 2901 5964
rect 2912 5963 2913 5964
rect 2906 5965 2907 5966
rect 3351 5965 3352 5966
rect 2912 5967 2913 5968
rect 2918 5967 2919 5968
rect 2918 5969 2919 5970
rect 2924 5969 2925 5970
rect 2924 5971 2925 5972
rect 2930 5971 2931 5972
rect 2930 5973 2931 5974
rect 2936 5973 2937 5974
rect 2936 5975 2937 5976
rect 2942 5975 2943 5976
rect 2942 5977 2943 5978
rect 2972 5977 2973 5978
rect 2948 5979 2949 5980
rect 3444 5979 3445 5980
rect 2948 5981 2949 5982
rect 2954 5981 2955 5982
rect 2954 5983 2955 5984
rect 2960 5983 2961 5984
rect 2960 5985 2961 5986
rect 2966 5985 2967 5986
rect 2966 5987 2967 5988
rect 3032 5987 3033 5988
rect 2972 5989 2973 5990
rect 2978 5989 2979 5990
rect 2975 5991 2976 5992
rect 2981 5991 2982 5992
rect 2978 5993 2979 5994
rect 2984 5993 2985 5994
rect 2984 5995 2985 5996
rect 2990 5995 2991 5996
rect 2990 5997 2991 5998
rect 3393 5997 3394 5998
rect 2996 5999 2997 6000
rect 3044 5999 3045 6000
rect 3011 6001 3012 6002
rect 3035 6001 3036 6002
rect 3020 6003 3021 6004
rect 3062 6003 3063 6004
rect 3026 6005 3027 6006
rect 3068 6005 3069 6006
rect 3044 6007 3045 6008
rect 3074 6007 3075 6008
rect 3062 6009 3063 6010
rect 3110 6009 3111 6010
rect 3068 6011 3069 6012
rect 3095 6011 3096 6012
rect 3074 6013 3075 6014
rect 3092 6013 3093 6014
rect 3086 6015 3087 6016
rect 3128 6015 3129 6016
rect 3092 6017 3093 6018
rect 3116 6017 3117 6018
rect 3098 6019 3099 6020
rect 3134 6019 3135 6020
rect 3104 6021 3105 6022
rect 3110 6021 3111 6022
rect 3104 6023 3105 6024
rect 3140 6023 3141 6024
rect 3107 6025 3108 6026
rect 3113 6025 3114 6026
rect 3134 6025 3135 6026
rect 3182 6025 3183 6026
rect 3140 6027 3141 6028
rect 3188 6027 3189 6028
rect 3152 6029 3153 6030
rect 3422 6029 3423 6030
rect 2126 6031 2127 6032
rect 3423 6031 3424 6032
rect 2096 6033 2097 6034
rect 2126 6033 2127 6034
rect 2096 6035 2097 6036
rect 2150 6035 2151 6036
rect 2138 6037 2139 6038
rect 2150 6037 2151 6038
rect 2138 6039 2139 6040
rect 2162 6039 2163 6040
rect 2162 6041 2163 6042
rect 2168 6041 2169 6042
rect 2168 6043 2169 6044
rect 2174 6043 2175 6044
rect 1447 6045 1448 6046
rect 2174 6045 2175 6046
rect 1448 6047 1449 6048
rect 2552 6047 2553 6048
rect 3146 6047 3147 6048
rect 3152 6047 3153 6048
rect 3146 6049 3147 6050
rect 3194 6049 3195 6050
rect 3158 6051 3159 6052
rect 3402 6051 3403 6052
rect 3158 6053 3159 6054
rect 3206 6053 3207 6054
rect 3164 6055 3165 6056
rect 3282 6055 3283 6056
rect 3164 6057 3165 6058
rect 3200 6057 3201 6058
rect 3176 6059 3177 6060
rect 3224 6059 3225 6060
rect 3182 6061 3183 6062
rect 3230 6061 3231 6062
rect 3188 6063 3189 6064
rect 3430 6063 3431 6064
rect 3200 6065 3201 6066
rect 3248 6065 3249 6066
rect 3203 6067 3204 6068
rect 3251 6067 3252 6068
rect 3206 6069 3207 6070
rect 3218 6069 3219 6070
rect 3209 6071 3210 6072
rect 3221 6071 3222 6072
rect 3218 6073 3219 6074
rect 3260 6073 3261 6074
rect 3221 6075 3222 6076
rect 3263 6075 3264 6076
rect 3224 6077 3225 6078
rect 3266 6077 3267 6078
rect 3230 6079 3231 6080
rect 3272 6079 3273 6080
rect 2588 6081 2589 6082
rect 3272 6081 3273 6082
rect 2588 6083 2589 6084
rect 2732 6083 2733 6084
rect 2732 6085 2733 6086
rect 2738 6085 2739 6086
rect 2738 6087 2739 6088
rect 2744 6087 2745 6088
rect 2744 6089 2745 6090
rect 2750 6089 2751 6090
rect 3233 6089 3234 6090
rect 3275 6089 3276 6090
rect 1640 6091 1641 6092
rect 3275 6091 3276 6092
rect 1634 6093 1635 6094
rect 1640 6093 1641 6094
rect 3242 6093 3243 6094
rect 3284 6093 3285 6094
rect 3248 6095 3249 6096
rect 3290 6095 3291 6096
rect 3260 6097 3261 6098
rect 3308 6097 3309 6098
rect 3263 6099 3264 6100
rect 3311 6099 3312 6100
rect 3266 6101 3267 6102
rect 3314 6101 3315 6102
rect 3285 6103 3286 6104
rect 3333 6103 3334 6104
rect 3291 6105 3292 6106
rect 3339 6105 3340 6106
rect 2030 6107 2031 6108
rect 3339 6107 3340 6108
rect 3296 6109 3297 6110
rect 3398 6109 3399 6110
rect 3309 6111 3310 6112
rect 3357 6111 3358 6112
rect 2066 6113 2067 6114
rect 3358 6113 3359 6114
rect 3315 6115 3316 6116
rect 3384 6115 3385 6116
rect 3321 6117 3322 6118
rect 3369 6117 3370 6118
rect 2666 6119 2667 6120
rect 3368 6119 3369 6120
rect 3324 6121 3325 6122
rect 3372 6121 3373 6122
rect 3342 6123 3343 6124
rect 3381 6123 3382 6124
rect 3345 6125 3346 6126
rect 3387 6125 3388 6126
rect 3348 6127 3349 6128
rect 3390 6127 3391 6128
rect 3371 6129 3372 6130
rect 3413 6129 3414 6130
rect 3374 6131 3375 6132
rect 3416 6131 3417 6132
rect 3377 6133 3378 6134
rect 3434 6133 3435 6134
rect 3389 6135 3390 6136
rect 3419 6135 3420 6136
rect 2342 6137 2343 6138
rect 3420 6137 3421 6138
rect 2342 6139 2343 6140
rect 2372 6139 2373 6140
rect 2372 6141 2373 6142
rect 3426 6141 3427 6142
rect 3236 6143 3237 6144
rect 3427 6143 3428 6144
rect 3236 6145 3237 6146
rect 3278 6145 3279 6146
rect 3116 6147 3117 6148
rect 3279 6147 3280 6148
rect 3410 6147 3411 6148
rect 3458 6147 3459 6148
rect 3414 6149 3415 6150
rect 3438 6149 3439 6150
rect 3392 6151 3393 6152
rect 3437 6151 3438 6152
rect 3417 6153 3418 6154
rect 3441 6153 3442 6154
rect 3014 6155 3015 6156
rect 3441 6155 3442 6156
rect 3014 6157 3015 6158
rect 3038 6157 3039 6158
rect 3038 6159 3039 6160
rect 3050 6159 3051 6160
rect 3050 6161 3051 6162
rect 3056 6161 3057 6162
rect 3056 6163 3057 6164
rect 3080 6163 3081 6164
rect 3080 6165 3081 6166
rect 3122 6165 3123 6166
rect 3122 6167 3123 6168
rect 3170 6167 3171 6168
rect 3170 6169 3171 6170
rect 3212 6169 3213 6170
rect 1417 6178 1418 6179
rect 1850 6178 1851 6179
rect 1417 6180 1418 6181
rect 1513 6180 1514 6181
rect 1420 6182 1421 6183
rect 2186 6182 2187 6183
rect 1420 6184 1421 6185
rect 1668 6184 1669 6185
rect 1424 6186 1425 6187
rect 1812 6186 1813 6187
rect 1424 6188 1425 6189
rect 1604 6188 1605 6189
rect 1427 6190 1428 6191
rect 1482 6190 1483 6191
rect 1427 6192 1428 6193
rect 1598 6192 1599 6193
rect 1431 6194 1432 6195
rect 1674 6194 1675 6195
rect 1431 6196 1432 6197
rect 1692 6196 1693 6197
rect 1434 6198 1435 6199
rect 1730 6198 1731 6199
rect 1434 6200 1435 6201
rect 1441 6200 1442 6201
rect 1438 6202 1439 6203
rect 2166 6202 2167 6203
rect 1438 6204 1439 6205
rect 1686 6204 1687 6205
rect 1441 6206 1442 6207
rect 1742 6206 1743 6207
rect 1448 6208 1449 6209
rect 2288 6208 2289 6209
rect 1448 6210 1449 6211
rect 2844 6210 2845 6211
rect 1457 6212 1458 6213
rect 1475 6212 1476 6213
rect 1457 6214 1458 6215
rect 1463 6214 1464 6215
rect 1463 6216 1464 6217
rect 1469 6216 1470 6217
rect 1469 6218 1470 6219
rect 2807 6218 2808 6219
rect 1472 6220 1473 6221
rect 2636 6220 2637 6221
rect 1476 6222 1477 6223
rect 1746 6222 1747 6223
rect 1478 6224 1479 6225
rect 2438 6224 2439 6225
rect 1479 6226 1480 6227
rect 1628 6226 1629 6227
rect 1485 6228 1486 6229
rect 2522 6228 2523 6229
rect 1489 6230 1490 6231
rect 2546 6230 2547 6231
rect 1492 6232 1493 6233
rect 1766 6232 1767 6233
rect 1494 6234 1495 6235
rect 1501 6234 1502 6235
rect 1500 6236 1501 6237
rect 1644 6236 1645 6237
rect 1503 6238 1504 6239
rect 1700 6238 1701 6239
rect 1512 6240 1513 6241
rect 1547 6240 1548 6241
rect 1516 6242 1517 6243
rect 1889 6242 1890 6243
rect 1515 6244 1516 6245
rect 2180 6244 2181 6245
rect 1518 6246 1519 6247
rect 1550 6246 1551 6247
rect 1525 6248 1526 6249
rect 1676 6248 1677 6249
rect 1524 6250 1525 6251
rect 1556 6250 1557 6251
rect 1528 6252 1529 6253
rect 2096 6252 2097 6253
rect 1532 6254 1533 6255
rect 3011 6254 3012 6255
rect 1539 6256 1540 6257
rect 1770 6256 1771 6257
rect 1542 6258 1543 6259
rect 1580 6258 1581 6259
rect 1554 6260 1555 6261
rect 1592 6260 1593 6261
rect 1560 6262 1561 6263
rect 1610 6262 1611 6263
rect 1566 6264 1567 6265
rect 1616 6264 1617 6265
rect 1572 6266 1573 6267
rect 1622 6266 1623 6267
rect 1584 6268 1585 6269
rect 2726 6268 2727 6269
rect 1587 6270 1588 6271
rect 2804 6270 2805 6271
rect 1596 6272 1597 6273
rect 1646 6272 1647 6273
rect 1608 6274 1609 6275
rect 2648 6274 2649 6275
rect 1611 6276 1612 6277
rect 2340 6276 2341 6277
rect 1614 6278 1615 6279
rect 1664 6278 1665 6279
rect 1620 6280 1621 6281
rect 1682 6280 1683 6281
rect 1626 6282 1627 6283
rect 1688 6282 1689 6283
rect 1632 6284 1633 6285
rect 1694 6284 1695 6285
rect 1652 6286 1653 6287
rect 2033 6286 2034 6287
rect 1656 6288 1657 6289
rect 1712 6288 1713 6289
rect 1662 6290 1663 6291
rect 1724 6290 1725 6291
rect 1680 6292 1681 6293
rect 1736 6292 1737 6293
rect 1698 6294 1699 6295
rect 1718 6294 1719 6295
rect 1710 6296 1711 6297
rect 1754 6296 1755 6297
rect 1716 6298 1717 6299
rect 1796 6298 1797 6299
rect 1722 6300 1723 6301
rect 1790 6300 1791 6301
rect 1728 6302 1729 6303
rect 2564 6302 2565 6303
rect 1734 6304 1735 6305
rect 1760 6304 1761 6305
rect 1740 6306 1741 6307
rect 2474 6306 2475 6307
rect 1752 6308 1753 6309
rect 2456 6308 2457 6309
rect 1758 6310 1759 6311
rect 1772 6310 1773 6311
rect 1764 6312 1765 6313
rect 1778 6312 1779 6313
rect 1776 6314 1777 6315
rect 2360 6314 2361 6315
rect 1782 6316 1783 6317
rect 1784 6316 1785 6317
rect 1788 6316 1789 6317
rect 2462 6316 2463 6317
rect 1794 6318 1795 6319
rect 2588 6318 2589 6319
rect 1800 6320 1801 6321
rect 1868 6320 1869 6321
rect 1802 6322 1803 6323
rect 1836 6322 1837 6323
rect 1806 6324 1807 6325
rect 1808 6324 1809 6325
rect 1814 6324 1815 6325
rect 1818 6324 1819 6325
rect 1820 6324 1821 6325
rect 1842 6324 1843 6325
rect 1824 6326 1825 6327
rect 2292 6326 2293 6327
rect 1826 6328 1827 6329
rect 1848 6328 1849 6329
rect 1827 6330 1828 6331
rect 2540 6330 2541 6331
rect 1829 6332 1830 6333
rect 1851 6332 1852 6333
rect 1830 6334 1831 6335
rect 1832 6334 1833 6335
rect 1838 6334 1839 6335
rect 1854 6334 1855 6335
rect 1844 6336 1845 6337
rect 1890 6336 1891 6337
rect 1856 6338 1857 6339
rect 1878 6338 1879 6339
rect 1860 6340 1861 6341
rect 2798 6340 2799 6341
rect 1862 6342 1863 6343
rect 1884 6342 1885 6343
rect 1866 6344 1867 6345
rect 2216 6344 2217 6345
rect 1872 6346 1873 6347
rect 2222 6346 2223 6347
rect 1874 6348 1875 6349
rect 2016 6348 2017 6349
rect 1880 6350 1881 6351
rect 2088 6350 2089 6351
rect 1886 6352 1887 6353
rect 3451 6352 3452 6353
rect 1568 6354 1569 6355
rect 1887 6354 1888 6355
rect 1892 6354 1893 6355
rect 1950 6354 1951 6355
rect 1896 6356 1897 6357
rect 1916 6356 1917 6357
rect 1898 6358 1899 6359
rect 1908 6358 1909 6359
rect 1902 6360 1903 6361
rect 1910 6360 1911 6361
rect 1904 6362 1905 6363
rect 1938 6362 1939 6363
rect 1905 6364 1906 6365
rect 1919 6364 1920 6365
rect 1914 6366 1915 6367
rect 1940 6366 1941 6367
rect 1920 6368 1921 6369
rect 1922 6368 1923 6369
rect 1928 6368 1929 6369
rect 2082 6368 2083 6369
rect 1932 6370 1933 6371
rect 1934 6370 1935 6371
rect 1944 6370 1945 6371
rect 1946 6370 1947 6371
rect 1956 6370 1957 6371
rect 1958 6370 1959 6371
rect 1962 6370 1963 6371
rect 1970 6370 1971 6371
rect 1964 6372 1965 6373
rect 1980 6372 1981 6373
rect 1974 6374 1975 6375
rect 1994 6374 1995 6375
rect 1976 6376 1977 6377
rect 2064 6376 2065 6377
rect 1982 6378 1983 6379
rect 1992 6378 1993 6379
rect 1986 6380 1987 6381
rect 2000 6380 2001 6381
rect 1998 6382 1999 6383
rect 2018 6382 2019 6383
rect 1925 6384 1926 6385
rect 2019 6384 2020 6385
rect 1445 6386 1446 6387
rect 1926 6386 1927 6387
rect 1445 6388 1446 6389
rect 1952 6388 1953 6389
rect 2004 6388 2005 6389
rect 2006 6388 2007 6389
rect 2010 6388 2011 6389
rect 2012 6388 2013 6389
rect 2022 6388 2023 6389
rect 2024 6388 2025 6389
rect 2028 6388 2029 6389
rect 2048 6388 2049 6389
rect 2030 6390 2031 6391
rect 2234 6390 2235 6391
rect 2034 6392 2035 6393
rect 2072 6392 2073 6393
rect 2036 6394 2037 6395
rect 2070 6394 2071 6395
rect 2040 6396 2041 6397
rect 2060 6396 2061 6397
rect 2042 6398 2043 6399
rect 2052 6398 2053 6399
rect 2046 6400 2047 6401
rect 2054 6400 2055 6401
rect 2058 6400 2059 6401
rect 3361 6400 3362 6401
rect 2066 6402 2067 6403
rect 3402 6402 3403 6403
rect 2076 6404 2077 6405
rect 2090 6404 2091 6405
rect 1967 6406 1968 6407
rect 2091 6406 2092 6407
rect 1968 6408 1969 6409
rect 1988 6408 1989 6409
rect 2078 6408 2079 6409
rect 3227 6408 3228 6409
rect 2084 6410 2085 6411
rect 2160 6410 2161 6411
rect 2094 6412 2095 6413
rect 2102 6412 2103 6413
rect 2100 6414 2101 6415
rect 2108 6414 2109 6415
rect 2106 6416 2107 6417
rect 2114 6416 2115 6417
rect 2112 6418 2113 6419
rect 2126 6418 2127 6419
rect 2118 6420 2119 6421
rect 2144 6420 2145 6421
rect 2120 6422 2121 6423
rect 3289 6422 3290 6423
rect 2124 6424 2125 6425
rect 3423 6424 3424 6425
rect 2130 6426 2131 6427
rect 2132 6426 2133 6427
rect 2136 6426 2137 6427
rect 2192 6426 2193 6427
rect 2138 6428 2139 6429
rect 2172 6428 2173 6429
rect 2142 6430 2143 6431
rect 2156 6430 2157 6431
rect 2148 6432 2149 6433
rect 2150 6432 2151 6433
rect 2154 6432 2155 6433
rect 2162 6432 2163 6433
rect 2168 6432 2169 6433
rect 2178 6432 2179 6433
rect 2174 6434 2175 6435
rect 2184 6434 2185 6435
rect 2181 6436 2182 6437
rect 2567 6436 2568 6437
rect 2190 6438 2191 6439
rect 2204 6438 2205 6439
rect 2196 6440 2197 6441
rect 2324 6440 2325 6441
rect 2198 6442 2199 6443
rect 2214 6442 2215 6443
rect 2202 6444 2203 6445
rect 2318 6444 2319 6445
rect 2208 6446 2209 6447
rect 2210 6446 2211 6447
rect 2220 6446 2221 6447
rect 2228 6446 2229 6447
rect 2223 6448 2224 6449
rect 2591 6448 2592 6449
rect 2226 6450 2227 6451
rect 2294 6450 2295 6451
rect 2232 6452 2233 6453
rect 2300 6452 2301 6453
rect 2238 6454 2239 6455
rect 2354 6454 2355 6455
rect 2240 6456 2241 6457
rect 2268 6456 2269 6457
rect 2244 6458 2245 6459
rect 2264 6458 2265 6459
rect 2246 6460 2247 6461
rect 2262 6460 2263 6461
rect 2250 6462 2251 6463
rect 2252 6462 2253 6463
rect 2256 6462 2257 6463
rect 2258 6462 2259 6463
rect 2270 6462 2271 6463
rect 2274 6462 2275 6463
rect 2276 6462 2277 6463
rect 2286 6462 2287 6463
rect 2282 6464 2283 6465
rect 2298 6464 2299 6465
rect 2304 6464 2305 6465
rect 2330 6464 2331 6465
rect 2306 6466 2307 6467
rect 2310 6466 2311 6467
rect 2307 6468 2308 6469
rect 2333 6468 2334 6469
rect 2312 6470 2313 6471
rect 2316 6470 2317 6471
rect 2322 6470 2323 6471
rect 2390 6470 2391 6471
rect 2328 6472 2329 6473
rect 3405 6472 3406 6473
rect 2334 6474 2335 6475
rect 2414 6474 2415 6475
rect 2336 6476 2337 6477
rect 2346 6476 2347 6477
rect 2337 6478 2338 6479
rect 2801 6478 2802 6479
rect 2342 6480 2343 6481
rect 3444 6480 3445 6481
rect 2348 6482 2349 6483
rect 2352 6482 2353 6483
rect 2358 6482 2359 6483
rect 2660 6482 2661 6483
rect 2364 6484 2365 6485
rect 2408 6484 2409 6485
rect 2366 6486 2367 6487
rect 2376 6486 2377 6487
rect 2370 6488 2371 6489
rect 2420 6488 2421 6489
rect 2372 6490 2373 6491
rect 2394 6490 2395 6491
rect 2378 6492 2379 6493
rect 2382 6492 2383 6493
rect 2384 6492 2385 6493
rect 3268 6492 3269 6493
rect 2396 6494 2397 6495
rect 2406 6494 2407 6495
rect 2400 6496 2401 6497
rect 2402 6496 2403 6497
rect 2412 6496 2413 6497
rect 3420 6496 3421 6497
rect 2418 6498 2419 6499
rect 3300 6498 3301 6499
rect 2424 6500 2425 6501
rect 2450 6500 2451 6501
rect 2426 6502 2427 6503
rect 2430 6502 2431 6503
rect 1640 6504 1641 6505
rect 2427 6504 2428 6505
rect 2432 6504 2433 6505
rect 2436 6504 2437 6505
rect 2442 6504 2443 6505
rect 2480 6504 2481 6505
rect 2444 6506 2445 6507
rect 2448 6506 2449 6507
rect 2454 6506 2455 6507
rect 2468 6506 2469 6507
rect 2460 6508 2461 6509
rect 2708 6508 2709 6509
rect 2466 6510 2467 6511
rect 2858 6510 2859 6511
rect 2472 6512 2473 6513
rect 2486 6512 2487 6513
rect 2478 6514 2479 6515
rect 2624 6514 2625 6515
rect 2484 6516 2485 6517
rect 2582 6516 2583 6517
rect 2490 6518 2491 6519
rect 2504 6518 2505 6519
rect 2492 6520 2493 6521
rect 3395 6520 3396 6521
rect 2496 6522 2497 6523
rect 2510 6522 2511 6523
rect 2498 6524 2499 6525
rect 3398 6524 3399 6525
rect 2502 6526 2503 6527
rect 2552 6526 2553 6527
rect 2508 6528 2509 6529
rect 2528 6528 2529 6529
rect 2514 6530 2515 6531
rect 2558 6530 2559 6531
rect 2516 6532 2517 6533
rect 2520 6532 2521 6533
rect 2526 6532 2527 6533
rect 2570 6532 2571 6533
rect 2532 6534 2533 6535
rect 2576 6534 2577 6535
rect 2534 6536 2535 6537
rect 3351 6536 3352 6537
rect 2538 6538 2539 6539
rect 3275 6538 3276 6539
rect 2544 6540 2545 6541
rect 2822 6540 2823 6541
rect 2550 6542 2551 6543
rect 2762 6542 2763 6543
rect 2556 6544 2557 6545
rect 2600 6544 2601 6545
rect 2562 6546 2563 6547
rect 3166 6546 3167 6547
rect 2568 6548 2569 6549
rect 2606 6548 2607 6549
rect 2574 6550 2575 6551
rect 2618 6550 2619 6551
rect 2580 6552 2581 6553
rect 2942 6552 2943 6553
rect 2586 6554 2587 6555
rect 2630 6554 2631 6555
rect 2592 6556 2593 6557
rect 2642 6556 2643 6557
rect 2594 6558 2595 6559
rect 3156 6558 3157 6559
rect 2598 6560 2599 6561
rect 2654 6560 2655 6561
rect 2604 6562 2605 6563
rect 2666 6562 2667 6563
rect 2610 6564 2611 6565
rect 2702 6564 2703 6565
rect 2616 6566 2617 6567
rect 2672 6566 2673 6567
rect 2622 6568 2623 6569
rect 2678 6568 2679 6569
rect 2628 6570 2629 6571
rect 2684 6570 2685 6571
rect 2634 6572 2635 6573
rect 2690 6572 2691 6573
rect 2640 6574 2641 6575
rect 3358 6574 3359 6575
rect 2646 6576 2647 6577
rect 2696 6576 2697 6577
rect 2652 6578 2653 6579
rect 3365 6578 3366 6579
rect 2658 6580 2659 6581
rect 3368 6580 3369 6581
rect 2664 6582 2665 6583
rect 2714 6582 2715 6583
rect 2670 6584 2671 6585
rect 2720 6584 2721 6585
rect 2676 6586 2677 6587
rect 2732 6586 2733 6587
rect 2682 6588 2683 6589
rect 2738 6588 2739 6589
rect 2688 6590 2689 6591
rect 2744 6590 2745 6591
rect 2706 6592 2707 6593
rect 2774 6592 2775 6593
rect 2712 6594 2713 6595
rect 2864 6594 2865 6595
rect 2718 6596 2719 6597
rect 2870 6596 2871 6597
rect 2724 6598 2725 6599
rect 2786 6598 2787 6599
rect 2730 6600 2731 6601
rect 2792 6600 2793 6601
rect 2736 6602 2737 6603
rect 2810 6602 2811 6603
rect 2742 6604 2743 6605
rect 2816 6604 2817 6605
rect 2748 6606 2749 6607
rect 2828 6606 2829 6607
rect 2754 6608 2755 6609
rect 2834 6608 2835 6609
rect 2766 6610 2767 6611
rect 2840 6610 2841 6611
rect 2772 6612 2773 6613
rect 2846 6612 2847 6613
rect 2778 6614 2779 6615
rect 2900 6614 2901 6615
rect 2784 6616 2785 6617
rect 2906 6616 2907 6617
rect 2790 6618 2791 6619
rect 2912 6618 2913 6619
rect 1535 6620 1536 6621
rect 2913 6620 2914 6621
rect 1536 6622 1537 6623
rect 2768 6622 2769 6623
rect 2796 6622 2797 6623
rect 2876 6622 2877 6623
rect 2802 6624 2803 6625
rect 2882 6624 2883 6625
rect 2808 6626 2809 6627
rect 2888 6626 2889 6627
rect 2820 6628 2821 6629
rect 2918 6628 2919 6629
rect 2826 6630 2827 6631
rect 2924 6630 2925 6631
rect 2832 6632 2833 6633
rect 2930 6632 2931 6633
rect 2838 6634 2839 6635
rect 2936 6634 2937 6635
rect 2850 6636 2851 6637
rect 2948 6636 2949 6637
rect 2856 6638 2857 6639
rect 2954 6638 2955 6639
rect 2859 6640 2860 6641
rect 2957 6640 2958 6641
rect 2862 6642 2863 6643
rect 2960 6642 2961 6643
rect 2868 6644 2869 6645
rect 2966 6644 2967 6645
rect 2874 6646 2875 6647
rect 2972 6646 2973 6647
rect 2877 6648 2878 6649
rect 3296 6648 3297 6649
rect 2880 6650 2881 6651
rect 2978 6650 2979 6651
rect 2886 6652 2887 6653
rect 2990 6652 2991 6653
rect 2892 6654 2893 6655
rect 3002 6654 3003 6655
rect 2898 6656 2899 6657
rect 2996 6656 2997 6657
rect 2904 6658 2905 6659
rect 3014 6658 3015 6659
rect 1748 6660 1749 6661
rect 3015 6660 3016 6661
rect 2910 6662 2911 6663
rect 3008 6662 3009 6663
rect 2916 6664 2917 6665
rect 3020 6664 3021 6665
rect 2922 6666 2923 6667
rect 3026 6666 3027 6667
rect 2928 6668 2929 6669
rect 3441 6668 3442 6669
rect 2940 6670 2941 6671
rect 3044 6670 3045 6671
rect 2946 6672 2947 6673
rect 3056 6672 3057 6673
rect 2952 6674 2953 6675
rect 3050 6674 3051 6675
rect 2958 6676 2959 6677
rect 3038 6676 3039 6677
rect 2964 6678 2965 6679
rect 3068 6678 3069 6679
rect 2970 6680 2971 6681
rect 3074 6680 3075 6681
rect 2975 6682 2976 6683
rect 3293 6682 3294 6683
rect 2976 6684 2977 6685
rect 3062 6684 3063 6685
rect 2982 6686 2983 6687
rect 3080 6686 3081 6687
rect 2988 6688 2989 6689
rect 3086 6688 3087 6689
rect 2994 6690 2995 6691
rect 3092 6690 3093 6691
rect 3000 6692 3001 6693
rect 3098 6692 3099 6693
rect 3006 6694 3007 6695
rect 3104 6694 3105 6695
rect 3012 6696 3013 6697
rect 3110 6696 3111 6697
rect 3018 6698 3019 6699
rect 3116 6698 3117 6699
rect 2852 6700 2853 6701
rect 3117 6700 3118 6701
rect 3024 6702 3025 6703
rect 3122 6702 3123 6703
rect 3036 6704 3037 6705
rect 3239 6704 3240 6705
rect 3048 6706 3049 6707
rect 3134 6706 3135 6707
rect 3054 6708 3055 6709
rect 3152 6708 3153 6709
rect 3060 6710 3061 6711
rect 3164 6710 3165 6711
rect 3066 6712 3067 6713
rect 3170 6712 3171 6713
rect 3078 6714 3079 6715
rect 3206 6714 3207 6715
rect 3081 6716 3082 6717
rect 3209 6716 3210 6717
rect 3090 6718 3091 6719
rect 3176 6718 3177 6719
rect 3102 6720 3103 6721
rect 3188 6720 3189 6721
rect 3105 6722 3106 6723
rect 3182 6722 3183 6723
rect 3108 6724 3109 6725
rect 3218 6724 3219 6725
rect 3111 6726 3112 6727
rect 3221 6726 3222 6727
rect 3113 6728 3114 6729
rect 3354 6728 3355 6729
rect 3114 6730 3115 6731
rect 3224 6730 3225 6731
rect 2780 6732 2781 6733
rect 3224 6732 3225 6733
rect 3120 6734 3121 6735
rect 3230 6734 3231 6735
rect 3123 6736 3124 6737
rect 3233 6736 3234 6737
rect 3126 6738 3127 6739
rect 3236 6738 3237 6739
rect 3030 6740 3031 6741
rect 3236 6740 3237 6741
rect 3132 6742 3133 6743
rect 3248 6742 3249 6743
rect 3140 6744 3141 6745
rect 3279 6744 3280 6745
rect 3144 6746 3145 6747
rect 3260 6746 3261 6747
rect 2756 6748 2757 6749
rect 3261 6748 3262 6749
rect 3146 6750 3147 6751
rect 3282 6750 3283 6751
rect 3147 6752 3148 6753
rect 3263 6752 3264 6753
rect 2700 6754 2701 6755
rect 3264 6754 3265 6755
rect 3150 6756 3151 6757
rect 3266 6756 3267 6757
rect 3158 6758 3159 6759
rect 3233 6758 3234 6759
rect 2984 6760 2985 6761
rect 3159 6760 3160 6761
rect 3163 6760 3164 6761
rect 3303 6760 3304 6761
rect 3169 6762 3170 6763
rect 3285 6762 3286 6763
rect 2280 6764 2281 6765
rect 3286 6764 3287 6765
rect 3181 6766 3182 6767
rect 3309 6766 3310 6767
rect 3187 6768 3188 6769
rect 3315 6768 3316 6769
rect 3193 6770 3194 6771
rect 3321 6770 3322 6771
rect 3196 6772 3197 6773
rect 3324 6772 3325 6773
rect 3200 6774 3201 6775
rect 3430 6774 3431 6775
rect 1544 6776 1545 6777
rect 3199 6776 3200 6777
rect 3203 6776 3204 6777
rect 3427 6776 3428 6777
rect 2612 6778 2613 6779
rect 3202 6778 3203 6779
rect 3211 6778 3212 6779
rect 3339 6778 3340 6779
rect 3214 6780 3215 6781
rect 3342 6780 3343 6781
rect 3217 6782 3218 6783
rect 3348 6782 3349 6783
rect 3220 6784 3221 6785
rect 3345 6784 3346 6785
rect 3230 6786 3231 6787
rect 3371 6786 3372 6787
rect 3242 6788 3243 6789
rect 3272 6788 3273 6789
rect 2388 6790 2389 6791
rect 3271 6790 3272 6791
rect 3243 6792 3244 6793
rect 3291 6792 3292 6793
rect 3246 6794 3247 6795
rect 3374 6794 3375 6795
rect 3255 6796 3256 6797
rect 3392 6796 3393 6797
rect 3258 6798 3259 6799
rect 3377 6798 3378 6799
rect 3280 6800 3281 6801
rect 3414 6800 3415 6801
rect 3283 6802 3284 6803
rect 3417 6802 3418 6803
rect 3389 6804 3390 6805
rect 3437 6804 3438 6805
rect 3434 6806 3435 6807
rect 3448 6806 3449 6807
rect 1427 6815 1428 6816
rect 1554 6815 1555 6816
rect 1434 6817 1435 6818
rect 1530 6817 1531 6818
rect 1438 6819 1439 6820
rect 1668 6819 1669 6820
rect 1441 6821 1442 6822
rect 1662 6821 1663 6822
rect 1445 6823 1446 6824
rect 2064 6823 2065 6824
rect 1448 6825 1449 6826
rect 1851 6825 1852 6826
rect 1454 6827 1455 6828
rect 1914 6827 1915 6828
rect 1472 6829 1473 6830
rect 1920 6829 1921 6830
rect 1476 6831 1477 6832
rect 2166 6831 2167 6832
rect 1417 6833 1418 6834
rect 1475 6833 1476 6834
rect 1479 6833 1480 6834
rect 2226 6833 2227 6834
rect 1478 6835 1479 6836
rect 2160 6835 2161 6836
rect 1482 6837 1483 6838
rect 2490 6837 2491 6838
rect 1503 6839 1504 6840
rect 1614 6839 1615 6840
rect 1512 6841 1513 6842
rect 2154 6841 2155 6842
rect 1512 6843 1513 6844
rect 2223 6843 2224 6844
rect 1536 6845 1537 6846
rect 2010 6845 2011 6846
rect 1524 6847 1525 6848
rect 1536 6847 1537 6848
rect 1518 6849 1519 6850
rect 1524 6849 1525 6850
rect 1542 6849 1543 6850
rect 1554 6849 1555 6850
rect 1548 6851 1549 6852
rect 2496 6851 2497 6852
rect 1551 6853 1552 6854
rect 1992 6853 1993 6854
rect 1566 6855 1567 6856
rect 1578 6855 1579 6856
rect 1424 6857 1425 6858
rect 1566 6857 1567 6858
rect 1599 6857 1600 6858
rect 2106 6857 2107 6858
rect 1608 6859 1609 6860
rect 1611 6859 1612 6860
rect 1596 6861 1597 6862
rect 1608 6861 1609 6862
rect 1596 6863 1597 6864
rect 1956 6863 1957 6864
rect 1469 6865 1470 6866
rect 1956 6865 1957 6866
rect 1463 6867 1464 6868
rect 1469 6867 1470 6868
rect 1457 6869 1458 6870
rect 1463 6869 1464 6870
rect 1620 6869 1621 6870
rect 1638 6869 1639 6870
rect 1620 6871 1621 6872
rect 2790 6871 2791 6872
rect 1623 6873 1624 6874
rect 2094 6873 2095 6874
rect 1632 6875 1633 6876
rect 1650 6875 1651 6876
rect 1644 6877 1645 6878
rect 1662 6877 1663 6878
rect 1626 6879 1627 6880
rect 1644 6879 1645 6880
rect 1500 6881 1501 6882
rect 1626 6881 1627 6882
rect 1494 6883 1495 6884
rect 1500 6883 1501 6884
rect 1698 6883 1699 6884
rect 1704 6883 1705 6884
rect 1692 6885 1693 6886
rect 1698 6885 1699 6886
rect 1431 6887 1432 6888
rect 1692 6887 1693 6888
rect 1430 6889 1431 6890
rect 1764 6889 1765 6890
rect 1749 6891 1750 6892
rect 2484 6891 2485 6892
rect 1764 6893 1765 6894
rect 1770 6893 1771 6894
rect 1433 6895 1434 6896
rect 1770 6895 1771 6896
rect 1836 6895 1837 6896
rect 3327 6895 3328 6896
rect 1836 6897 1837 6898
rect 1872 6897 1873 6898
rect 1740 6899 1741 6900
rect 1872 6899 1873 6900
rect 1423 6901 1424 6902
rect 1740 6901 1741 6902
rect 1866 6901 1867 6902
rect 1914 6901 1915 6902
rect 1806 6903 1807 6904
rect 1866 6903 1867 6904
rect 1788 6905 1789 6906
rect 1806 6905 1807 6906
rect 1776 6907 1777 6908
rect 1788 6907 1789 6908
rect 1758 6909 1759 6910
rect 1776 6909 1777 6910
rect 1746 6911 1747 6912
rect 1758 6911 1759 6912
rect 1887 6911 1888 6912
rect 1959 6911 1960 6912
rect 1905 6913 1906 6914
rect 1971 6913 1972 6914
rect 1656 6915 1657 6916
rect 1905 6915 1906 6916
rect 1920 6915 1921 6916
rect 2442 6915 2443 6916
rect 1950 6917 1951 6918
rect 1992 6917 1993 6918
rect 1878 6919 1879 6920
rect 1950 6919 1951 6920
rect 1728 6921 1729 6922
rect 1878 6921 1879 6922
rect 1728 6923 1729 6924
rect 1734 6923 1735 6924
rect 1426 6925 1427 6926
rect 1734 6925 1735 6926
rect 1980 6925 1981 6926
rect 2010 6925 2011 6926
rect 1938 6927 1939 6928
rect 1980 6927 1981 6928
rect 1884 6929 1885 6930
rect 1938 6929 1939 6930
rect 1884 6931 1885 6932
rect 3202 6931 3203 6932
rect 2001 6933 2002 6934
rect 2019 6933 2020 6934
rect 2025 6933 2026 6934
rect 2307 6933 2308 6934
rect 2034 6935 2035 6936
rect 2106 6935 2107 6936
rect 1962 6937 1963 6938
rect 2034 6937 2035 6938
rect 1902 6939 1903 6940
rect 1962 6939 1963 6940
rect 1848 6941 1849 6942
rect 1902 6941 1903 6942
rect 1812 6943 1813 6944
rect 1848 6943 1849 6944
rect 1800 6945 1801 6946
rect 1812 6945 1813 6946
rect 1800 6947 1801 6948
rect 3156 6947 3157 6948
rect 2043 6949 2044 6950
rect 2091 6949 2092 6950
rect 2058 6951 2059 6952
rect 2154 6951 2155 6952
rect 1974 6953 1975 6954
rect 2058 6953 2059 6954
rect 1974 6955 1975 6956
rect 2016 6955 2017 6956
rect 1944 6957 1945 6958
rect 2016 6957 2017 6958
rect 1944 6959 1945 6960
rect 2136 6959 2137 6960
rect 2040 6961 2041 6962
rect 2136 6961 2137 6962
rect 2040 6963 2041 6964
rect 2088 6963 2089 6964
rect 2064 6965 2065 6966
rect 3189 6965 3190 6966
rect 2070 6967 2071 6968
rect 2094 6967 2095 6968
rect 1986 6969 1987 6970
rect 2070 6969 2071 6970
rect 1908 6971 1909 6972
rect 1986 6971 1987 6972
rect 1437 6973 1438 6974
rect 1908 6973 1909 6974
rect 2100 6973 2101 6974
rect 2166 6973 2167 6974
rect 2004 6975 2005 6976
rect 2100 6975 2101 6976
rect 1932 6977 1933 6978
rect 2004 6977 2005 6978
rect 1890 6979 1891 6980
rect 1932 6979 1933 6980
rect 1854 6981 1855 6982
rect 1890 6981 1891 6982
rect 1440 6983 1441 6984
rect 1854 6983 1855 6984
rect 2112 6983 2113 6984
rect 3286 6983 3287 6984
rect 2022 6985 2023 6986
rect 2112 6985 2113 6986
rect 1451 6987 1452 6988
rect 2022 6987 2023 6988
rect 2130 6987 2131 6988
rect 2160 6987 2161 6988
rect 2046 6989 2047 6990
rect 2130 6989 2131 6990
rect 1420 6991 1421 6992
rect 2046 6991 2047 6992
rect 2181 6991 2182 6992
rect 2193 6991 2194 6992
rect 2184 6993 2185 6994
rect 2226 6993 2227 6994
rect 1485 6995 1486 6996
rect 2184 6995 2185 6996
rect 2235 6995 2236 6996
rect 3236 6995 3237 6996
rect 2280 6997 2281 6998
rect 3266 6997 3267 6998
rect 2280 6999 2281 7000
rect 2322 6999 2323 7000
rect 2286 7001 2287 7002
rect 2322 7001 2323 7002
rect 2250 7003 2251 7004
rect 2286 7003 2287 7004
rect 2190 7005 2191 7006
rect 2250 7005 2251 7006
rect 2178 7007 2179 7008
rect 2190 7007 2191 7008
rect 2178 7009 2179 7010
rect 3289 7009 3290 7010
rect 2310 7011 2311 7012
rect 3331 7011 3332 7012
rect 2262 7013 2263 7014
rect 2310 7013 2311 7014
rect 2214 7015 2215 7016
rect 2262 7015 2263 7016
rect 1515 7017 1516 7018
rect 2214 7017 2215 7018
rect 2316 7017 2317 7018
rect 3334 7017 3335 7018
rect 2274 7019 2275 7020
rect 2316 7019 2317 7020
rect 2274 7021 2275 7022
rect 2298 7021 2299 7022
rect 2244 7023 2245 7024
rect 2298 7023 2299 7024
rect 2232 7025 2233 7026
rect 2244 7025 2245 7026
rect 2220 7027 2221 7028
rect 2232 7027 2233 7028
rect 2142 7029 2143 7030
rect 2220 7029 2221 7030
rect 2052 7031 2053 7032
rect 2142 7031 2143 7032
rect 1968 7033 1969 7034
rect 2052 7033 2053 7034
rect 1896 7035 1897 7036
rect 1968 7035 1969 7036
rect 1842 7037 1843 7038
rect 1896 7037 1897 7038
rect 1842 7039 1843 7040
rect 2304 7039 2305 7040
rect 2268 7041 2269 7042
rect 2304 7041 2305 7042
rect 2268 7043 2269 7044
rect 2868 7043 2869 7044
rect 2337 7045 2338 7046
rect 2769 7045 2770 7046
rect 2358 7047 2359 7048
rect 3199 7047 3200 7048
rect 2340 7049 2341 7050
rect 2358 7049 2359 7050
rect 1827 7051 1828 7052
rect 2340 7051 2341 7052
rect 2391 7051 2392 7052
rect 2427 7051 2428 7052
rect 2406 7053 2407 7054
rect 2442 7053 2443 7054
rect 2376 7055 2377 7056
rect 2406 7055 2407 7056
rect 2352 7057 2353 7058
rect 2376 7057 2377 7058
rect 2328 7059 2329 7060
rect 2352 7059 2353 7060
rect 2292 7061 2293 7062
rect 2328 7061 2329 7062
rect 2256 7063 2257 7064
rect 2292 7063 2293 7064
rect 2238 7065 2239 7066
rect 2256 7065 2257 7066
rect 2208 7067 2209 7068
rect 2238 7067 2239 7068
rect 2118 7069 2119 7070
rect 2208 7069 2209 7070
rect 2118 7071 2119 7072
rect 2202 7071 2203 7072
rect 2124 7073 2125 7074
rect 2202 7073 2203 7074
rect 2028 7075 2029 7076
rect 2124 7075 2125 7076
rect 2028 7077 2029 7078
rect 2082 7077 2083 7078
rect 1998 7079 1999 7080
rect 2082 7079 2083 7080
rect 1926 7081 1927 7082
rect 1998 7081 1999 7082
rect 1926 7083 1927 7084
rect 3300 7083 3301 7084
rect 2448 7085 2449 7086
rect 3276 7085 3277 7086
rect 2418 7087 2419 7088
rect 2448 7087 2449 7088
rect 2394 7089 2395 7090
rect 2418 7089 2419 7090
rect 2364 7091 2365 7092
rect 2394 7091 2395 7092
rect 2364 7093 2365 7094
rect 2370 7093 2371 7094
rect 2346 7095 2347 7096
rect 2370 7095 2371 7096
rect 2334 7097 2335 7098
rect 2346 7097 2347 7098
rect 1824 7099 1825 7100
rect 2334 7099 2335 7100
rect 1824 7101 1825 7102
rect 1830 7101 1831 7102
rect 1521 7103 1522 7104
rect 1830 7103 1831 7104
rect 2472 7103 2473 7104
rect 2490 7103 2491 7104
rect 2454 7105 2455 7106
rect 2472 7105 2473 7106
rect 2436 7107 2437 7108
rect 2454 7107 2455 7108
rect 2412 7109 2413 7110
rect 2436 7109 2437 7110
rect 2382 7111 2383 7112
rect 2412 7111 2413 7112
rect 2382 7113 2383 7114
rect 3303 7113 3304 7114
rect 2478 7115 2479 7116
rect 3159 7115 3160 7116
rect 2478 7117 2479 7118
rect 2520 7117 2521 7118
rect 2484 7119 2485 7120
rect 3273 7119 3274 7120
rect 2496 7121 2497 7122
rect 2538 7121 2539 7122
rect 2502 7123 2503 7124
rect 2520 7123 2521 7124
rect 1584 7125 1585 7126
rect 2502 7125 2503 7126
rect 1572 7127 1573 7128
rect 1584 7127 1585 7128
rect 1560 7129 1561 7130
rect 1572 7129 1573 7130
rect 2526 7129 2527 7130
rect 2538 7129 2539 7130
rect 2526 7131 2527 7132
rect 2562 7131 2563 7132
rect 2466 7133 2467 7134
rect 2562 7133 2563 7134
rect 1746 7135 1747 7136
rect 2466 7135 2467 7136
rect 2568 7135 2569 7136
rect 3163 7135 3164 7136
rect 2568 7137 2569 7138
rect 3288 7137 3289 7138
rect 2574 7139 2575 7140
rect 3285 7139 3286 7140
rect 2556 7141 2557 7142
rect 2574 7141 2575 7142
rect 1587 7143 1588 7144
rect 2556 7143 2557 7144
rect 2616 7143 2617 7144
rect 3302 7143 3303 7144
rect 2616 7145 2617 7146
rect 2628 7145 2629 7146
rect 2628 7147 2629 7148
rect 2646 7147 2647 7148
rect 2646 7149 2647 7150
rect 2664 7149 2665 7150
rect 2664 7151 2665 7152
rect 2682 7151 2683 7152
rect 2676 7153 2677 7154
rect 3268 7153 3269 7154
rect 2676 7155 2677 7156
rect 3317 7155 3318 7156
rect 2694 7157 2695 7158
rect 3264 7157 3265 7158
rect 2712 7159 2713 7160
rect 2790 7159 2791 7160
rect 2712 7161 2713 7162
rect 2724 7161 2725 7162
rect 2706 7163 2707 7164
rect 2724 7163 2725 7164
rect 2706 7165 2707 7166
rect 3320 7165 3321 7166
rect 2760 7167 2761 7168
rect 3117 7167 3118 7168
rect 2838 7169 2839 7170
rect 2868 7169 2869 7170
rect 1447 7171 1448 7172
rect 2838 7171 2839 7172
rect 2859 7171 2860 7172
rect 2889 7171 2890 7172
rect 2862 7173 2863 7174
rect 3296 7173 3297 7174
rect 2832 7175 2833 7176
rect 2862 7175 2863 7176
rect 2778 7177 2779 7178
rect 2832 7177 2833 7178
rect 2772 7179 2773 7180
rect 2778 7179 2779 7180
rect 2766 7181 2767 7182
rect 2772 7181 2773 7182
rect 1860 7183 1861 7184
rect 2766 7183 2767 7184
rect 1818 7185 1819 7186
rect 1860 7185 1861 7186
rect 1518 7187 1519 7188
rect 1818 7187 1819 7188
rect 2877 7187 2878 7188
rect 2907 7187 2908 7188
rect 2886 7189 2887 7190
rect 3224 7189 3225 7190
rect 2856 7191 2857 7192
rect 2886 7191 2887 7192
rect 2826 7193 2827 7194
rect 2856 7193 2857 7194
rect 2718 7195 2719 7196
rect 2826 7195 2827 7196
rect 2544 7197 2545 7198
rect 2718 7197 2719 7198
rect 2532 7199 2533 7200
rect 2544 7199 2545 7200
rect 2508 7201 2509 7202
rect 2532 7201 2533 7202
rect 2508 7203 2509 7204
rect 2550 7203 2551 7204
rect 1444 7205 1445 7206
rect 2550 7205 2551 7206
rect 2895 7205 2896 7206
rect 2913 7205 2914 7206
rect 2904 7207 2905 7208
rect 2934 7207 2935 7208
rect 2874 7209 2875 7210
rect 2904 7209 2905 7210
rect 2844 7211 2845 7212
rect 2874 7211 2875 7212
rect 2784 7213 2785 7214
rect 2844 7213 2845 7214
rect 2580 7215 2581 7216
rect 2784 7215 2785 7216
rect 2580 7217 2581 7218
rect 2592 7217 2593 7218
rect 2592 7219 2593 7220
rect 2598 7219 2599 7220
rect 2598 7221 2599 7222
rect 2610 7221 2611 7222
rect 2610 7223 2611 7224
rect 2622 7223 2623 7224
rect 2622 7225 2623 7226
rect 2640 7225 2641 7226
rect 2640 7227 2641 7228
rect 2652 7227 2653 7228
rect 2652 7229 2653 7230
rect 2670 7229 2671 7230
rect 2670 7231 2671 7232
rect 2700 7231 2701 7232
rect 2700 7233 2701 7234
rect 2730 7233 2731 7234
rect 2730 7235 2731 7236
rect 2736 7235 2737 7236
rect 2736 7237 2737 7238
rect 2742 7237 2743 7238
rect 1539 7239 1540 7240
rect 2742 7239 2743 7240
rect 2940 7239 2941 7240
rect 3295 7239 3296 7240
rect 2898 7241 2899 7242
rect 2940 7241 2941 7242
rect 2892 7243 2893 7244
rect 2898 7243 2899 7244
rect 2892 7245 2893 7246
rect 2910 7245 2911 7246
rect 2880 7247 2881 7248
rect 2910 7247 2911 7248
rect 2850 7249 2851 7250
rect 2880 7249 2881 7250
rect 2820 7251 2821 7252
rect 2850 7251 2851 7252
rect 2802 7253 2803 7254
rect 2820 7253 2821 7254
rect 2796 7255 2797 7256
rect 2802 7255 2803 7256
rect 2796 7257 2797 7258
rect 3261 7257 3262 7258
rect 2964 7259 2965 7260
rect 2991 7259 2992 7260
rect 2946 7261 2947 7262
rect 2964 7261 2965 7262
rect 2916 7263 2917 7264
rect 2946 7263 2947 7264
rect 2916 7265 2917 7266
rect 3262 7265 3263 7266
rect 3006 7267 3007 7268
rect 3042 7267 3043 7268
rect 3006 7269 3007 7270
rect 3012 7269 3013 7270
rect 2982 7271 2983 7272
rect 3012 7271 3013 7272
rect 3009 7273 3010 7274
rect 3015 7273 3016 7274
rect 3030 7273 3031 7274
rect 3072 7273 3073 7274
rect 3030 7275 3031 7276
rect 3299 7275 3300 7276
rect 3036 7277 3037 7278
rect 3141 7277 3142 7278
rect 3000 7279 3001 7280
rect 3036 7279 3037 7280
rect 2958 7281 2959 7282
rect 3000 7281 3001 7282
rect 3048 7281 3049 7282
rect 3084 7281 3085 7282
rect 2976 7283 2977 7284
rect 3048 7283 3049 7284
rect 2922 7285 2923 7286
rect 2976 7285 2977 7286
rect 3066 7285 3067 7286
rect 3096 7285 3097 7286
rect 3024 7287 3025 7288
rect 3066 7287 3067 7288
rect 2994 7289 2995 7290
rect 3024 7289 3025 7290
rect 2994 7291 2995 7292
rect 3081 7291 3082 7292
rect 3078 7293 3079 7294
rect 3156 7293 3157 7294
rect 3105 7295 3106 7296
rect 3135 7295 3136 7296
rect 3108 7297 3109 7298
rect 3138 7297 3139 7298
rect 3111 7299 3112 7300
rect 3239 7299 3240 7300
rect 3123 7301 3124 7302
rect 3153 7301 3154 7302
rect 3132 7303 3133 7304
rect 3162 7303 3163 7304
rect 3102 7305 3103 7306
rect 3132 7305 3133 7306
rect 3102 7307 3103 7308
rect 3233 7307 3234 7308
rect 3144 7309 3145 7310
rect 3174 7309 3175 7310
rect 3147 7311 3148 7312
rect 3177 7311 3178 7312
rect 3159 7313 3160 7314
rect 3227 7313 3228 7314
rect 3166 7315 3167 7316
rect 3311 7315 3312 7316
rect 3169 7317 3170 7318
rect 3199 7317 3200 7318
rect 3181 7319 3182 7320
rect 3223 7319 3224 7320
rect 3150 7321 3151 7322
rect 3180 7321 3181 7322
rect 3120 7323 3121 7324
rect 3150 7323 3151 7324
rect 3090 7325 3091 7326
rect 3120 7325 3121 7326
rect 3060 7327 3061 7328
rect 3090 7327 3091 7328
rect 3054 7329 3055 7330
rect 3060 7329 3061 7330
rect 3018 7331 3019 7332
rect 3054 7331 3055 7332
rect 2988 7333 2989 7334
rect 3018 7333 3019 7334
rect 2970 7335 2971 7336
rect 2988 7335 2989 7336
rect 2952 7337 2953 7338
rect 2970 7337 2971 7338
rect 2928 7339 2929 7340
rect 2952 7339 2953 7340
rect 3193 7339 3194 7340
rect 3235 7339 3236 7340
rect 2922 7341 2923 7342
rect 3193 7341 3194 7342
rect 3196 7341 3197 7342
rect 3238 7341 3239 7342
rect 2928 7343 2929 7344
rect 3196 7343 3197 7344
rect 3205 7343 3206 7344
rect 3243 7343 3244 7344
rect 3114 7345 3115 7346
rect 3244 7345 3245 7346
rect 3211 7347 3212 7348
rect 3253 7347 3254 7348
rect 3217 7349 3218 7350
rect 3241 7349 3242 7350
rect 3220 7351 3221 7352
rect 3269 7351 3270 7352
rect 3255 7353 3256 7354
rect 3324 7353 3325 7354
rect 3214 7355 3215 7356
rect 3256 7355 3257 7356
rect 3258 7355 3259 7356
rect 3271 7355 3272 7356
rect 3126 7357 3127 7358
rect 3259 7357 3260 7358
rect 3280 7357 3281 7358
rect 3293 7357 3294 7358
rect 2958 7359 2959 7360
rect 3292 7359 3293 7360
rect 3230 7361 3231 7362
rect 3279 7361 3280 7362
rect 3187 7363 3188 7364
rect 3229 7363 3230 7364
rect 2088 7365 2089 7366
rect 3186 7365 3187 7366
rect 3283 7365 3284 7366
rect 3314 7365 3315 7366
rect 3246 7367 3247 7368
rect 3282 7367 3283 7368
rect 1423 7376 1424 7377
rect 1728 7376 1729 7377
rect 1423 7378 1424 7379
rect 1848 7378 1849 7379
rect 1430 7380 1431 7381
rect 1776 7380 1777 7381
rect 1433 7382 1434 7383
rect 1644 7382 1645 7383
rect 1437 7384 1438 7385
rect 1463 7384 1464 7385
rect 1438 7386 1439 7387
rect 1986 7386 1987 7387
rect 1444 7388 1445 7389
rect 1469 7388 1470 7389
rect 1445 7390 1446 7391
rect 1572 7390 1573 7391
rect 1447 7392 1448 7393
rect 2760 7392 2761 7393
rect 1449 7394 1450 7395
rect 1536 7394 1537 7395
rect 1451 7396 1452 7397
rect 2106 7396 2107 7397
rect 1452 7398 1453 7399
rect 1530 7398 1531 7399
rect 1454 7400 1455 7401
rect 1794 7400 1795 7401
rect 1461 7402 1462 7403
rect 1728 7402 1729 7403
rect 1464 7404 1465 7405
rect 1806 7404 1807 7405
rect 1468 7406 1469 7407
rect 1752 7406 1753 7407
rect 1475 7408 1476 7409
rect 1571 7408 1572 7409
rect 1478 7410 1479 7411
rect 2190 7410 2191 7411
rect 1480 7412 1481 7413
rect 1500 7412 1501 7413
rect 1482 7414 1483 7415
rect 1980 7414 1981 7415
rect 1485 7416 1486 7417
rect 2895 7416 2896 7417
rect 1492 7418 1493 7419
rect 3081 7418 3082 7419
rect 1504 7420 1505 7421
rect 1512 7420 1513 7421
rect 1510 7422 1511 7423
rect 1554 7422 1555 7423
rect 1442 7424 1443 7425
rect 1553 7424 1554 7425
rect 1513 7426 1514 7427
rect 2214 7426 2215 7427
rect 1518 7428 1519 7429
rect 2994 7428 2995 7429
rect 1517 7430 1518 7431
rect 1638 7430 1639 7431
rect 1521 7432 1522 7433
rect 1524 7432 1525 7433
rect 1523 7434 1524 7435
rect 1620 7434 1621 7435
rect 1551 7436 1552 7437
rect 2532 7436 2533 7437
rect 1559 7438 1560 7439
rect 1578 7438 1579 7439
rect 1580 7438 1581 7439
rect 2880 7438 2881 7439
rect 1589 7440 1590 7441
rect 1608 7440 1609 7441
rect 1599 7442 1600 7443
rect 2160 7442 2161 7443
rect 1602 7444 1603 7445
rect 2298 7444 2299 7445
rect 1605 7446 1606 7447
rect 2256 7446 2257 7447
rect 1614 7448 1615 7449
rect 1626 7448 1627 7449
rect 1623 7450 1624 7451
rect 2478 7450 2479 7451
rect 1626 7452 1627 7453
rect 1662 7452 1663 7453
rect 1644 7454 1645 7455
rect 3000 7454 3001 7455
rect 1656 7456 1657 7457
rect 2268 7456 2269 7457
rect 1662 7458 1663 7459
rect 2562 7458 2563 7459
rect 1520 7460 1521 7461
rect 2562 7460 2563 7461
rect 1668 7462 1669 7463
rect 1716 7462 1717 7463
rect 1692 7464 1693 7465
rect 1752 7464 1753 7465
rect 1710 7466 1711 7467
rect 2367 7466 2368 7467
rect 1686 7468 1687 7469
rect 1710 7468 1711 7469
rect 1650 7470 1651 7471
rect 1686 7470 1687 7471
rect 1650 7472 1651 7473
rect 3006 7472 3007 7473
rect 1716 7474 1717 7475
rect 3090 7474 3091 7475
rect 1746 7476 1747 7477
rect 2634 7476 2635 7477
rect 1746 7478 1747 7479
rect 2916 7478 2917 7479
rect 1749 7480 1750 7481
rect 2910 7480 2911 7481
rect 1776 7482 1777 7483
rect 2784 7482 2785 7483
rect 1782 7484 1783 7485
rect 1848 7484 1849 7485
rect 1782 7486 1783 7487
rect 2868 7486 2869 7487
rect 1794 7488 1795 7489
rect 2862 7488 2863 7489
rect 1806 7490 1807 7491
rect 2718 7490 2719 7491
rect 1824 7492 1825 7493
rect 1986 7492 1987 7493
rect 1722 7494 1723 7495
rect 1824 7494 1825 7495
rect 1722 7496 1723 7497
rect 2940 7496 2941 7497
rect 1896 7498 1897 7499
rect 2106 7498 2107 7499
rect 1788 7500 1789 7501
rect 1896 7500 1897 7501
rect 1471 7502 1472 7503
rect 1788 7502 1789 7503
rect 1905 7502 1906 7503
rect 2115 7502 2116 7503
rect 1959 7504 1960 7505
rect 2283 7504 2284 7505
rect 1974 7506 1975 7507
rect 2160 7506 2161 7507
rect 1974 7508 1975 7509
rect 2832 7508 2833 7509
rect 1980 7510 1981 7511
rect 2850 7510 2851 7511
rect 2001 7512 2002 7513
rect 2277 7512 2278 7513
rect 2016 7514 2017 7515
rect 2298 7514 2299 7515
rect 2016 7516 2017 7517
rect 2466 7516 2467 7517
rect 2025 7518 2026 7519
rect 2313 7518 2314 7519
rect 2028 7520 2029 7521
rect 2256 7520 2257 7521
rect 2028 7522 2029 7523
rect 2736 7522 2737 7523
rect 2043 7524 2044 7525
rect 2289 7524 2290 7525
rect 2100 7526 2101 7527
rect 3184 7526 3185 7527
rect 2100 7528 2101 7529
rect 2388 7528 2389 7529
rect 2088 7530 2089 7531
rect 2388 7530 2389 7531
rect 1890 7532 1891 7533
rect 2088 7532 2089 7533
rect 1764 7534 1765 7535
rect 1890 7534 1891 7535
rect 2190 7534 2191 7535
rect 2358 7534 2359 7535
rect 2064 7536 2065 7537
rect 2358 7536 2359 7537
rect 2064 7538 2065 7539
rect 2640 7538 2641 7539
rect 2193 7540 2194 7541
rect 2295 7540 2296 7541
rect 2208 7542 2209 7543
rect 2478 7542 2479 7543
rect 1950 7544 1951 7545
rect 2208 7544 2209 7545
rect 1812 7546 1813 7547
rect 1950 7546 1951 7547
rect 1812 7548 1813 7549
rect 1878 7548 1879 7549
rect 1818 7550 1819 7551
rect 1878 7550 1879 7551
rect 1548 7552 1549 7553
rect 1818 7552 1819 7553
rect 1547 7554 1548 7555
rect 1566 7554 1567 7555
rect 1565 7556 1566 7557
rect 1584 7556 1585 7557
rect 2214 7556 2215 7557
rect 2550 7556 2551 7557
rect 2235 7558 2236 7559
rect 2355 7558 2356 7559
rect 1971 7560 1972 7561
rect 2235 7560 2236 7561
rect 2238 7560 2239 7561
rect 2466 7560 2467 7561
rect 1992 7562 1993 7563
rect 2238 7562 2239 7563
rect 1836 7564 1837 7565
rect 1992 7564 1993 7565
rect 1598 7566 1599 7567
rect 1836 7566 1837 7567
rect 2244 7566 2245 7567
rect 3186 7566 3187 7567
rect 1440 7568 1441 7569
rect 2244 7568 2245 7569
rect 2268 7568 2269 7569
rect 2274 7568 2275 7569
rect 1998 7570 1999 7571
rect 2274 7570 2275 7571
rect 1842 7572 1843 7573
rect 1998 7572 1999 7573
rect 1758 7574 1759 7575
rect 1842 7574 1843 7575
rect 1698 7576 1699 7577
rect 1758 7576 1759 7577
rect 1698 7578 1699 7579
rect 1704 7578 1705 7579
rect 2286 7578 2287 7579
rect 2532 7578 2533 7579
rect 2004 7580 2005 7581
rect 2286 7580 2287 7581
rect 2004 7582 2005 7583
rect 2724 7582 2725 7583
rect 2316 7584 2317 7585
rect 3189 7584 3190 7585
rect 2316 7586 2317 7587
rect 2352 7586 2353 7587
rect 2052 7588 2053 7589
rect 2352 7588 2353 7589
rect 1854 7590 1855 7591
rect 2052 7590 2053 7591
rect 1426 7592 1427 7593
rect 1854 7592 1855 7593
rect 1426 7594 1427 7595
rect 1866 7594 1867 7595
rect 1740 7596 1741 7597
rect 1866 7596 1867 7597
rect 1680 7598 1681 7599
rect 1740 7598 1741 7599
rect 1680 7600 1681 7601
rect 2892 7600 2893 7601
rect 2337 7602 2338 7603
rect 2391 7602 2392 7603
rect 2361 7604 2362 7605
rect 2769 7604 2770 7605
rect 2406 7606 2407 7607
rect 3276 7606 3277 7607
rect 2166 7608 2167 7609
rect 2406 7608 2407 7609
rect 2166 7610 2167 7611
rect 2280 7610 2281 7611
rect 2280 7612 2281 7613
rect 3187 7612 3188 7613
rect 2412 7614 2413 7615
rect 3212 7614 3213 7615
rect 2124 7616 2125 7617
rect 2412 7616 2413 7617
rect 1926 7618 1927 7619
rect 2124 7618 2125 7619
rect 1926 7620 1927 7621
rect 2556 7620 2557 7621
rect 2394 7622 2395 7623
rect 2556 7622 2557 7623
rect 2130 7624 2131 7625
rect 2394 7624 2395 7625
rect 2076 7626 2077 7627
rect 2130 7626 2131 7627
rect 1914 7628 1915 7629
rect 2076 7628 2077 7629
rect 1914 7630 1915 7631
rect 2742 7630 2743 7631
rect 2454 7632 2455 7633
rect 2550 7632 2551 7633
rect 2322 7634 2323 7635
rect 2454 7634 2455 7635
rect 2034 7636 2035 7637
rect 2322 7636 2323 7637
rect 2034 7638 2035 7639
rect 3170 7638 3171 7639
rect 2460 7640 2461 7641
rect 3266 7640 3267 7641
rect 2172 7642 2173 7643
rect 2460 7642 2461 7643
rect 1938 7644 1939 7645
rect 2172 7644 2173 7645
rect 1938 7646 1939 7647
rect 2790 7646 2791 7647
rect 2472 7648 2473 7649
rect 3262 7648 3263 7649
rect 2202 7650 2203 7651
rect 2472 7650 2473 7651
rect 1956 7652 1957 7653
rect 2202 7652 2203 7653
rect 1920 7654 1921 7655
rect 1956 7654 1957 7655
rect 1920 7656 1921 7657
rect 2502 7656 2503 7657
rect 2340 7658 2341 7659
rect 2502 7658 2503 7659
rect 2046 7660 2047 7661
rect 2340 7660 2341 7661
rect 1435 7662 1436 7663
rect 2046 7662 2047 7663
rect 2490 7662 2491 7663
rect 2640 7662 2641 7663
rect 2262 7664 2263 7665
rect 2490 7664 2491 7665
rect 2040 7666 2041 7667
rect 2262 7666 2263 7667
rect 2040 7668 2041 7669
rect 2526 7668 2527 7669
rect 2508 7670 2509 7671
rect 3166 7670 3167 7671
rect 2304 7672 2305 7673
rect 2508 7672 2509 7673
rect 2094 7674 2095 7675
rect 2304 7674 2305 7675
rect 1908 7676 1909 7677
rect 2094 7676 2095 7677
rect 1770 7678 1771 7679
rect 1908 7678 1909 7679
rect 1770 7680 1771 7681
rect 2874 7680 2875 7681
rect 2514 7682 2515 7683
rect 3144 7682 3145 7683
rect 2514 7684 2515 7685
rect 2544 7684 2545 7685
rect 2310 7686 2311 7687
rect 2544 7686 2545 7687
rect 2022 7688 2023 7689
rect 2310 7688 2311 7689
rect 2022 7690 2023 7691
rect 2496 7690 2497 7691
rect 2250 7692 2251 7693
rect 2496 7692 2497 7693
rect 2010 7694 2011 7695
rect 2250 7694 2251 7695
rect 2010 7696 2011 7697
rect 2838 7696 2839 7697
rect 2526 7698 2527 7699
rect 3269 7698 3270 7699
rect 2538 7700 2539 7701
rect 2634 7700 2635 7701
rect 2292 7702 2293 7703
rect 2538 7702 2539 7703
rect 2184 7704 2185 7705
rect 2292 7704 2293 7705
rect 2184 7706 2185 7707
rect 2232 7706 2233 7707
rect 1968 7708 1969 7709
rect 2232 7708 2233 7709
rect 1968 7710 1969 7711
rect 3273 7710 3274 7711
rect 2610 7712 2611 7713
rect 3299 7712 3300 7713
rect 2424 7714 2425 7715
rect 2610 7714 2611 7715
rect 2136 7716 2137 7717
rect 2424 7716 2425 7717
rect 2118 7718 2119 7719
rect 2136 7718 2137 7719
rect 2118 7720 2119 7721
rect 2364 7720 2365 7721
rect 1596 7722 1597 7723
rect 2364 7722 2365 7723
rect 1595 7724 1596 7725
rect 2832 7724 2833 7725
rect 2616 7726 2617 7727
rect 3302 7726 3303 7727
rect 2436 7728 2437 7729
rect 2616 7728 2617 7729
rect 2196 7730 2197 7731
rect 2436 7730 2437 7731
rect 2196 7732 2197 7733
rect 2580 7732 2581 7733
rect 2370 7734 2371 7735
rect 2580 7734 2581 7735
rect 2646 7734 2647 7735
rect 2724 7734 2725 7735
rect 2664 7736 2665 7737
rect 2736 7736 2737 7737
rect 2568 7738 2569 7739
rect 2664 7738 2665 7739
rect 2568 7740 2569 7741
rect 3327 7740 3328 7741
rect 2670 7742 2671 7743
rect 2742 7742 2743 7743
rect 2670 7744 2671 7745
rect 3288 7744 3289 7745
rect 2682 7746 2683 7747
rect 3324 7746 3325 7747
rect 2688 7748 2689 7749
rect 3320 7748 3321 7749
rect 2574 7750 2575 7751
rect 2688 7750 2689 7751
rect 2520 7752 2521 7753
rect 2574 7752 2575 7753
rect 2484 7754 2485 7755
rect 2520 7754 2521 7755
rect 2220 7756 2221 7757
rect 2484 7756 2485 7757
rect 2148 7758 2149 7759
rect 2220 7758 2221 7759
rect 1932 7760 1933 7761
rect 2148 7760 2149 7761
rect 1932 7762 1933 7763
rect 2400 7762 2401 7763
rect 2142 7764 2143 7765
rect 2400 7764 2401 7765
rect 2142 7766 2143 7767
rect 3334 7766 3335 7767
rect 2694 7768 2695 7769
rect 3147 7768 3148 7769
rect 2604 7770 2605 7771
rect 2694 7770 2695 7771
rect 2604 7772 2605 7773
rect 3209 7772 3210 7773
rect 2700 7774 2701 7775
rect 2718 7774 2719 7775
rect 2622 7776 2623 7777
rect 2700 7776 2701 7777
rect 2442 7778 2443 7779
rect 2622 7778 2623 7779
rect 2334 7780 2335 7781
rect 2442 7780 2443 7781
rect 2058 7782 2059 7783
rect 2334 7782 2335 7783
rect 1860 7784 1861 7785
rect 2058 7784 2059 7785
rect 1734 7786 1735 7787
rect 1860 7786 1861 7787
rect 1674 7788 1675 7789
rect 1734 7788 1735 7789
rect 1577 7790 1578 7791
rect 1674 7790 1675 7791
rect 2706 7790 2707 7791
rect 2760 7790 2761 7791
rect 2628 7792 2629 7793
rect 2706 7792 2707 7793
rect 2448 7794 2449 7795
rect 2628 7794 2629 7795
rect 2178 7796 2179 7797
rect 2448 7796 2449 7797
rect 2178 7798 2179 7799
rect 2346 7798 2347 7799
rect 2070 7800 2071 7801
rect 2346 7800 2347 7801
rect 1884 7802 1885 7803
rect 2070 7802 2071 7803
rect 1800 7804 1801 7805
rect 1884 7804 1885 7805
rect 1800 7806 1801 7807
rect 2856 7806 2857 7807
rect 2754 7808 2755 7809
rect 3015 7808 3016 7809
rect 2784 7810 2785 7811
rect 2844 7810 2845 7811
rect 2790 7812 2791 7813
rect 2796 7812 2797 7813
rect 2772 7814 2773 7815
rect 2796 7814 2797 7815
rect 2748 7816 2749 7817
rect 2772 7816 2773 7817
rect 2676 7818 2677 7819
rect 2748 7818 2749 7819
rect 2586 7820 2587 7821
rect 2676 7820 2677 7821
rect 2376 7822 2377 7823
rect 2586 7822 2587 7823
rect 2112 7824 2113 7825
rect 2376 7824 2377 7825
rect 1902 7826 1903 7827
rect 2112 7826 2113 7827
rect 1830 7828 1831 7829
rect 1902 7828 1903 7829
rect 1830 7830 1831 7831
rect 1872 7830 1873 7831
rect 1872 7832 1873 7833
rect 2766 7832 2767 7833
rect 2712 7834 2713 7835
rect 2766 7834 2767 7835
rect 2658 7836 2659 7837
rect 2712 7836 2713 7837
rect 2592 7838 2593 7839
rect 2658 7838 2659 7839
rect 2418 7840 2419 7841
rect 2592 7840 2593 7841
rect 2328 7842 2329 7843
rect 2418 7842 2419 7843
rect 2226 7844 2227 7845
rect 2328 7844 2329 7845
rect 1962 7846 1963 7847
rect 2226 7846 2227 7847
rect 1962 7848 1963 7849
rect 3331 7848 3332 7849
rect 2814 7850 2815 7851
rect 2820 7850 2821 7851
rect 2835 7850 2836 7851
rect 3009 7850 3010 7851
rect 2838 7852 2839 7853
rect 2946 7852 2947 7853
rect 2844 7854 2845 7855
rect 2976 7854 2977 7855
rect 2850 7856 2851 7857
rect 2898 7856 2899 7857
rect 2856 7858 2857 7859
rect 2922 7858 2923 7859
rect 2862 7860 2863 7861
rect 2886 7860 2887 7861
rect 2865 7862 2866 7863
rect 2889 7862 2890 7863
rect 2868 7864 2869 7865
rect 2928 7864 2929 7865
rect 2874 7866 2875 7867
rect 3096 7866 3097 7867
rect 2880 7868 2881 7869
rect 2904 7868 2905 7869
rect 2883 7870 2884 7871
rect 2907 7870 2908 7871
rect 2886 7872 2887 7873
rect 3129 7872 3130 7873
rect 2892 7874 2893 7875
rect 3156 7874 3157 7875
rect 2895 7876 2896 7877
rect 3159 7876 3160 7877
rect 2898 7878 2899 7879
rect 3012 7878 3013 7879
rect 2904 7880 2905 7881
rect 2958 7880 2959 7881
rect 2910 7882 2911 7883
rect 2952 7882 2953 7883
rect 2916 7884 2917 7885
rect 3295 7884 3296 7885
rect 2922 7886 2923 7887
rect 2970 7886 2971 7887
rect 2928 7888 2929 7889
rect 3018 7888 3019 7889
rect 2934 7890 2935 7891
rect 3196 7890 3197 7891
rect 2940 7892 2941 7893
rect 2988 7892 2989 7893
rect 2943 7894 2944 7895
rect 2991 7894 2992 7895
rect 2946 7896 2947 7897
rect 3030 7896 3031 7897
rect 2952 7898 2953 7899
rect 3259 7898 3260 7899
rect 2958 7900 2959 7901
rect 3024 7900 3025 7901
rect 2964 7902 2965 7903
rect 3292 7902 3293 7903
rect 2964 7904 2965 7905
rect 3317 7904 3318 7905
rect 2970 7906 2971 7907
rect 3036 7906 3037 7907
rect 2976 7908 2977 7909
rect 3042 7908 3043 7909
rect 2982 7910 2983 7911
rect 3066 7910 3067 7911
rect 2370 7912 2371 7913
rect 3066 7912 3067 7913
rect 2988 7914 2989 7915
rect 3072 7914 3073 7915
rect 2994 7916 2995 7917
rect 3141 7916 3142 7917
rect 3000 7918 3001 7919
rect 3084 7918 3085 7919
rect 3006 7920 3007 7921
rect 3150 7920 3151 7921
rect 3009 7922 3010 7923
rect 3054 7922 3055 7923
rect 3012 7924 3013 7925
rect 3244 7924 3245 7925
rect 3018 7926 3019 7927
rect 3102 7926 3103 7927
rect 3030 7928 3031 7929
rect 3138 7928 3139 7929
rect 3033 7930 3034 7931
rect 3069 7930 3070 7931
rect 3036 7932 3037 7933
rect 3120 7932 3121 7933
rect 3048 7934 3049 7935
rect 3126 7934 3127 7935
rect 3048 7936 3049 7937
rect 3132 7936 3133 7937
rect 3051 7938 3052 7939
rect 3135 7938 3136 7939
rect 3054 7940 3055 7941
rect 3162 7940 3163 7941
rect 3060 7942 3061 7943
rect 3163 7942 3164 7943
rect 3060 7944 3061 7945
rect 3177 7944 3178 7945
rect 3063 7946 3064 7947
rect 3174 7946 3175 7947
rect 2730 7948 2731 7949
rect 3173 7948 3174 7949
rect 2652 7950 2653 7951
rect 2730 7950 2731 7951
rect 2652 7952 2653 7953
rect 3202 7952 3203 7953
rect 3072 7954 3073 7955
rect 3180 7954 3181 7955
rect 2646 7956 2647 7957
rect 3180 7956 3181 7957
rect 3078 7958 3079 7959
rect 3153 7958 3154 7959
rect 3084 7960 3085 7961
rect 3199 7960 3200 7961
rect 3096 7962 3097 7963
rect 3205 7962 3206 7963
rect 2382 7964 2383 7965
rect 3205 7964 3206 7965
rect 2082 7966 2083 7967
rect 2382 7966 2383 7967
rect 2082 7968 2083 7969
rect 2598 7968 2599 7969
rect 2430 7970 2431 7971
rect 2598 7970 2599 7971
rect 2154 7972 2155 7973
rect 2430 7972 2431 7973
rect 1944 7974 1945 7975
rect 2154 7974 2155 7975
rect 1944 7976 1945 7977
rect 2826 7976 2827 7977
rect 2808 7978 2809 7979
rect 2826 7978 2827 7979
rect 2802 7980 2803 7981
rect 2808 7980 2809 7981
rect 2778 7982 2779 7983
rect 2802 7982 2803 7983
rect 3108 7982 3109 7983
rect 3223 7982 3224 7983
rect 3114 7984 3115 7985
rect 3229 7984 3230 7985
rect 3120 7986 3121 7987
rect 3235 7986 3236 7987
rect 3123 7988 3124 7989
rect 3238 7988 3239 7989
rect 3138 7990 3139 7991
rect 3253 7990 3254 7991
rect 3141 7992 3142 7993
rect 3151 7992 3152 7993
rect 3154 7992 3155 7993
rect 3256 7992 3257 7993
rect 3157 7994 3158 7995
rect 3279 7994 3280 7995
rect 3160 7996 3161 7997
rect 3282 7996 3283 7997
rect 3177 7998 3178 7999
rect 3241 7998 3242 7999
rect 3193 8000 3194 8001
rect 3285 8000 3286 8001
rect 3196 8002 3197 8003
rect 3311 8002 3312 8003
rect 3199 8004 3200 8005
rect 3314 8004 3315 8005
rect 1423 8013 1424 8014
rect 1440 8013 1441 8014
rect 1423 8015 1424 8016
rect 2208 8015 2209 8016
rect 1426 8017 1427 8018
rect 2046 8017 2047 8018
rect 1430 8019 1431 8020
rect 1488 8019 1489 8020
rect 1433 8021 1434 8022
rect 1492 8021 1493 8022
rect 1438 8023 1439 8024
rect 1926 8023 1927 8024
rect 1445 8025 1446 8026
rect 2289 8025 2290 8026
rect 1444 8027 1445 8028
rect 2322 8027 2323 8028
rect 1452 8029 1453 8030
rect 1523 8029 1524 8030
rect 1454 8031 1455 8032
rect 1890 8031 1891 8032
rect 1461 8033 1462 8034
rect 1830 8033 1831 8034
rect 1464 8035 1465 8036
rect 1812 8035 1813 8036
rect 1463 8037 1464 8038
rect 1896 8037 1897 8038
rect 1437 8039 1438 8040
rect 1896 8039 1897 8040
rect 1466 8041 1467 8042
rect 1812 8041 1813 8042
rect 1468 8043 1469 8044
rect 1547 8043 1548 8044
rect 1471 8045 1472 8046
rect 1575 8045 1576 8046
rect 1480 8047 1481 8048
rect 1494 8047 1495 8048
rect 1504 8047 1505 8048
rect 1506 8047 1507 8048
rect 1510 8047 1511 8048
rect 2370 8047 2371 8048
rect 1520 8049 1521 8050
rect 2358 8049 2359 8050
rect 1524 8051 1525 8052
rect 1764 8051 1765 8052
rect 1527 8053 1528 8054
rect 1914 8053 1915 8054
rect 1548 8055 1549 8056
rect 1553 8055 1554 8056
rect 1554 8057 1555 8058
rect 1559 8057 1560 8058
rect 1560 8059 1561 8060
rect 1565 8059 1566 8060
rect 1566 8061 1567 8062
rect 1571 8061 1572 8062
rect 1572 8063 1573 8064
rect 1650 8063 1651 8064
rect 1577 8065 1578 8066
rect 3051 8065 3052 8066
rect 1584 8067 1585 8068
rect 1589 8067 1590 8068
rect 1590 8069 1591 8070
rect 1626 8069 1627 8070
rect 1593 8071 1594 8072
rect 3054 8071 3055 8072
rect 1595 8073 1596 8074
rect 1800 8073 1801 8074
rect 1598 8075 1599 8076
rect 1794 8075 1795 8076
rect 1602 8077 1603 8078
rect 2454 8077 2455 8078
rect 1602 8079 1603 8080
rect 1614 8079 1615 8080
rect 1614 8081 1615 8082
rect 1674 8081 1675 8082
rect 1620 8083 1621 8084
rect 1686 8083 1687 8084
rect 1638 8085 1639 8086
rect 1698 8085 1699 8086
rect 1650 8087 1651 8088
rect 1734 8087 1735 8088
rect 1656 8089 1657 8090
rect 1692 8089 1693 8090
rect 1656 8091 1657 8092
rect 1740 8091 1741 8092
rect 1662 8093 1663 8094
rect 1698 8093 1699 8094
rect 1662 8095 1663 8096
rect 1668 8095 1669 8096
rect 1668 8097 1669 8098
rect 1752 8097 1753 8098
rect 1674 8099 1675 8100
rect 1758 8099 1759 8100
rect 1686 8101 1687 8102
rect 1728 8101 1729 8102
rect 1704 8103 1705 8104
rect 1788 8103 1789 8104
rect 1716 8105 1717 8106
rect 2778 8105 2779 8106
rect 1716 8107 1717 8108
rect 1776 8107 1777 8108
rect 1722 8109 1723 8110
rect 2745 8109 2746 8110
rect 1722 8111 1723 8112
rect 1806 8111 1807 8112
rect 1451 8113 1452 8114
rect 1806 8113 1807 8114
rect 1728 8115 1729 8116
rect 1818 8115 1819 8116
rect 1734 8117 1735 8118
rect 1824 8117 1825 8118
rect 1740 8119 1741 8120
rect 1782 8119 1783 8120
rect 1752 8121 1753 8122
rect 1842 8121 1843 8122
rect 1758 8123 1759 8124
rect 1848 8123 1849 8124
rect 1776 8125 1777 8126
rect 1854 8125 1855 8126
rect 1782 8127 1783 8128
rect 1860 8127 1861 8128
rect 1788 8129 1789 8130
rect 1866 8129 1867 8130
rect 1794 8131 1795 8132
rect 1902 8131 1903 8132
rect 1800 8133 1801 8134
rect 1884 8133 1885 8134
rect 1818 8135 1819 8136
rect 1878 8135 1879 8136
rect 1824 8137 1825 8138
rect 1920 8137 1921 8138
rect 1830 8139 1831 8140
rect 1944 8139 1945 8140
rect 1842 8141 1843 8142
rect 1908 8141 1909 8142
rect 1836 8143 1837 8144
rect 1908 8143 1909 8144
rect 1836 8145 1837 8146
rect 1932 8145 1933 8146
rect 1848 8147 1849 8148
rect 1974 8147 1975 8148
rect 1854 8149 1855 8150
rect 1980 8149 1981 8150
rect 1860 8151 1861 8152
rect 2010 8151 2011 8152
rect 1866 8153 1867 8154
rect 2784 8153 2785 8154
rect 1878 8155 1879 8156
rect 1962 8155 1963 8156
rect 1884 8157 1885 8158
rect 1968 8157 1969 8158
rect 1890 8159 1891 8160
rect 1950 8159 1951 8160
rect 1902 8161 1903 8162
rect 2004 8161 2005 8162
rect 1473 8163 1474 8164
rect 2004 8163 2005 8164
rect 1914 8165 1915 8166
rect 2772 8165 2773 8166
rect 1926 8167 1927 8168
rect 2034 8167 2035 8168
rect 1932 8169 1933 8170
rect 3184 8169 3185 8170
rect 1944 8171 1945 8172
rect 1992 8171 1993 8172
rect 1950 8173 1951 8174
rect 1998 8173 1999 8174
rect 1962 8175 1963 8176
rect 2016 8175 2017 8176
rect 1968 8177 1969 8178
rect 2022 8177 2023 8178
rect 1974 8179 1975 8180
rect 2760 8179 2761 8180
rect 1980 8181 1981 8182
rect 2040 8181 2041 8182
rect 1992 8183 1993 8184
rect 2052 8183 2053 8184
rect 1998 8185 1999 8186
rect 2058 8185 2059 8186
rect 2010 8187 2011 8188
rect 2082 8187 2083 8188
rect 2016 8189 2017 8190
rect 2070 8189 2071 8190
rect 2022 8191 2023 8192
rect 2076 8191 2077 8192
rect 2028 8193 2029 8194
rect 3170 8193 3171 8194
rect 2028 8195 2029 8196
rect 2682 8195 2683 8196
rect 2034 8197 2035 8198
rect 2100 8197 2101 8198
rect 2040 8199 2041 8200
rect 2088 8199 2089 8200
rect 2046 8201 2047 8202
rect 2106 8201 2107 8202
rect 2052 8203 2053 8204
rect 2112 8203 2113 8204
rect 2055 8205 2056 8206
rect 2115 8205 2116 8206
rect 2058 8207 2059 8208
rect 2094 8207 2095 8208
rect 2064 8209 2065 8210
rect 3041 8209 3042 8210
rect 2064 8211 2065 8212
rect 2118 8211 2119 8212
rect 1447 8213 1448 8214
rect 2118 8213 2119 8214
rect 2070 8215 2071 8216
rect 2142 8215 2143 8216
rect 2076 8217 2077 8218
rect 2124 8217 2125 8218
rect 2082 8219 2083 8220
rect 2130 8219 2131 8220
rect 2088 8221 2089 8222
rect 2136 8221 2137 8222
rect 2094 8223 2095 8224
rect 2154 8223 2155 8224
rect 2100 8225 2101 8226
rect 2148 8225 2149 8226
rect 2106 8227 2107 8228
rect 2178 8227 2179 8228
rect 2112 8229 2113 8230
rect 2160 8229 2161 8230
rect 1580 8231 1581 8232
rect 2160 8231 2161 8232
rect 2124 8233 2125 8234
rect 2196 8233 2197 8234
rect 2130 8235 2131 8236
rect 2184 8235 2185 8236
rect 2136 8237 2137 8238
rect 3023 8237 3024 8238
rect 2142 8239 2143 8240
rect 2190 8239 2191 8240
rect 1426 8241 1427 8242
rect 2190 8241 2191 8242
rect 2148 8243 2149 8244
rect 2172 8243 2173 8244
rect 2154 8245 2155 8246
rect 2652 8245 2653 8246
rect 2166 8247 2167 8248
rect 3202 8247 3203 8248
rect 2166 8249 2167 8250
rect 2268 8249 2269 8250
rect 2172 8251 2173 8252
rect 2214 8251 2215 8252
rect 1435 8253 1436 8254
rect 2214 8253 2215 8254
rect 2178 8255 2179 8256
rect 2520 8255 2521 8256
rect 2184 8257 2185 8258
rect 2202 8257 2203 8258
rect 2196 8259 2197 8260
rect 2220 8259 2221 8260
rect 2202 8261 2203 8262
rect 2514 8261 2515 8262
rect 2208 8263 2209 8264
rect 2292 8263 2293 8264
rect 2220 8265 2221 8266
rect 2226 8265 2227 8266
rect 2226 8267 2227 8268
rect 2232 8267 2233 8268
rect 2229 8269 2230 8270
rect 2235 8269 2236 8270
rect 2232 8271 2233 8272
rect 2238 8271 2239 8272
rect 2238 8273 2239 8274
rect 2244 8273 2245 8274
rect 2244 8275 2245 8276
rect 2250 8275 2251 8276
rect 2250 8277 2251 8278
rect 2256 8277 2257 8278
rect 2256 8279 2257 8280
rect 2262 8279 2263 8280
rect 2262 8281 2263 8282
rect 2502 8281 2503 8282
rect 2268 8283 2269 8284
rect 2274 8283 2275 8284
rect 2271 8285 2272 8286
rect 2277 8285 2278 8286
rect 1442 8287 1443 8288
rect 2277 8287 2278 8288
rect 2274 8289 2275 8290
rect 2286 8289 2287 8290
rect 2280 8291 2281 8292
rect 2286 8291 2287 8292
rect 1515 8293 1516 8294
rect 2280 8293 2281 8294
rect 2283 8293 2284 8294
rect 2289 8293 2290 8294
rect 2292 8293 2293 8294
rect 2304 8293 2305 8294
rect 2298 8295 2299 8296
rect 2304 8295 2305 8296
rect 2298 8297 2299 8298
rect 2418 8297 2419 8298
rect 2313 8299 2314 8300
rect 2331 8299 2332 8300
rect 2316 8301 2317 8302
rect 3069 8301 3070 8302
rect 2316 8303 2317 8304
rect 2364 8303 2365 8304
rect 2319 8305 2320 8306
rect 3075 8305 3076 8306
rect 2322 8307 2323 8308
rect 2442 8307 2443 8308
rect 1605 8309 1606 8310
rect 2442 8309 2443 8310
rect 2337 8311 2338 8312
rect 2349 8311 2350 8312
rect 2295 8313 2296 8314
rect 2337 8313 2338 8314
rect 2346 8313 2347 8314
rect 2358 8313 2359 8314
rect 2334 8315 2335 8316
rect 2346 8315 2347 8316
rect 1470 8317 1471 8318
rect 2334 8317 2335 8318
rect 2352 8317 2353 8318
rect 2364 8317 2365 8318
rect 2340 8319 2341 8320
rect 2352 8319 2353 8320
rect 2340 8321 2341 8322
rect 2376 8321 2377 8322
rect 2370 8323 2371 8324
rect 2394 8323 2395 8324
rect 2376 8325 2377 8326
rect 2400 8325 2401 8326
rect 2382 8327 2383 8328
rect 2394 8327 2395 8328
rect 2382 8329 2383 8330
rect 2550 8329 2551 8330
rect 2400 8331 2401 8332
rect 2490 8331 2491 8332
rect 2418 8333 2419 8334
rect 2430 8333 2431 8334
rect 2424 8335 2425 8336
rect 2430 8335 2431 8336
rect 2412 8337 2413 8338
rect 2424 8337 2425 8338
rect 2412 8339 2413 8340
rect 3147 8339 3148 8340
rect 2454 8341 2455 8342
rect 2466 8341 2467 8342
rect 2466 8343 2467 8344
rect 2556 8343 2557 8344
rect 2490 8345 2491 8346
rect 2508 8345 2509 8346
rect 2496 8347 2497 8348
rect 2956 8347 2957 8348
rect 2496 8349 2497 8350
rect 2562 8349 2563 8350
rect 2502 8351 2503 8352
rect 2574 8351 2575 8352
rect 2508 8353 2509 8354
rect 2526 8353 2527 8354
rect 2514 8355 2515 8356
rect 2568 8355 2569 8356
rect 2520 8357 2521 8358
rect 2532 8357 2533 8358
rect 2526 8359 2527 8360
rect 2538 8359 2539 8360
rect 2532 8361 2533 8362
rect 2598 8361 2599 8362
rect 2538 8363 2539 8364
rect 3180 8363 3181 8364
rect 2544 8365 2545 8366
rect 3020 8365 3021 8366
rect 2544 8367 2545 8368
rect 2592 8367 2593 8368
rect 2550 8369 2551 8370
rect 2616 8369 2617 8370
rect 2556 8371 2557 8372
rect 2610 8371 2611 8372
rect 2562 8373 2563 8374
rect 2580 8373 2581 8374
rect 2568 8375 2569 8376
rect 2586 8375 2587 8376
rect 2574 8377 2575 8378
rect 2622 8377 2623 8378
rect 2586 8379 2587 8380
rect 2604 8379 2605 8380
rect 2592 8381 2593 8382
rect 2628 8381 2629 8382
rect 2604 8383 2605 8384
rect 2640 8383 2641 8384
rect 2610 8385 2611 8386
rect 2646 8385 2647 8386
rect 2616 8387 2617 8388
rect 2658 8387 2659 8388
rect 2622 8389 2623 8390
rect 2670 8389 2671 8390
rect 2628 8391 2629 8392
rect 2664 8391 2665 8392
rect 2640 8393 2641 8394
rect 2694 8393 2695 8394
rect 2646 8395 2647 8396
rect 2700 8395 2701 8396
rect 2652 8397 2653 8398
rect 2706 8397 2707 8398
rect 2658 8399 2659 8400
rect 2736 8399 2737 8400
rect 2664 8401 2665 8402
rect 2742 8401 2743 8402
rect 1746 8403 1747 8404
rect 2742 8403 2743 8404
rect 1746 8405 1747 8406
rect 1872 8405 1873 8406
rect 1872 8407 1873 8408
rect 1956 8407 1957 8408
rect 1956 8409 1957 8410
rect 2718 8409 2719 8410
rect 2670 8411 2671 8412
rect 2724 8411 2725 8412
rect 2682 8413 2683 8414
rect 2748 8413 2749 8414
rect 2694 8415 2695 8416
rect 2796 8415 2797 8416
rect 2700 8417 2701 8418
rect 2802 8417 2803 8418
rect 2706 8419 2707 8420
rect 2808 8419 2809 8420
rect 2724 8421 2725 8422
rect 2826 8421 2827 8422
rect 2733 8423 2734 8424
rect 2835 8423 2836 8424
rect 2736 8425 2737 8426
rect 2850 8425 2851 8426
rect 1517 8427 1518 8428
rect 2850 8427 2851 8428
rect 1449 8429 1450 8430
rect 1518 8429 1519 8430
rect 2748 8429 2749 8430
rect 2862 8429 2863 8430
rect 2751 8431 2752 8432
rect 2865 8431 2866 8432
rect 2754 8433 2755 8434
rect 2868 8433 2869 8434
rect 2769 8435 2770 8436
rect 3209 8435 3210 8436
rect 2772 8437 2773 8438
rect 2844 8437 2845 8438
rect 2775 8439 2776 8440
rect 2838 8439 2839 8440
rect 2784 8441 2785 8442
rect 2886 8441 2887 8442
rect 2796 8443 2797 8444
rect 2910 8443 2911 8444
rect 2802 8445 2803 8446
rect 3126 8445 3127 8446
rect 2808 8447 2809 8448
rect 2922 8447 2923 8448
rect 2826 8449 2827 8450
rect 2940 8449 2941 8450
rect 2829 8451 2830 8452
rect 2943 8451 2944 8452
rect 2832 8453 2833 8454
rect 3173 8453 3174 8454
rect 2832 8455 2833 8456
rect 2970 8455 2971 8456
rect 2838 8457 2839 8458
rect 2946 8457 2947 8458
rect 2856 8459 2857 8460
rect 3066 8459 3067 8460
rect 2856 8461 2857 8462
rect 2976 8461 2977 8462
rect 2862 8463 2863 8464
rect 2874 8463 2875 8464
rect 2874 8465 2875 8466
rect 3000 8465 3001 8466
rect 2883 8467 2884 8468
rect 3205 8467 3206 8468
rect 2898 8469 2899 8470
rect 3166 8469 3167 8470
rect 2898 8471 2899 8472
rect 3012 8471 3013 8472
rect 2598 8473 2599 8474
rect 3011 8473 3012 8474
rect 2901 8475 2902 8476
rect 3015 8475 3016 8476
rect 2910 8477 2911 8478
rect 3018 8477 3019 8478
rect 2916 8479 2917 8480
rect 3177 8479 3178 8480
rect 2916 8481 2917 8482
rect 3033 8481 3034 8482
rect 2712 8483 2713 8484
rect 3034 8483 3035 8484
rect 2712 8485 2713 8486
rect 2814 8485 2815 8486
rect 2814 8487 2815 8488
rect 2928 8487 2929 8488
rect 2919 8489 2920 8490
rect 2994 8489 2995 8490
rect 2928 8491 2929 8492
rect 3048 8491 3049 8492
rect 2931 8493 2932 8494
rect 2964 8493 2965 8494
rect 2934 8495 2935 8496
rect 3063 8495 3064 8496
rect 2937 8497 2938 8498
rect 2949 8497 2950 8498
rect 2940 8499 2941 8500
rect 3072 8499 3073 8500
rect 2730 8501 2731 8502
rect 3072 8501 3073 8502
rect 1644 8503 1645 8504
rect 2730 8503 2731 8504
rect 1644 8505 1645 8506
rect 1710 8505 1711 8506
rect 1680 8507 1681 8508
rect 1710 8507 1711 8508
rect 1680 8509 1681 8510
rect 2367 8509 2368 8510
rect 2355 8511 2356 8512
rect 2367 8511 2368 8512
rect 2946 8511 2947 8512
rect 3060 8511 3061 8512
rect 2952 8513 2953 8514
rect 3068 8513 3069 8514
rect 2406 8515 2407 8516
rect 2953 8515 2954 8516
rect 2388 8517 2389 8518
rect 2406 8517 2407 8518
rect 2388 8519 2389 8520
rect 2436 8519 2437 8520
rect 2436 8521 2437 8522
rect 3144 8521 3145 8522
rect 2958 8523 2959 8524
rect 3065 8523 3066 8524
rect 2959 8525 2960 8526
rect 3084 8525 3085 8526
rect 2971 8527 2972 8528
rect 3123 8527 3124 8528
rect 2986 8529 2987 8530
rect 3001 8529 3002 8530
rect 2995 8531 2996 8532
rect 3151 8531 3152 8532
rect 2998 8533 2999 8534
rect 3141 8533 3142 8534
rect 3004 8535 3005 8536
rect 3120 8535 3121 8536
rect 3006 8537 3007 8538
rect 3081 8537 3082 8538
rect 2982 8539 2983 8540
rect 3082 8539 3083 8540
rect 3009 8541 3010 8542
rect 3129 8541 3130 8542
rect 2634 8543 2635 8544
rect 3008 8543 3009 8544
rect 2634 8545 2635 8546
rect 2676 8545 2677 8546
rect 1770 8547 1771 8548
rect 2676 8547 2677 8548
rect 1770 8549 1771 8550
rect 1938 8549 1939 8550
rect 1938 8551 1939 8552
rect 1986 8551 1987 8552
rect 1986 8553 1987 8554
rect 2766 8553 2767 8554
rect 2766 8555 2767 8556
rect 2880 8555 2881 8556
rect 2880 8557 2881 8558
rect 2988 8557 2989 8558
rect 3014 8557 3015 8558
rect 3157 8557 3158 8558
rect 3017 8559 3018 8560
rect 3160 8559 3161 8560
rect 3027 8561 3028 8562
rect 3096 8561 3097 8562
rect 3036 8563 3037 8564
rect 3212 8563 3213 8564
rect 2983 8565 2984 8566
rect 3037 8565 3038 8566
rect 3044 8565 3045 8566
rect 3114 8565 3115 8566
rect 3047 8567 3048 8568
rect 3199 8567 3200 8568
rect 3059 8569 3060 8570
rect 3078 8569 3079 8570
rect 2688 8571 2689 8572
rect 3079 8571 3080 8572
rect 2688 8573 2689 8574
rect 2790 8573 2791 8574
rect 2790 8575 2791 8576
rect 2904 8575 2905 8576
rect 2904 8577 2905 8578
rect 3163 8577 3164 8578
rect 3062 8579 3063 8580
rect 3196 8579 3197 8580
rect 3108 8581 3109 8582
rect 3187 8581 3188 8582
rect 3138 8583 3139 8584
rect 3154 8583 3155 8584
rect 1423 8592 1424 8593
rect 2184 8592 2185 8593
rect 1423 8594 1424 8595
rect 2004 8594 2005 8595
rect 1426 8596 1427 8597
rect 1680 8596 1681 8597
rect 1426 8598 1427 8599
rect 1998 8598 1999 8599
rect 1430 8600 1431 8601
rect 2188 8600 2189 8601
rect 1430 8602 1431 8603
rect 2226 8602 2227 8603
rect 1433 8604 1434 8605
rect 2229 8604 2230 8605
rect 1437 8606 1438 8607
rect 2232 8606 2233 8607
rect 1440 8608 1441 8609
rect 1444 8608 1445 8609
rect 1444 8610 1445 8611
rect 1656 8610 1657 8611
rect 1447 8612 1448 8613
rect 1758 8612 1759 8613
rect 1433 8614 1434 8615
rect 1447 8614 1448 8615
rect 1451 8614 1452 8615
rect 1692 8614 1693 8615
rect 1451 8616 1452 8617
rect 1770 8616 1771 8617
rect 1454 8618 1455 8619
rect 1693 8618 1694 8619
rect 1454 8620 1455 8621
rect 1776 8620 1777 8621
rect 1461 8622 1462 8623
rect 2733 8622 2734 8623
rect 1466 8624 1467 8625
rect 1800 8624 1801 8625
rect 1470 8626 1471 8627
rect 2358 8626 2359 8627
rect 1470 8628 1471 8629
rect 1938 8628 1939 8629
rect 1473 8630 1474 8631
rect 1939 8630 1940 8631
rect 1473 8632 1474 8633
rect 2244 8632 2245 8633
rect 1458 8634 1459 8635
rect 2245 8634 2246 8635
rect 1494 8636 1495 8637
rect 1500 8636 1501 8637
rect 1488 8638 1489 8639
rect 1494 8638 1495 8639
rect 1512 8638 1513 8639
rect 1980 8638 1981 8639
rect 1506 8640 1507 8641
rect 1512 8640 1513 8641
rect 1506 8642 1507 8643
rect 3037 8642 3038 8643
rect 1515 8644 1516 8645
rect 1534 8644 1535 8645
rect 1524 8646 1525 8647
rect 1746 8646 1747 8647
rect 1531 8648 1532 8649
rect 1962 8648 1963 8649
rect 1543 8650 1544 8651
rect 1566 8650 1567 8651
rect 1552 8652 1553 8653
rect 1884 8652 1885 8653
rect 1560 8654 1561 8655
rect 1567 8654 1568 8655
rect 1554 8656 1555 8657
rect 1561 8656 1562 8657
rect 1584 8656 1585 8657
rect 1597 8656 1598 8657
rect 1588 8658 1589 8659
rect 1627 8658 1628 8659
rect 1602 8660 1603 8661
rect 1609 8660 1610 8661
rect 1620 8660 1621 8661
rect 2266 8660 2267 8661
rect 1614 8662 1615 8663
rect 1621 8662 1622 8663
rect 1644 8662 1645 8663
rect 1657 8662 1658 8663
rect 1638 8664 1639 8665
rect 1645 8664 1646 8665
rect 1674 8664 1675 8665
rect 1681 8664 1682 8665
rect 1668 8666 1669 8667
rect 1675 8666 1676 8667
rect 1662 8668 1663 8669
rect 1669 8668 1670 8669
rect 1650 8670 1651 8671
rect 1663 8670 1664 8671
rect 1585 8672 1586 8673
rect 1651 8672 1652 8673
rect 1722 8672 1723 8673
rect 1747 8672 1748 8673
rect 1723 8674 1724 8675
rect 1734 8674 1735 8675
rect 1716 8676 1717 8677
rect 1735 8676 1736 8677
rect 1717 8678 1718 8679
rect 1728 8678 1729 8679
rect 1729 8680 1730 8681
rect 2730 8680 2731 8681
rect 1740 8682 1741 8683
rect 1801 8682 1802 8683
rect 1741 8684 1742 8685
rect 1752 8684 1753 8685
rect 1527 8686 1528 8687
rect 1753 8686 1754 8687
rect 1527 8688 1528 8689
rect 2289 8688 2290 8689
rect 1759 8690 1760 8691
rect 1782 8690 1783 8691
rect 1764 8692 1765 8693
rect 1771 8692 1772 8693
rect 1765 8694 1766 8695
rect 1788 8694 1789 8695
rect 1463 8696 1464 8697
rect 1789 8696 1790 8697
rect 1777 8698 1778 8699
rect 1794 8698 1795 8699
rect 1783 8700 1784 8701
rect 1806 8700 1807 8701
rect 1795 8702 1796 8703
rect 1818 8702 1819 8703
rect 1807 8704 1808 8705
rect 1824 8704 1825 8705
rect 1819 8706 1820 8707
rect 1830 8706 1831 8707
rect 1825 8708 1826 8709
rect 1854 8708 1855 8709
rect 1831 8710 1832 8711
rect 1908 8710 1909 8711
rect 1848 8712 1849 8713
rect 2975 8712 2976 8713
rect 1849 8714 1850 8715
rect 1866 8714 1867 8715
rect 1855 8716 1856 8717
rect 1878 8716 1879 8717
rect 1867 8718 1868 8719
rect 1896 8718 1897 8719
rect 1879 8720 1880 8721
rect 1902 8720 1903 8721
rect 1894 8722 1895 8723
rect 1914 8722 1915 8723
rect 1897 8724 1898 8725
rect 2676 8724 2677 8725
rect 1903 8726 1904 8727
rect 1926 8726 1927 8727
rect 1909 8728 1910 8729
rect 1932 8728 1933 8729
rect 1915 8730 1916 8731
rect 1944 8730 1945 8731
rect 1921 8732 1922 8733
rect 1950 8732 1951 8733
rect 1927 8734 1928 8735
rect 1956 8734 1957 8735
rect 1933 8736 1934 8737
rect 1974 8736 1975 8737
rect 1945 8738 1946 8739
rect 1968 8738 1969 8739
rect 1951 8740 1952 8741
rect 2010 8740 2011 8741
rect 1957 8742 1958 8743
rect 1992 8742 1993 8743
rect 1963 8744 1964 8745
rect 2028 8744 2029 8745
rect 1969 8746 1970 8747
rect 2016 8746 2017 8747
rect 1975 8748 1976 8749
rect 2022 8748 2023 8749
rect 1981 8750 1982 8751
rect 2923 8750 2924 8751
rect 1993 8752 1994 8753
rect 2064 8752 2065 8753
rect 1572 8754 1573 8755
rect 2065 8754 2066 8755
rect 1548 8756 1549 8757
rect 1573 8756 1574 8757
rect 1549 8758 1550 8759
rect 1812 8758 1813 8759
rect 1813 8760 1814 8761
rect 1842 8760 1843 8761
rect 1843 8762 1844 8763
rect 1860 8762 1861 8763
rect 1861 8764 1862 8765
rect 1890 8764 1891 8765
rect 1999 8764 2000 8765
rect 2040 8764 2041 8765
rect 2005 8766 2006 8767
rect 2046 8766 2047 8767
rect 2011 8768 2012 8769
rect 2052 8768 2053 8769
rect 2014 8770 2015 8771
rect 2055 8770 2056 8771
rect 2017 8772 2018 8773
rect 2058 8772 2059 8773
rect 2023 8774 2024 8775
rect 2034 8774 2035 8775
rect 2029 8776 2030 8777
rect 2106 8776 2107 8777
rect 2032 8778 2033 8779
rect 2361 8778 2362 8779
rect 2035 8780 2036 8781
rect 2076 8780 2077 8781
rect 2041 8782 2042 8783
rect 2082 8782 2083 8783
rect 2047 8784 2048 8785
rect 2094 8784 2095 8785
rect 2053 8786 2054 8787
rect 2100 8786 2101 8787
rect 2059 8788 2060 8789
rect 2088 8788 2089 8789
rect 2070 8790 2071 8791
rect 2101 8790 2102 8791
rect 2071 8792 2072 8793
rect 2112 8792 2113 8793
rect 2077 8794 2078 8795
rect 2118 8794 2119 8795
rect 2083 8796 2084 8797
rect 2646 8796 2647 8797
rect 2089 8798 2090 8799
rect 2130 8798 2131 8799
rect 2095 8800 2096 8801
rect 2136 8800 2137 8801
rect 1440 8802 1441 8803
rect 2137 8802 2138 8803
rect 2107 8804 2108 8805
rect 2142 8804 2143 8805
rect 2113 8806 2114 8807
rect 2160 8806 2161 8807
rect 2119 8808 2120 8809
rect 2166 8808 2167 8809
rect 2124 8810 2125 8811
rect 2131 8810 2132 8811
rect 2125 8812 2126 8813
rect 2148 8812 2149 8813
rect 2143 8814 2144 8815
rect 2178 8814 2179 8815
rect 2149 8816 2150 8817
rect 2616 8816 2617 8817
rect 2161 8818 2162 8819
rect 2196 8818 2197 8819
rect 2167 8820 2168 8821
rect 2190 8820 2191 8821
rect 2179 8822 2180 8823
rect 2322 8822 2323 8823
rect 2185 8824 2186 8825
rect 2214 8824 2215 8825
rect 2191 8826 2192 8827
rect 2208 8826 2209 8827
rect 2197 8828 2198 8829
rect 2256 8828 2257 8829
rect 2202 8830 2203 8831
rect 3011 8830 3012 8831
rect 2203 8832 2204 8833
rect 2280 8832 2281 8833
rect 2209 8834 2210 8835
rect 2298 8834 2299 8835
rect 2215 8836 2216 8837
rect 2466 8836 2467 8837
rect 2227 8838 2228 8839
rect 2310 8838 2311 8839
rect 2233 8840 2234 8841
rect 2292 8840 2293 8841
rect 1593 8842 1594 8843
rect 2293 8842 2294 8843
rect 2250 8844 2251 8845
rect 3044 8844 3045 8845
rect 2251 8846 2252 8847
rect 2268 8846 2269 8847
rect 2254 8848 2255 8849
rect 2271 8848 2272 8849
rect 2257 8850 2258 8851
rect 2274 8850 2275 8851
rect 2260 8852 2261 8853
rect 2277 8852 2278 8853
rect 2262 8854 2263 8855
rect 2852 8854 2853 8855
rect 2263 8856 2264 8857
rect 2286 8856 2287 8857
rect 2269 8858 2270 8859
rect 2502 8858 2503 8859
rect 2275 8860 2276 8861
rect 2442 8860 2443 8861
rect 2281 8862 2282 8863
rect 2316 8862 2317 8863
rect 1575 8864 1576 8865
rect 2317 8864 2318 8865
rect 2287 8866 2288 8867
rect 2304 8866 2305 8867
rect 2299 8868 2300 8869
rect 2956 8868 2957 8869
rect 2305 8870 2306 8871
rect 2334 8870 2335 8871
rect 2308 8872 2309 8873
rect 2337 8872 2338 8873
rect 2311 8874 2312 8875
rect 2328 8874 2329 8875
rect 2314 8876 2315 8877
rect 2331 8876 2332 8877
rect 2319 8878 2320 8879
rect 2356 8878 2357 8879
rect 2323 8880 2324 8881
rect 2346 8880 2347 8881
rect 2326 8882 2327 8883
rect 2349 8882 2350 8883
rect 2329 8884 2330 8885
rect 2340 8884 2341 8885
rect 2335 8886 2336 8887
rect 2352 8886 2353 8887
rect 2341 8888 2342 8889
rect 2364 8888 2365 8889
rect 2344 8890 2345 8891
rect 2367 8890 2368 8891
rect 2347 8892 2348 8893
rect 2388 8892 2389 8893
rect 2353 8894 2354 8895
rect 2961 8894 2962 8895
rect 2359 8896 2360 8897
rect 2370 8896 2371 8897
rect 2365 8898 2366 8899
rect 2376 8898 2377 8899
rect 2371 8900 2372 8901
rect 2394 8900 2395 8901
rect 2377 8902 2378 8903
rect 2490 8902 2491 8903
rect 2389 8904 2390 8905
rect 2454 8904 2455 8905
rect 2395 8906 2396 8907
rect 2412 8906 2413 8907
rect 2400 8908 2401 8909
rect 2953 8908 2954 8909
rect 2401 8910 2402 8911
rect 2418 8910 2419 8911
rect 2413 8912 2414 8913
rect 2430 8912 2431 8913
rect 2419 8914 2420 8915
rect 2436 8914 2437 8915
rect 2431 8916 2432 8917
rect 2448 8916 2449 8917
rect 2437 8918 2438 8919
rect 2460 8918 2461 8919
rect 2443 8920 2444 8921
rect 2514 8920 2515 8921
rect 2449 8922 2450 8923
rect 2508 8922 2509 8923
rect 2455 8924 2456 8925
rect 2484 8924 2485 8925
rect 2461 8926 2462 8927
rect 2472 8926 2473 8927
rect 2467 8928 2468 8929
rect 2478 8928 2479 8929
rect 2473 8930 2474 8931
rect 2544 8930 2545 8931
rect 2479 8932 2480 8933
rect 2532 8932 2533 8933
rect 2485 8934 2486 8935
rect 2550 8934 2551 8935
rect 2491 8936 2492 8937
rect 2520 8936 2521 8937
rect 2496 8938 2497 8939
rect 3008 8938 3009 8939
rect 2497 8940 2498 8941
rect 2526 8940 2527 8941
rect 2503 8942 2504 8943
rect 2538 8942 2539 8943
rect 2509 8944 2510 8945
rect 2556 8944 2557 8945
rect 2515 8946 2516 8947
rect 2592 8946 2593 8947
rect 2521 8948 2522 8949
rect 2562 8948 2563 8949
rect 2527 8950 2528 8951
rect 2568 8950 2569 8951
rect 2533 8952 2534 8953
rect 2598 8952 2599 8953
rect 2536 8954 2537 8955
rect 2901 8954 2902 8955
rect 2539 8956 2540 8957
rect 2769 8956 2770 8957
rect 2545 8958 2546 8959
rect 2586 8958 2587 8959
rect 2551 8960 2552 8961
rect 2604 8960 2605 8961
rect 2557 8962 2558 8963
rect 2610 8962 2611 8963
rect 2563 8964 2564 8965
rect 2622 8964 2623 8965
rect 2569 8966 2570 8967
rect 2628 8966 2629 8967
rect 2574 8968 2575 8969
rect 3034 8968 3035 8969
rect 2575 8970 2576 8971
rect 2634 8970 2635 8971
rect 2581 8972 2582 8973
rect 2652 8972 2653 8973
rect 2593 8974 2594 8975
rect 2664 8974 2665 8975
rect 2605 8976 2606 8977
rect 3079 8976 3080 8977
rect 2611 8978 2612 8979
rect 2670 8978 2671 8979
rect 2617 8980 2618 8981
rect 2800 8980 2801 8981
rect 2620 8982 2621 8983
rect 2895 8982 2896 8983
rect 2623 8984 2624 8985
rect 2688 8984 2689 8985
rect 2629 8986 2630 8987
rect 2694 8986 2695 8987
rect 2635 8988 2636 8989
rect 2700 8988 2701 8989
rect 2653 8990 2654 8991
rect 2751 8990 2752 8991
rect 2656 8992 2657 8993
rect 2724 8992 2725 8993
rect 2658 8994 2659 8995
rect 3072 8994 3073 8995
rect 2659 8996 2660 8997
rect 2848 8996 2849 8997
rect 2665 8998 2666 8999
rect 2736 8998 2737 8999
rect 2671 9000 2672 9001
rect 2742 9000 2743 9001
rect 2677 9002 2678 9003
rect 2754 9002 2755 9003
rect 2695 9004 2696 9005
rect 2766 9004 2767 9005
rect 2698 9006 2699 9007
rect 3082 9006 3083 9007
rect 2701 9008 2702 9009
rect 2772 9008 2773 9009
rect 2704 9010 2705 9011
rect 2775 9010 2776 9011
rect 2719 9012 2720 9013
rect 2796 9012 2797 9013
rect 2722 9014 2723 9015
rect 2901 9014 2902 9015
rect 2725 9016 2726 9017
rect 2862 9016 2863 9017
rect 2731 9018 2732 9019
rect 2968 9018 2969 9019
rect 2737 9020 2738 9021
rect 2808 9020 2809 9021
rect 2743 9022 2744 9023
rect 2784 9022 2785 9023
rect 2761 9024 2762 9025
rect 2826 9024 2827 9025
rect 2764 9026 2765 9027
rect 2829 9026 2830 9027
rect 2767 9028 2768 9029
rect 2832 9028 2833 9029
rect 2773 9030 2774 9031
rect 2850 9030 2851 9031
rect 2785 9032 2786 9033
rect 2802 9032 2803 9033
rect 2797 9034 2798 9035
rect 2892 9034 2893 9035
rect 2818 9036 2819 9037
rect 2919 9036 2920 9037
rect 2332 9038 2333 9039
rect 2920 9038 2921 9039
rect 2821 9040 2822 9041
rect 2904 9040 2905 9041
rect 2682 9042 2683 9043
rect 2904 9042 2905 9043
rect 2683 9044 2684 9045
rect 2745 9044 2746 9045
rect 2827 9044 2828 9045
rect 2910 9044 2911 9045
rect 2833 9046 2834 9047
rect 2949 9046 2950 9047
rect 2836 9048 2837 9049
rect 2937 9048 2938 9049
rect 2790 9050 2791 9051
rect 2937 9050 2938 9051
rect 2838 9052 2839 9053
rect 3065 9052 3066 9053
rect 2839 9054 2840 9055
rect 2940 9054 2941 9055
rect 2845 9056 2846 9057
rect 3075 9056 3076 9057
rect 2856 9058 2857 9059
rect 2891 9058 2892 9059
rect 2220 9060 2221 9061
rect 2855 9060 2856 9061
rect 2221 9062 2222 9063
rect 2238 9062 2239 9063
rect 1524 9064 1525 9065
rect 2239 9064 2240 9065
rect 2858 9064 2859 9065
rect 2959 9064 2960 9065
rect 2748 9066 2749 9067
rect 2958 9066 2959 9067
rect 2749 9068 2750 9069
rect 2814 9068 2815 9069
rect 2815 9070 2816 9071
rect 3030 9070 3031 9071
rect 2870 9072 2871 9073
rect 2971 9072 2972 9073
rect 2712 9074 2713 9075
rect 2972 9074 2973 9075
rect 2880 9076 2881 9077
rect 3020 9076 3021 9077
rect 2882 9078 2883 9079
rect 3001 9078 3002 9079
rect 2885 9080 2886 9081
rect 2986 9080 2987 9081
rect 2888 9082 2889 9083
rect 2995 9082 2996 9083
rect 2894 9084 2895 9085
rect 2898 9084 2899 9085
rect 1836 9086 1837 9087
rect 2897 9086 2898 9087
rect 1437 9088 1438 9089
rect 1837 9088 1838 9089
rect 2907 9088 2908 9089
rect 3014 9088 3015 9089
rect 2910 9090 2911 9091
rect 3017 9090 3018 9091
rect 2913 9092 2914 9093
rect 3023 9092 3024 9093
rect 2916 9094 2917 9095
rect 3027 9094 3028 9095
rect 2154 9096 2155 9097
rect 2916 9096 2917 9097
rect 2155 9098 2156 9099
rect 2172 9098 2173 9099
rect 2173 9100 2174 9101
rect 2382 9100 2383 9101
rect 2383 9102 2384 9103
rect 2406 9102 2407 9103
rect 2407 9104 2408 9105
rect 2424 9104 2425 9105
rect 1590 9106 1591 9107
rect 2425 9106 2426 9107
rect 2928 9106 2929 9107
rect 3041 9106 3042 9107
rect 1986 9108 1987 9109
rect 2927 9108 2928 9109
rect 1987 9110 1988 9111
rect 2640 9110 2641 9111
rect 2641 9112 2642 9113
rect 2706 9112 2707 9113
rect 2707 9114 2708 9115
rect 2778 9114 2779 9115
rect 2931 9114 2932 9115
rect 3068 9114 3069 9115
rect 2587 9116 2588 9117
rect 2930 9116 2931 9117
rect 2934 9116 2935 9117
rect 2946 9116 2947 9117
rect 2874 9118 2875 9119
rect 2934 9118 2935 9119
rect 2940 9118 2941 9119
rect 3047 9118 3048 9119
rect 2952 9120 2953 9121
rect 3059 9120 3060 9121
rect 2955 9122 2956 9123
rect 3062 9122 3063 9123
rect 2965 9124 2966 9125
rect 2998 9124 2999 9125
rect 2983 9126 2984 9127
rect 3004 9126 3005 9127
rect 1426 9135 1427 9136
rect 1957 9135 1958 9136
rect 1426 9137 1427 9138
rect 2263 9137 2264 9138
rect 1430 9139 1431 9140
rect 1783 9139 1784 9140
rect 1430 9141 1431 9142
rect 2185 9141 2186 9142
rect 1437 9143 1438 9144
rect 2260 9143 2261 9144
rect 1440 9145 1441 9146
rect 1813 9145 1814 9146
rect 1444 9147 1445 9148
rect 2521 9147 2522 9148
rect 1444 9149 1445 9150
rect 2257 9149 2258 9150
rect 1451 9151 1452 9152
rect 2617 9151 2618 9152
rect 1458 9153 1459 9154
rect 2593 9153 2594 9154
rect 1458 9155 1459 9156
rect 2209 9155 2210 9156
rect 1461 9157 1462 9158
rect 2305 9157 2306 9158
rect 1461 9159 1462 9160
rect 1795 9159 1796 9160
rect 1470 9161 1471 9162
rect 1534 9161 1535 9162
rect 1470 9163 1471 9164
rect 2059 9163 2060 9164
rect 1473 9165 1474 9166
rect 2341 9165 2342 9166
rect 1473 9167 1474 9168
rect 2041 9167 2042 9168
rect 1531 9169 1532 9170
rect 1891 9169 1892 9170
rect 1531 9171 1532 9172
rect 2125 9171 2126 9172
rect 1534 9173 1535 9174
rect 1573 9173 1574 9174
rect 1537 9175 1538 9176
rect 1561 9175 1562 9176
rect 1543 9177 1544 9178
rect 1555 9177 1556 9178
rect 1543 9179 1544 9180
rect 1567 9179 1568 9180
rect 1549 9181 1550 9182
rect 1873 9181 1874 9182
rect 1552 9183 1553 9184
rect 1597 9183 1598 9184
rect 1564 9185 1565 9186
rect 1699 9185 1700 9186
rect 1576 9187 1577 9188
rect 2855 9187 2856 9188
rect 1585 9189 1586 9190
rect 2548 9189 2549 9190
rect 1588 9191 1589 9192
rect 2332 9191 2333 9192
rect 1603 9193 1604 9194
rect 1657 9193 1658 9194
rect 1609 9195 1610 9196
rect 1633 9195 1634 9196
rect 1609 9197 1610 9198
rect 1663 9197 1664 9198
rect 1437 9199 1438 9200
rect 1663 9199 1664 9200
rect 1615 9201 1616 9202
rect 1645 9201 1646 9202
rect 1621 9203 1622 9204
rect 1858 9203 1859 9204
rect 1621 9205 1622 9206
rect 1675 9205 1676 9206
rect 1627 9207 1628 9208
rect 2521 9207 2522 9208
rect 1627 9209 1628 9210
rect 1681 9209 1682 9210
rect 1639 9211 1640 9212
rect 1693 9211 1694 9212
rect 1645 9213 1646 9214
rect 1687 9213 1688 9214
rect 1657 9215 1658 9216
rect 1717 9215 1718 9216
rect 1675 9217 1676 9218
rect 1765 9217 1766 9218
rect 1681 9219 1682 9220
rect 1723 9219 1724 9220
rect 1687 9221 1688 9222
rect 1741 9221 1742 9222
rect 1693 9223 1694 9224
rect 1711 9223 1712 9224
rect 1423 9225 1424 9226
rect 1711 9225 1712 9226
rect 1423 9227 1424 9228
rect 2293 9227 2294 9228
rect 1717 9229 1718 9230
rect 2005 9229 2006 9230
rect 1723 9231 1724 9232
rect 2011 9231 2012 9232
rect 1726 9233 1727 9234
rect 2014 9233 2015 9234
rect 1741 9235 1742 9236
rect 1999 9235 2000 9236
rect 1747 9237 1748 9238
rect 2257 9237 2258 9238
rect 1747 9239 1748 9240
rect 2053 9239 2054 9240
rect 1765 9241 1766 9242
rect 2065 9241 2066 9242
rect 1777 9243 1778 9244
rect 2209 9243 2210 9244
rect 1777 9245 1778 9246
rect 2137 9245 2138 9246
rect 1783 9247 1784 9248
rect 1915 9247 1916 9248
rect 1795 9249 1796 9250
rect 2167 9249 2168 9250
rect 1798 9251 1799 9252
rect 2266 9251 2267 9252
rect 1813 9253 1814 9254
rect 2191 9253 2192 9254
rect 1825 9255 1826 9256
rect 2341 9255 2342 9256
rect 1825 9257 1826 9258
rect 2089 9257 2090 9258
rect 1846 9259 1847 9260
rect 2254 9259 2255 9260
rect 1852 9261 1853 9262
rect 2188 9261 2189 9262
rect 1873 9263 1874 9264
rect 2311 9263 2312 9264
rect 1885 9265 1886 9266
rect 2335 9265 2336 9266
rect 1888 9267 1889 9268
rect 2344 9267 2345 9268
rect 1894 9269 1895 9270
rect 2386 9269 2387 9270
rect 1903 9271 1904 9272
rect 2897 9271 2898 9272
rect 1524 9273 1525 9274
rect 1903 9273 1904 9274
rect 1440 9275 1441 9276
rect 1524 9275 1525 9276
rect 1915 9275 1916 9276
rect 2371 9275 2372 9276
rect 1927 9277 1928 9278
rect 2930 9277 2931 9278
rect 1927 9279 1928 9280
rect 2383 9279 2384 9280
rect 1933 9281 1934 9282
rect 2927 9281 2928 9282
rect 1933 9283 1934 9284
rect 2233 9283 2234 9284
rect 1957 9285 1958 9286
rect 2407 9285 2408 9286
rect 1999 9287 2000 9288
rect 2347 9287 2348 9288
rect 2005 9289 2006 9290
rect 2437 9289 2438 9290
rect 1735 9291 1736 9292
rect 2437 9291 2438 9292
rect 1735 9293 1736 9294
rect 2017 9293 2018 9294
rect 2011 9295 2012 9296
rect 2299 9295 2300 9296
rect 2017 9297 2018 9298
rect 2431 9297 2432 9298
rect 2023 9299 2024 9300
rect 2191 9299 2192 9300
rect 1433 9301 1434 9302
rect 2023 9301 2024 9302
rect 2032 9301 2033 9302
rect 2416 9301 2417 9302
rect 2041 9303 2042 9304
rect 2461 9303 2462 9304
rect 2053 9305 2054 9306
rect 2675 9305 2676 9306
rect 2059 9307 2060 9308
rect 2113 9307 2114 9308
rect 2029 9309 2030 9310
rect 2113 9309 2114 9310
rect 2029 9311 2030 9312
rect 2389 9311 2390 9312
rect 1849 9313 1850 9314
rect 2389 9313 2390 9314
rect 1849 9315 1850 9316
rect 2961 9315 2962 9316
rect 2065 9317 2066 9318
rect 2449 9317 2450 9318
rect 1897 9319 1898 9320
rect 2449 9319 2450 9320
rect 1897 9321 1898 9322
rect 2323 9321 2324 9322
rect 1819 9323 1820 9324
rect 2323 9323 2324 9324
rect 1819 9325 1820 9326
rect 2197 9325 2198 9326
rect 1789 9327 1790 9328
rect 2197 9327 2198 9328
rect 1789 9329 1790 9330
rect 2047 9329 2048 9330
rect 2083 9329 2084 9330
rect 2734 9329 2735 9330
rect 2083 9331 2084 9332
rect 2491 9331 2492 9332
rect 2089 9333 2090 9334
rect 2497 9333 2498 9334
rect 2098 9335 2099 9336
rect 2455 9335 2456 9336
rect 2101 9337 2102 9338
rect 2916 9337 2917 9338
rect 1969 9339 1970 9340
rect 2101 9339 2102 9340
rect 1969 9341 1970 9342
rect 2119 9341 2120 9342
rect 2119 9343 2120 9344
rect 2527 9343 2528 9344
rect 2125 9345 2126 9346
rect 2509 9345 2510 9346
rect 2131 9347 2132 9348
rect 2913 9347 2914 9348
rect 2095 9349 2096 9350
rect 2131 9349 2132 9350
rect 2095 9351 2096 9352
rect 2503 9351 2504 9352
rect 2137 9353 2138 9354
rect 2545 9353 2546 9354
rect 1651 9355 1652 9356
rect 2545 9355 2546 9356
rect 1651 9357 1652 9358
rect 1669 9357 1670 9358
rect 1669 9359 1670 9360
rect 1759 9359 1760 9360
rect 1759 9361 1760 9362
rect 2071 9361 2072 9362
rect 2071 9363 2072 9364
rect 2443 9363 2444 9364
rect 1573 9365 1574 9366
rect 2443 9365 2444 9366
rect 2143 9367 2144 9368
rect 2626 9367 2627 9368
rect 2143 9369 2144 9370
rect 2473 9369 2474 9370
rect 2149 9371 2150 9372
rect 2920 9371 2921 9372
rect 2107 9373 2108 9374
rect 2149 9373 2150 9374
rect 1939 9375 1940 9376
rect 2107 9375 2108 9376
rect 1939 9377 1940 9378
rect 2227 9377 2228 9378
rect 1945 9379 1946 9380
rect 2227 9379 2228 9380
rect 1945 9381 1946 9382
rect 2329 9381 2330 9382
rect 1951 9383 1952 9384
rect 2329 9383 2330 9384
rect 1951 9385 1952 9386
rect 2179 9385 2180 9386
rect 1993 9387 1994 9388
rect 2179 9387 2180 9388
rect 1993 9389 1994 9390
rect 2395 9389 2396 9390
rect 1843 9391 1844 9392
rect 2395 9391 2396 9392
rect 1843 9393 1844 9394
rect 2251 9393 2252 9394
rect 1771 9395 1772 9396
rect 2251 9395 2252 9396
rect 1454 9397 1455 9398
rect 1771 9397 1772 9398
rect 1454 9399 1455 9400
rect 1500 9399 1501 9400
rect 1451 9401 1452 9402
rect 1500 9401 1501 9402
rect 2161 9401 2162 9402
rect 2778 9401 2779 9402
rect 1921 9403 1922 9404
rect 2161 9403 2162 9404
rect 1921 9405 1922 9406
rect 2239 9405 2240 9406
rect 1561 9407 1562 9408
rect 2239 9407 2240 9408
rect 2164 9409 2165 9410
rect 2314 9409 2315 9410
rect 2167 9411 2168 9412
rect 2515 9411 2516 9412
rect 2173 9413 2174 9414
rect 2185 9413 2186 9414
rect 1837 9415 1838 9416
rect 2173 9415 2174 9416
rect 1837 9417 1838 9418
rect 2245 9417 2246 9418
rect 2200 9419 2201 9420
rect 2308 9419 2309 9420
rect 2212 9421 2213 9422
rect 2326 9421 2327 9422
rect 2215 9423 2216 9424
rect 2901 9423 2902 9424
rect 1855 9425 1856 9426
rect 2215 9425 2216 9426
rect 2233 9425 2234 9426
rect 2269 9425 2270 9426
rect 2155 9427 2156 9428
rect 2269 9427 2270 9428
rect 2155 9429 2156 9430
rect 2425 9429 2426 9430
rect 2245 9431 2246 9432
rect 2533 9431 2534 9432
rect 2293 9433 2294 9434
rect 2563 9433 2564 9434
rect 2299 9435 2300 9436
rect 2569 9435 2570 9436
rect 2305 9437 2306 9438
rect 2575 9437 2576 9438
rect 2311 9439 2312 9440
rect 2715 9439 2716 9440
rect 2317 9441 2318 9442
rect 2894 9441 2895 9442
rect 1801 9443 1802 9444
rect 2317 9443 2318 9444
rect 1433 9445 1434 9446
rect 1801 9445 1802 9446
rect 2335 9445 2336 9446
rect 2581 9445 2582 9446
rect 2347 9447 2348 9448
rect 2611 9447 2612 9448
rect 2356 9449 2357 9450
rect 2470 9449 2471 9450
rect 2359 9451 2360 9452
rect 2668 9451 2669 9452
rect 1831 9453 1832 9454
rect 2359 9453 2360 9454
rect 1831 9455 1832 9456
rect 2221 9455 2222 9456
rect 1753 9457 1754 9458
rect 2221 9457 2222 9458
rect 1753 9459 1754 9460
rect 2077 9459 2078 9460
rect 1527 9461 1528 9462
rect 2077 9461 2078 9462
rect 1527 9463 1528 9464
rect 2785 9463 2786 9464
rect 2371 9465 2372 9466
rect 2587 9465 2588 9466
rect 2383 9467 2384 9468
rect 2536 9467 2537 9468
rect 2407 9469 2408 9470
rect 2635 9469 2636 9470
rect 2419 9471 2420 9472
rect 2711 9471 2712 9472
rect 2419 9473 2420 9474
rect 2623 9473 2624 9474
rect 2425 9475 2426 9476
rect 2641 9475 2642 9476
rect 2431 9477 2432 9478
rect 2904 9477 2905 9478
rect 2455 9479 2456 9480
rect 2659 9479 2660 9480
rect 2461 9481 2462 9482
rect 2848 9481 2849 9482
rect 2467 9483 2468 9484
rect 2972 9483 2973 9484
rect 1705 9485 1706 9486
rect 2467 9485 2468 9486
rect 1705 9487 1706 9488
rect 1867 9487 1868 9488
rect 1867 9489 1868 9490
rect 2287 9489 2288 9490
rect 2473 9489 2474 9490
rect 2695 9489 2696 9490
rect 2476 9491 2477 9492
rect 2698 9491 2699 9492
rect 2485 9493 2486 9494
rect 2741 9493 2742 9494
rect 2485 9495 2486 9496
rect 2671 9495 2672 9496
rect 2497 9497 2498 9498
rect 2719 9497 2720 9498
rect 1963 9499 1964 9500
rect 2718 9499 2719 9500
rect 1963 9501 1964 9502
rect 2281 9501 2282 9502
rect 1981 9503 1982 9504
rect 2281 9503 2282 9504
rect 1447 9505 1448 9506
rect 1981 9505 1982 9506
rect 1447 9507 1448 9508
rect 1855 9507 1856 9508
rect 2500 9507 2501 9508
rect 2722 9507 2723 9508
rect 2515 9509 2516 9510
rect 2701 9509 2702 9510
rect 2518 9511 2519 9512
rect 2704 9511 2705 9512
rect 2527 9513 2528 9514
rect 2731 9513 2732 9514
rect 2263 9515 2264 9516
rect 2730 9515 2731 9516
rect 2533 9517 2534 9518
rect 2965 9517 2966 9518
rect 2539 9519 2540 9520
rect 2852 9519 2853 9520
rect 1729 9521 1730 9522
rect 2539 9521 2540 9522
rect 1729 9523 1730 9524
rect 1861 9523 1862 9524
rect 1861 9525 1862 9526
rect 2035 9525 2036 9526
rect 2035 9527 2036 9528
rect 2377 9527 2378 9528
rect 1909 9529 1910 9530
rect 2377 9529 2378 9530
rect 1909 9531 1910 9532
rect 2353 9531 2354 9532
rect 1879 9533 1880 9534
rect 2353 9533 2354 9534
rect 1879 9535 1880 9536
rect 2203 9535 2204 9536
rect 2551 9535 2552 9536
rect 2672 9535 2673 9536
rect 2551 9537 2552 9538
rect 2751 9537 2752 9538
rect 2557 9539 2558 9540
rect 2727 9539 2728 9540
rect 2563 9541 2564 9542
rect 2761 9541 2762 9542
rect 2566 9543 2567 9544
rect 2764 9543 2765 9544
rect 2569 9545 2570 9546
rect 2749 9545 2750 9546
rect 2575 9547 2576 9548
rect 2767 9547 2768 9548
rect 2581 9549 2582 9550
rect 2773 9549 2774 9550
rect 2593 9551 2594 9552
rect 2743 9551 2744 9552
rect 2479 9553 2480 9554
rect 2744 9553 2745 9554
rect 2479 9555 2480 9556
rect 2677 9555 2678 9556
rect 2599 9557 2600 9558
rect 2707 9557 2708 9558
rect 2401 9559 2402 9560
rect 2708 9559 2709 9560
rect 2401 9561 2402 9562
rect 2629 9561 2630 9562
rect 2605 9563 2606 9564
rect 2748 9563 2749 9564
rect 2605 9565 2606 9566
rect 2725 9565 2726 9566
rect 2611 9567 2612 9568
rect 2800 9567 2801 9568
rect 2614 9569 2615 9570
rect 2683 9569 2684 9570
rect 2620 9571 2621 9572
rect 2797 9571 2798 9572
rect 2635 9573 2636 9574
rect 2815 9573 2816 9574
rect 2638 9575 2639 9576
rect 2818 9575 2819 9576
rect 2641 9577 2642 9578
rect 2821 9577 2822 9578
rect 2647 9579 2648 9580
rect 2827 9579 2828 9580
rect 2653 9581 2654 9582
rect 2937 9581 2938 9582
rect 2653 9583 2654 9584
rect 2833 9583 2834 9584
rect 2656 9585 2657 9586
rect 2934 9585 2935 9586
rect 2656 9587 2657 9588
rect 2836 9587 2837 9588
rect 2659 9589 2660 9590
rect 2839 9589 2840 9590
rect 2665 9591 2666 9592
rect 2845 9591 2846 9592
rect 2365 9593 2366 9594
rect 2665 9593 2666 9594
rect 2678 9593 2679 9594
rect 2870 9593 2871 9594
rect 2696 9595 2697 9596
rect 2882 9595 2883 9596
rect 2699 9597 2700 9598
rect 2885 9597 2886 9598
rect 2702 9599 2703 9600
rect 2888 9599 2889 9600
rect 2705 9601 2706 9602
rect 2891 9601 2892 9602
rect 2721 9603 2722 9604
rect 2907 9603 2908 9604
rect 2724 9605 2725 9606
rect 2910 9605 2911 9606
rect 2737 9607 2738 9608
rect 2968 9607 2969 9608
rect 1987 9609 1988 9610
rect 2737 9609 2738 9610
rect 1987 9611 1988 9612
rect 2275 9611 2276 9612
rect 1807 9613 1808 9614
rect 2275 9613 2276 9614
rect 1807 9615 1808 9616
rect 1975 9615 1976 9616
rect 1975 9617 1976 9618
rect 2413 9617 2414 9618
rect 2413 9619 2414 9620
rect 2623 9619 2624 9620
rect 2754 9619 2755 9620
rect 2940 9619 2941 9620
rect 2760 9621 2761 9622
rect 2955 9621 2956 9622
rect 2772 9623 2773 9624
rect 2958 9623 2959 9624
rect 2775 9625 2776 9626
rect 2952 9625 2953 9626
rect 2781 9627 2782 9628
rect 2975 9627 2976 9628
rect 2858 9629 2859 9630
rect 2923 9629 2924 9630
rect 1423 9638 1424 9639
rect 1518 9638 1519 9639
rect 1423 9640 1424 9641
rect 1615 9640 1616 9641
rect 1426 9642 1427 9643
rect 1831 9642 1832 9643
rect 1426 9644 1427 9645
rect 2263 9644 2264 9645
rect 1430 9646 1431 9647
rect 1777 9646 1778 9647
rect 1430 9648 1431 9649
rect 2059 9648 2060 9649
rect 1433 9650 1434 9651
rect 2527 9650 2528 9651
rect 1433 9652 1434 9653
rect 2275 9652 2276 9653
rect 1437 9654 1438 9655
rect 1603 9654 1604 9655
rect 1437 9656 1438 9657
rect 1633 9656 1634 9657
rect 1440 9658 1441 9659
rect 1602 9658 1603 9659
rect 1440 9660 1441 9661
rect 2699 9660 2700 9661
rect 1444 9662 1445 9663
rect 1711 9662 1712 9663
rect 1444 9664 1445 9665
rect 2212 9664 2213 9665
rect 1447 9666 1448 9667
rect 1698 9666 1699 9667
rect 1447 9668 1448 9669
rect 1609 9668 1610 9669
rect 1451 9670 1452 9671
rect 1899 9670 1900 9671
rect 1454 9672 1455 9673
rect 2164 9672 2165 9673
rect 1456 9674 1457 9675
rect 1879 9674 1880 9675
rect 1458 9676 1459 9677
rect 1537 9676 1538 9677
rect 1459 9678 1460 9679
rect 2098 9678 2099 9679
rect 1463 9680 1464 9681
rect 1639 9680 1640 9681
rect 1466 9682 1467 9683
rect 1645 9682 1646 9683
rect 1473 9684 1474 9685
rect 1861 9684 1862 9685
rect 1481 9686 1482 9687
rect 1494 9686 1495 9687
rect 1487 9688 1488 9689
rect 1500 9688 1501 9689
rect 1493 9690 1494 9691
rect 1512 9690 1513 9691
rect 1496 9692 1497 9693
rect 1506 9692 1507 9693
rect 1499 9694 1500 9695
rect 1543 9694 1544 9695
rect 1511 9696 1512 9697
rect 2386 9696 2387 9697
rect 1518 9698 1519 9699
rect 2413 9698 2414 9699
rect 1524 9700 1525 9701
rect 2545 9700 2546 9701
rect 1527 9702 1528 9703
rect 1632 9702 1633 9703
rect 1566 9704 1567 9705
rect 1627 9704 1628 9705
rect 1573 9706 1574 9707
rect 2449 9706 2450 9707
rect 1572 9708 1573 9709
rect 1626 9708 1627 9709
rect 1578 9710 1579 9711
rect 1651 9710 1652 9711
rect 1590 9712 1591 9713
rect 1657 9712 1658 9713
rect 1521 9714 1522 9715
rect 1656 9714 1657 9715
rect 1596 9716 1597 9717
rect 1681 9716 1682 9717
rect 1611 9718 1612 9719
rect 2065 9718 2066 9719
rect 1614 9720 1615 9721
rect 1669 9720 1670 9721
rect 1638 9722 1639 9723
rect 1687 9722 1688 9723
rect 1644 9724 1645 9725
rect 1771 9724 1772 9725
rect 1650 9726 1651 9727
rect 2197 9726 2198 9727
rect 1663 9728 1664 9729
rect 2665 9728 2666 9729
rect 1662 9730 1663 9731
rect 1729 9730 1730 9731
rect 1668 9732 1669 9733
rect 1705 9732 1706 9733
rect 1680 9734 1681 9735
rect 1783 9734 1784 9735
rect 1686 9736 1687 9737
rect 2161 9736 2162 9737
rect 1693 9738 1694 9739
rect 2633 9738 2634 9739
rect 1692 9740 1693 9741
rect 2107 9740 2108 9741
rect 1704 9742 1705 9743
rect 1801 9742 1802 9743
rect 1710 9744 1711 9745
rect 2173 9744 2174 9745
rect 1726 9746 1727 9747
rect 1743 9746 1744 9747
rect 1728 9748 1729 9749
rect 2718 9748 2719 9749
rect 1753 9750 1754 9751
rect 1776 9750 1777 9751
rect 1747 9752 1748 9753
rect 1752 9752 1753 9753
rect 1741 9754 1742 9755
rect 1746 9754 1747 9755
rect 1723 9756 1724 9757
rect 1740 9756 1741 9757
rect 1722 9758 1723 9759
rect 1807 9758 1808 9759
rect 1759 9760 1760 9761
rect 1770 9760 1771 9761
rect 1735 9762 1736 9763
rect 1758 9762 1759 9763
rect 1717 9764 1718 9765
rect 1734 9764 1735 9765
rect 1716 9766 1717 9767
rect 2101 9766 2102 9767
rect 1798 9768 1799 9769
rect 1827 9768 1828 9769
rect 1800 9770 1801 9771
rect 2179 9770 2180 9771
rect 1806 9772 1807 9773
rect 2077 9772 2078 9773
rect 1830 9774 1831 9775
rect 1969 9774 1970 9775
rect 1843 9776 1844 9777
rect 1860 9776 1861 9777
rect 1819 9778 1820 9779
rect 1842 9778 1843 9779
rect 1461 9780 1462 9781
rect 1818 9780 1819 9781
rect 1846 9780 1847 9781
rect 1863 9780 1864 9781
rect 1858 9782 1859 9783
rect 1869 9782 1870 9783
rect 1867 9784 1868 9785
rect 1878 9784 1879 9785
rect 1855 9786 1856 9787
rect 1866 9786 1867 9787
rect 1837 9788 1838 9789
rect 1854 9788 1855 9789
rect 1836 9790 1837 9791
rect 2053 9790 2054 9791
rect 1888 9792 1889 9793
rect 1923 9792 1924 9793
rect 1852 9794 1853 9795
rect 1887 9794 1888 9795
rect 1851 9796 1852 9797
rect 2200 9796 2201 9797
rect 1921 9798 1922 9799
rect 2616 9798 2617 9799
rect 1885 9800 1886 9801
rect 1920 9800 1921 9801
rect 1849 9802 1850 9803
rect 1884 9802 1885 9803
rect 1813 9804 1814 9805
rect 1848 9804 1849 9805
rect 1812 9806 1813 9807
rect 1825 9806 1826 9807
rect 1795 9808 1796 9809
rect 1824 9808 1825 9809
rect 1789 9810 1790 9811
rect 1794 9810 1795 9811
rect 1470 9812 1471 9813
rect 1788 9812 1789 9813
rect 1968 9812 1969 9813
rect 2113 9812 2114 9813
rect 1981 9814 1982 9815
rect 2708 9814 2709 9815
rect 1980 9816 1981 9817
rect 2011 9816 2012 9817
rect 1987 9818 1988 9819
rect 2052 9818 2053 9819
rect 1957 9820 1958 9821
rect 1986 9820 1987 9821
rect 1927 9822 1928 9823
rect 1956 9822 1957 9823
rect 1903 9824 1904 9825
rect 1926 9824 1927 9825
rect 1902 9826 1903 9827
rect 2023 9826 2024 9827
rect 1993 9828 1994 9829
rect 2010 9828 2011 9829
rect 1992 9830 1993 9831
rect 2711 9830 2712 9831
rect 2005 9832 2006 9833
rect 2022 9832 2023 9833
rect 1951 9834 1952 9835
rect 2004 9834 2005 9835
rect 1915 9836 1916 9837
rect 1950 9836 1951 9837
rect 1897 9838 1898 9839
rect 1914 9838 1915 9839
rect 1873 9840 1874 9841
rect 1896 9840 1897 9841
rect 1531 9842 1532 9843
rect 1872 9842 1873 9843
rect 2029 9842 2030 9843
rect 2046 9842 2047 9843
rect 2035 9844 2036 9845
rect 2058 9844 2059 9845
rect 2041 9846 2042 9847
rect 2109 9846 2110 9847
rect 2017 9848 2018 9849
rect 2040 9848 2041 9849
rect 1999 9850 2000 9851
rect 2016 9850 2017 9851
rect 1975 9852 1976 9853
rect 1998 9852 1999 9853
rect 1963 9854 1964 9855
rect 1974 9854 1975 9855
rect 1945 9856 1946 9857
rect 1962 9856 1963 9857
rect 1939 9858 1940 9859
rect 1944 9858 1945 9859
rect 1909 9860 1910 9861
rect 1938 9860 1939 9861
rect 1891 9862 1892 9863
rect 1908 9862 1909 9863
rect 1534 9864 1535 9865
rect 1890 9864 1891 9865
rect 2071 9864 2072 9865
rect 2112 9864 2113 9865
rect 2070 9866 2071 9867
rect 2191 9866 2192 9867
rect 2073 9868 2074 9869
rect 2209 9868 2210 9869
rect 2076 9870 2077 9871
rect 2131 9870 2132 9871
rect 2083 9872 2084 9873
rect 2619 9872 2620 9873
rect 2082 9874 2083 9875
rect 2668 9874 2669 9875
rect 2095 9876 2096 9877
rect 2106 9876 2107 9877
rect 2089 9878 2090 9879
rect 2094 9878 2095 9879
rect 2088 9880 2089 9881
rect 2149 9880 2150 9881
rect 2100 9882 2101 9883
rect 2672 9882 2673 9883
rect 2125 9884 2126 9885
rect 2751 9884 2752 9885
rect 2124 9886 2125 9887
rect 2215 9886 2216 9887
rect 2130 9888 2131 9889
rect 2251 9888 2252 9889
rect 2133 9890 2134 9891
rect 2416 9890 2417 9891
rect 2148 9892 2149 9893
rect 2239 9892 2240 9893
rect 2155 9894 2156 9895
rect 2741 9894 2742 9895
rect 2137 9896 2138 9897
rect 2154 9896 2155 9897
rect 2119 9898 2120 9899
rect 2136 9898 2137 9899
rect 2118 9900 2119 9901
rect 2650 9900 2651 9901
rect 2160 9902 2161 9903
rect 2185 9902 2186 9903
rect 1564 9904 1565 9905
rect 2184 9904 2185 9905
rect 2167 9906 2168 9907
rect 2172 9906 2173 9907
rect 1561 9908 1562 9909
rect 2166 9908 2167 9909
rect 1560 9910 1561 9911
rect 1621 9910 1622 9911
rect 1620 9912 1621 9913
rect 1675 9912 1676 9913
rect 1608 9914 1609 9915
rect 1674 9914 1675 9915
rect 2178 9914 2179 9915
rect 2227 9914 2228 9915
rect 2190 9916 2191 9917
rect 2317 9916 2318 9917
rect 2196 9918 2197 9919
rect 2233 9918 2234 9919
rect 2202 9920 2203 9921
rect 2245 9920 2246 9921
rect 2208 9922 2209 9923
rect 2323 9922 2324 9923
rect 2214 9924 2215 9925
rect 2281 9924 2282 9925
rect 2221 9926 2222 9927
rect 2623 9926 2624 9927
rect 2034 9928 2035 9929
rect 2623 9928 2624 9929
rect 2220 9930 2221 9931
rect 2341 9930 2342 9931
rect 2226 9932 2227 9933
rect 2293 9932 2294 9933
rect 2232 9934 2233 9935
rect 2305 9934 2306 9935
rect 2238 9936 2239 9937
rect 2630 9936 2631 9937
rect 2250 9938 2251 9939
rect 2335 9938 2336 9939
rect 2257 9940 2258 9941
rect 2781 9940 2782 9941
rect 2256 9942 2257 9943
rect 2359 9942 2360 9943
rect 1514 9944 1515 9945
rect 2358 9944 2359 9945
rect 2262 9946 2263 9947
rect 2437 9946 2438 9947
rect 2269 9948 2270 9949
rect 2727 9948 2728 9949
rect 2268 9950 2269 9951
rect 2347 9950 2348 9951
rect 2274 9952 2275 9953
rect 2607 9952 2608 9953
rect 2280 9954 2281 9955
rect 2371 9954 2372 9955
rect 2286 9956 2287 9957
rect 2395 9956 2396 9957
rect 2299 9958 2300 9959
rect 2553 9958 2554 9959
rect 2298 9960 2299 9961
rect 2383 9960 2384 9961
rect 2301 9962 2302 9963
rect 2353 9962 2354 9963
rect 2304 9964 2305 9965
rect 2377 9964 2378 9965
rect 2311 9966 2312 9967
rect 2626 9966 2627 9967
rect 2310 9968 2311 9969
rect 2443 9968 2444 9969
rect 2316 9970 2317 9971
rect 2425 9970 2426 9971
rect 2322 9972 2323 9973
rect 2419 9972 2420 9973
rect 2329 9974 2330 9975
rect 2734 9974 2735 9975
rect 1576 9976 1577 9977
rect 2328 9976 2329 9977
rect 1575 9978 1576 9979
rect 2431 9978 2432 9979
rect 2334 9980 2335 9981
rect 2401 9980 2402 9981
rect 2346 9982 2347 9983
rect 2455 9982 2456 9983
rect 2352 9984 2353 9985
rect 2461 9984 2462 9985
rect 2364 9986 2365 9987
rect 2479 9986 2480 9987
rect 2370 9988 2371 9989
rect 2485 9988 2486 9989
rect 2382 9990 2383 9991
rect 2473 9990 2474 9991
rect 2385 9992 2386 9993
rect 2476 9992 2477 9993
rect 2394 9994 2395 9995
rect 2497 9994 2498 9995
rect 2397 9996 2398 9997
rect 2407 9996 2408 9997
rect 2400 9998 2401 9999
rect 2583 9998 2584 9999
rect 2412 10000 2413 10001
rect 2533 10000 2534 10001
rect 2418 10002 2419 10003
rect 2515 10002 2516 10003
rect 2421 10004 2422 10005
rect 2518 10004 2519 10005
rect 2424 10006 2425 10007
rect 2467 10006 2468 10007
rect 2427 10008 2428 10009
rect 2470 10008 2471 10009
rect 2430 10010 2431 10011
rect 2551 10010 2552 10011
rect 2028 10012 2029 10013
rect 2550 10012 2551 10013
rect 2442 10014 2443 10015
rect 2563 10014 2564 10015
rect 2445 10016 2446 10017
rect 2566 10016 2567 10017
rect 2454 10018 2455 10019
rect 2548 10018 2549 10019
rect 2457 10020 2458 10021
rect 2539 10020 2540 10021
rect 2460 10022 2461 10023
rect 2569 10022 2570 10023
rect 2466 10024 2467 10025
rect 2575 10024 2576 10025
rect 2472 10026 2473 10027
rect 2737 10026 2738 10027
rect 2478 10028 2479 10029
rect 2581 10028 2582 10029
rect 2490 10030 2491 10031
rect 2593 10030 2594 10031
rect 2496 10032 2497 10033
rect 2599 10032 2600 10033
rect 2500 10034 2501 10035
rect 2643 10034 2644 10035
rect 2502 10036 2503 10037
rect 2568 10036 2569 10037
rect 2508 10038 2509 10039
rect 2571 10038 2572 10039
rect 2526 10040 2527 10041
rect 2611 10040 2612 10041
rect 2529 10042 2530 10043
rect 2614 10042 2615 10043
rect 2532 10044 2533 10045
rect 2635 10044 2636 10045
rect 2535 10046 2536 10047
rect 2638 10046 2639 10047
rect 2544 10048 2545 10049
rect 2647 10048 2648 10049
rect 2521 10050 2522 10051
rect 2646 10050 2647 10051
rect 2556 10052 2557 10053
rect 2656 10052 2657 10053
rect 2559 10054 2560 10055
rect 2605 10054 2606 10055
rect 2389 10056 2390 10057
rect 2604 10056 2605 10057
rect 2388 10058 2389 10059
rect 2580 10058 2581 10059
rect 2574 10060 2575 10061
rect 2659 10060 2660 10061
rect 2592 10062 2593 10063
rect 2696 10062 2697 10063
rect 2595 10064 2596 10065
rect 2678 10064 2679 10065
rect 2598 10066 2599 10067
rect 2724 10066 2725 10067
rect 2601 10068 2602 10069
rect 2778 10068 2779 10069
rect 2610 10070 2611 10071
rect 2702 10070 2703 10071
rect 2613 10072 2614 10073
rect 2705 10072 2706 10073
rect 2626 10074 2627 10075
rect 2683 10074 2684 10075
rect 2637 10076 2638 10077
rect 2641 10076 2642 10077
rect 2538 10078 2539 10079
rect 2640 10078 2641 10079
rect 2656 10078 2657 10079
rect 2754 10078 2755 10079
rect 2662 10080 2663 10081
rect 2760 10080 2761 10081
rect 2668 10082 2669 10083
rect 2775 10082 2776 10083
rect 2675 10084 2676 10085
rect 2715 10084 2716 10085
rect 2680 10086 2681 10087
rect 2772 10086 2773 10087
rect 2721 10088 2722 10089
rect 2744 10088 2745 10089
rect 2730 10090 2731 10091
rect 2748 10090 2749 10091
rect 1423 10099 1424 10100
rect 1878 10099 1879 10100
rect 1426 10101 1427 10102
rect 1644 10101 1645 10102
rect 1430 10103 1431 10104
rect 2130 10103 2131 10104
rect 1429 10105 1430 10106
rect 1788 10105 1789 10106
rect 1433 10107 1434 10108
rect 1998 10107 1999 10108
rect 1432 10109 1433 10110
rect 1602 10109 1603 10110
rect 1437 10111 1438 10112
rect 1596 10111 1597 10112
rect 1436 10113 1437 10114
rect 1743 10113 1744 10114
rect 1440 10115 1441 10116
rect 1590 10115 1591 10116
rect 1439 10117 1440 10118
rect 1560 10117 1561 10118
rect 1447 10119 1448 10120
rect 1794 10119 1795 10120
rect 1446 10121 1447 10122
rect 1899 10121 1900 10122
rect 1459 10123 1460 10124
rect 2388 10123 2389 10124
rect 1463 10125 1464 10126
rect 2454 10125 2455 10126
rect 1462 10127 1463 10128
rect 1626 10127 1627 10128
rect 1466 10129 1467 10130
rect 2328 10129 2329 10130
rect 1465 10131 1466 10132
rect 1674 10131 1675 10132
rect 1481 10133 1482 10134
rect 2030 10133 2031 10134
rect 1480 10135 1481 10136
rect 1499 10135 1500 10136
rect 1487 10137 1488 10138
rect 2042 10137 2043 10138
rect 1486 10139 1487 10140
rect 1974 10139 1975 10140
rect 1489 10141 1490 10142
rect 1956 10141 1957 10142
rect 1493 10143 1494 10144
rect 2066 10143 2067 10144
rect 1496 10145 1497 10146
rect 1923 10145 1924 10146
rect 1498 10147 1499 10148
rect 2298 10147 2299 10148
rect 1501 10149 1502 10150
rect 2352 10149 2353 10150
rect 1505 10151 1506 10152
rect 1926 10151 1927 10152
rect 1508 10153 1509 10154
rect 2162 10153 2163 10154
rect 1511 10155 1512 10156
rect 1800 10155 1801 10156
rect 1514 10157 1515 10158
rect 2070 10157 2071 10158
rect 1518 10159 1519 10160
rect 1595 10159 1596 10160
rect 1521 10161 1522 10162
rect 1887 10161 1888 10162
rect 1523 10163 1524 10164
rect 1611 10163 1612 10164
rect 1535 10165 1536 10166
rect 1578 10165 1579 10166
rect 1541 10167 1542 10168
rect 1554 10167 1555 10168
rect 1553 10169 1554 10170
rect 2526 10169 2527 10170
rect 1556 10171 1557 10172
rect 2198 10171 2199 10172
rect 1566 10173 1567 10174
rect 1577 10173 1578 10174
rect 1568 10175 1569 10176
rect 2136 10175 2137 10176
rect 1572 10177 1573 10178
rect 2358 10177 2359 10178
rect 1458 10179 1459 10180
rect 1571 10179 1572 10180
rect 1575 10179 1576 10180
rect 2424 10179 2425 10180
rect 1583 10181 1584 10182
rect 1728 10181 1729 10182
rect 1589 10183 1590 10184
rect 2262 10183 2263 10184
rect 1601 10185 1602 10186
rect 1656 10185 1657 10186
rect 1620 10187 1621 10188
rect 1643 10187 1644 10188
rect 1619 10189 1620 10190
rect 1638 10189 1639 10190
rect 1614 10191 1615 10192
rect 1637 10191 1638 10192
rect 1613 10193 1614 10194
rect 1632 10193 1633 10194
rect 1650 10193 1651 10194
rect 1655 10193 1656 10194
rect 1649 10195 1650 10196
rect 2256 10195 2257 10196
rect 1664 10197 1665 10198
rect 2190 10197 2191 10198
rect 1673 10199 1674 10200
rect 2208 10199 2209 10200
rect 1680 10201 1681 10202
rect 2387 10201 2388 10202
rect 1679 10203 1680 10204
rect 2220 10203 2221 10204
rect 1686 10205 1687 10206
rect 1727 10205 1728 10206
rect 1722 10207 1723 10208
rect 1781 10207 1782 10208
rect 1721 10209 1722 10210
rect 2124 10209 2125 10210
rect 1734 10211 1735 10212
rect 1808 10211 1809 10212
rect 1733 10213 1734 10214
rect 2166 10213 2167 10214
rect 1787 10215 1788 10216
rect 2274 10215 2275 10216
rect 1793 10217 1794 10218
rect 2346 10217 2347 10218
rect 1827 10219 1828 10220
rect 1940 10219 1941 10220
rect 1832 10221 1833 10222
rect 2370 10221 2371 10222
rect 1836 10223 1837 10224
rect 1877 10223 1878 10224
rect 1764 10225 1765 10226
rect 1835 10225 1836 10226
rect 1698 10227 1699 10228
rect 1763 10227 1764 10228
rect 1697 10229 1698 10230
rect 2184 10229 2185 10230
rect 1848 10231 1849 10232
rect 1955 10231 1956 10232
rect 1776 10233 1777 10234
rect 1847 10233 1848 10234
rect 1716 10235 1717 10236
rect 1775 10235 1776 10236
rect 1668 10237 1669 10238
rect 1715 10237 1716 10238
rect 1851 10237 1852 10238
rect 1958 10237 1959 10238
rect 1854 10239 1855 10240
rect 1973 10239 1974 10240
rect 1853 10241 1854 10242
rect 2178 10241 2179 10242
rect 1863 10243 1864 10244
rect 1982 10243 1983 10244
rect 1869 10245 1870 10246
rect 2012 10245 2013 10246
rect 1920 10247 1921 10248
rect 2063 10247 2064 10248
rect 1925 10249 1926 10250
rect 2196 10249 2197 10250
rect 1932 10251 1933 10252
rect 2619 10251 2620 10252
rect 1931 10253 1932 10254
rect 2028 10253 2029 10254
rect 1884 10255 1885 10256
rect 2027 10255 2028 10256
rect 1883 10257 1884 10258
rect 1902 10257 1903 10258
rect 1901 10259 1902 10260
rect 2076 10259 2077 10260
rect 1938 10261 1939 10262
rect 2075 10261 2076 10262
rect 1824 10263 1825 10264
rect 1937 10263 1938 10264
rect 1752 10265 1753 10266
rect 1823 10265 1824 10266
rect 1444 10267 1445 10268
rect 1751 10267 1752 10268
rect 1443 10269 1444 10270
rect 2088 10269 2089 10270
rect 1950 10271 1951 10272
rect 2222 10271 2223 10272
rect 1872 10273 1873 10274
rect 1949 10273 1950 10274
rect 1812 10275 1813 10276
rect 1871 10275 1872 10276
rect 1746 10277 1747 10278
rect 1811 10277 1812 10278
rect 1704 10279 1705 10280
rect 1745 10279 1746 10280
rect 1703 10281 1704 10282
rect 2148 10281 2149 10282
rect 1952 10283 1953 10284
rect 2133 10283 2134 10284
rect 1997 10285 1998 10286
rect 2052 10285 2053 10286
rect 1914 10287 1915 10288
rect 2051 10287 2052 10288
rect 1818 10289 1819 10290
rect 1913 10289 1914 10290
rect 1758 10291 1759 10292
rect 1817 10291 1818 10292
rect 1757 10293 1758 10294
rect 2318 10293 2319 10294
rect 2016 10295 2017 10296
rect 2087 10295 2088 10296
rect 1908 10297 1909 10298
rect 2015 10297 2016 10298
rect 1907 10299 1908 10300
rect 2550 10299 2551 10300
rect 2024 10301 2025 10302
rect 2529 10301 2530 10302
rect 2034 10303 2035 10304
rect 2135 10303 2136 10304
rect 2033 10305 2034 10306
rect 2202 10305 2203 10306
rect 2040 10307 2041 10308
rect 2626 10307 2627 10308
rect 1896 10309 1897 10310
rect 2039 10309 2040 10310
rect 1895 10311 1896 10312
rect 2316 10311 2317 10312
rect 2046 10313 2047 10314
rect 2204 10313 2205 10314
rect 1608 10315 1609 10316
rect 2045 10315 2046 10316
rect 1565 10317 1566 10318
rect 1607 10317 1608 10318
rect 2054 10317 2055 10318
rect 2073 10317 2074 10318
rect 2058 10319 2059 10320
rect 2616 10319 2617 10320
rect 1962 10321 1963 10322
rect 2057 10321 2058 10322
rect 1842 10323 1843 10324
rect 1961 10323 1962 10324
rect 1770 10325 1771 10326
rect 1841 10325 1842 10326
rect 1769 10327 1770 10328
rect 2315 10327 2316 10328
rect 2060 10329 2061 10330
rect 2310 10329 2311 10330
rect 2069 10331 2070 10332
rect 2100 10331 2101 10332
rect 2078 10333 2079 10334
rect 2427 10333 2428 10334
rect 2082 10335 2083 10336
rect 2147 10335 2148 10336
rect 2081 10337 2082 10338
rect 2112 10337 2113 10338
rect 2010 10339 2011 10340
rect 2111 10339 2112 10340
rect 1456 10341 1457 10342
rect 2009 10341 2010 10342
rect 1455 10343 1456 10344
rect 1625 10343 1626 10344
rect 2094 10343 2095 10344
rect 2165 10343 2166 10344
rect 2093 10345 2094 10346
rect 2219 10345 2220 10346
rect 2106 10347 2107 10348
rect 2650 10347 2651 10348
rect 1992 10349 1993 10350
rect 2105 10349 2106 10350
rect 1991 10351 1992 10352
rect 2623 10351 2624 10352
rect 2118 10353 2119 10354
rect 2123 10353 2124 10354
rect 1986 10355 1987 10356
rect 2117 10355 2118 10356
rect 1866 10357 1867 10358
rect 1985 10357 1986 10358
rect 1806 10359 1807 10360
rect 1865 10359 1866 10360
rect 1740 10361 1741 10362
rect 1805 10361 1806 10362
rect 1692 10363 1693 10364
rect 1739 10363 1740 10364
rect 1691 10365 1692 10366
rect 1710 10365 1711 10366
rect 1662 10367 1663 10368
rect 1709 10367 1710 10368
rect 2129 10367 2130 10368
rect 2160 10367 2161 10368
rect 2154 10369 2155 10370
rect 2186 10369 2187 10370
rect 2153 10371 2154 10372
rect 2390 10371 2391 10372
rect 2159 10373 2160 10374
rect 2214 10373 2215 10374
rect 2168 10375 2169 10376
rect 2322 10375 2323 10376
rect 2172 10377 2173 10378
rect 2630 10377 2631 10378
rect 2174 10379 2175 10380
rect 2226 10379 2227 10380
rect 2180 10381 2181 10382
rect 2232 10381 2233 10382
rect 2192 10383 2193 10384
rect 2250 10383 2251 10384
rect 2201 10385 2202 10386
rect 2400 10385 2401 10386
rect 2207 10387 2208 10388
rect 2304 10387 2305 10388
rect 2225 10389 2226 10390
rect 2268 10389 2269 10390
rect 2231 10391 2232 10392
rect 2502 10391 2503 10392
rect 2238 10393 2239 10394
rect 2424 10393 2425 10394
rect 2243 10395 2244 10396
rect 2460 10395 2461 10396
rect 2249 10397 2250 10398
rect 2382 10397 2383 10398
rect 2252 10399 2253 10400
rect 2385 10399 2386 10400
rect 2255 10401 2256 10402
rect 2434 10401 2435 10402
rect 2261 10403 2262 10404
rect 2462 10403 2463 10404
rect 2267 10405 2268 10406
rect 2412 10405 2413 10406
rect 2273 10407 2274 10408
rect 2472 10407 2473 10408
rect 2286 10409 2287 10410
rect 2607 10409 2608 10410
rect 2291 10411 2292 10412
rect 2442 10411 2443 10412
rect 2294 10413 2295 10414
rect 2445 10413 2446 10414
rect 2022 10415 2023 10416
rect 2445 10415 2446 10416
rect 1980 10417 1981 10418
rect 2021 10417 2022 10418
rect 1860 10419 1861 10420
rect 1979 10419 1980 10420
rect 1859 10421 1860 10422
rect 1968 10421 1969 10422
rect 1967 10423 1968 10424
rect 2004 10423 2005 10424
rect 1944 10425 1945 10426
rect 2003 10425 2004 10426
rect 1890 10427 1891 10428
rect 1943 10427 1944 10428
rect 1830 10429 1831 10430
rect 1889 10429 1890 10430
rect 2297 10429 2298 10430
rect 2478 10429 2479 10430
rect 2301 10431 2302 10432
rect 2553 10431 2554 10432
rect 2309 10433 2310 10434
rect 2556 10433 2557 10434
rect 2312 10435 2313 10436
rect 2508 10435 2509 10436
rect 2321 10437 2322 10438
rect 2405 10437 2406 10438
rect 2334 10439 2335 10440
rect 2452 10439 2453 10440
rect 2333 10441 2334 10442
rect 2532 10441 2533 10442
rect 2336 10443 2337 10444
rect 2535 10443 2536 10444
rect 2339 10445 2340 10446
rect 2640 10445 2641 10446
rect 2345 10447 2346 10448
rect 2408 10447 2409 10448
rect 2351 10449 2352 10450
rect 2438 10449 2439 10450
rect 2357 10451 2358 10452
rect 2441 10451 2442 10452
rect 2364 10453 2365 10454
rect 2643 10453 2644 10454
rect 2369 10455 2370 10456
rect 2574 10455 2575 10456
rect 2375 10457 2376 10458
rect 2633 10457 2634 10458
rect 2381 10459 2382 10460
rect 2598 10459 2599 10460
rect 2384 10461 2385 10462
rect 2601 10461 2602 10462
rect 2394 10463 2395 10464
rect 2646 10463 2647 10464
rect 2397 10465 2398 10466
rect 2455 10465 2456 10466
rect 2399 10467 2400 10468
rect 2592 10467 2593 10468
rect 2402 10469 2403 10470
rect 2595 10469 2596 10470
rect 2411 10471 2412 10472
rect 2610 10471 2611 10472
rect 2414 10473 2415 10474
rect 2613 10473 2614 10474
rect 2418 10475 2419 10476
rect 2583 10475 2584 10476
rect 2109 10477 2110 10478
rect 2417 10477 2418 10478
rect 2421 10477 2422 10478
rect 2580 10477 2581 10478
rect 2280 10479 2281 10480
rect 2420 10479 2421 10480
rect 2279 10481 2280 10482
rect 2430 10481 2431 10482
rect 2427 10483 2428 10484
rect 2538 10483 2539 10484
rect 2431 10485 2432 10486
rect 2466 10485 2467 10486
rect 2448 10487 2449 10488
rect 2604 10487 2605 10488
rect 2457 10489 2458 10490
rect 2568 10489 2569 10490
rect 2459 10491 2460 10492
rect 2496 10491 2497 10492
rect 2465 10493 2466 10494
rect 2656 10493 2657 10494
rect 2471 10495 2472 10496
rect 2662 10495 2663 10496
rect 2477 10497 2478 10498
rect 2668 10497 2669 10498
rect 2490 10499 2491 10500
rect 2653 10499 2654 10500
rect 2489 10501 2490 10502
rect 2680 10501 2681 10502
rect 2492 10503 2493 10504
rect 2683 10503 2684 10504
rect 2544 10505 2545 10506
rect 2637 10505 2638 10506
rect 2559 10507 2560 10508
rect 2571 10507 2572 10508
rect 1429 10516 1430 10517
rect 1535 10516 1536 10517
rect 1432 10518 1433 10519
rect 2027 10518 2028 10519
rect 1436 10520 1437 10521
rect 1769 10520 1770 10521
rect 1439 10522 1440 10523
rect 1664 10522 1665 10523
rect 1441 10524 1442 10525
rect 1649 10524 1650 10525
rect 1443 10526 1444 10527
rect 2009 10526 2010 10527
rect 1444 10528 1445 10529
rect 1480 10528 1481 10529
rect 1448 10530 1449 10531
rect 1733 10530 1734 10531
rect 1451 10532 1452 10533
rect 1781 10532 1782 10533
rect 1455 10534 1456 10535
rect 1619 10534 1620 10535
rect 1455 10536 1456 10537
rect 1745 10536 1746 10537
rect 1458 10538 1459 10539
rect 1613 10538 1614 10539
rect 1465 10540 1466 10541
rect 1691 10540 1692 10541
rect 1467 10542 1468 10543
rect 1534 10542 1535 10543
rect 1470 10544 1471 10545
rect 2030 10544 2031 10545
rect 1479 10546 1480 10547
rect 1883 10546 1884 10547
rect 1482 10548 1483 10549
rect 1819 10548 1820 10549
rect 1486 10550 1487 10551
rect 2411 10550 2412 10551
rect 1486 10552 1487 10553
rect 1958 10552 1959 10553
rect 1489 10554 1490 10555
rect 1889 10554 1890 10555
rect 1489 10556 1490 10557
rect 1565 10556 1566 10557
rect 1498 10558 1499 10559
rect 2015 10558 2016 10559
rect 1498 10560 1499 10561
rect 1952 10560 1953 10561
rect 1505 10562 1506 10563
rect 1985 10562 1986 10563
rect 1504 10564 1505 10565
rect 1541 10564 1542 10565
rect 1510 10566 1511 10567
rect 1633 10566 1634 10567
rect 1523 10568 1524 10569
rect 1528 10568 1529 10569
rect 1462 10570 1463 10571
rect 1522 10570 1523 10571
rect 1537 10570 1538 10571
rect 1963 10570 1964 10571
rect 1553 10572 1554 10573
rect 1901 10572 1902 10573
rect 1552 10574 1553 10575
rect 2434 10574 2435 10575
rect 1556 10576 1557 10577
rect 2180 10576 2181 10577
rect 1558 10578 1559 10579
rect 2045 10578 2046 10579
rect 1561 10580 1562 10581
rect 1757 10580 1758 10581
rect 1568 10582 1569 10583
rect 2345 10582 2346 10583
rect 1577 10584 1578 10585
rect 1777 10584 1778 10585
rect 1576 10586 1577 10587
rect 1832 10586 1833 10587
rect 1612 10588 1613 10589
rect 1637 10588 1638 10589
rect 1618 10590 1619 10591
rect 1643 10590 1644 10591
rect 1630 10592 1631 10593
rect 2021 10592 2022 10593
rect 1651 10594 1652 10595
rect 1673 10594 1674 10595
rect 1655 10596 1656 10597
rect 2219 10596 2220 10597
rect 1654 10598 1655 10599
rect 2231 10598 2232 10599
rect 1660 10600 1661 10601
rect 1793 10600 1794 10601
rect 1666 10602 1667 10603
rect 2315 10602 2316 10603
rect 1672 10604 1673 10605
rect 1709 10604 1710 10605
rect 1684 10606 1685 10607
rect 1703 10606 1704 10607
rect 1446 10608 1447 10609
rect 1702 10608 1703 10609
rect 1690 10610 1691 10611
rect 1751 10610 1752 10611
rect 1708 10612 1709 10613
rect 1763 10612 1764 10613
rect 1727 10614 1728 10615
rect 2390 10614 2391 10615
rect 1697 10616 1698 10617
rect 1726 10616 1727 10617
rect 1732 10616 1733 10617
rect 1775 10616 1776 10617
rect 1735 10618 1736 10619
rect 2042 10618 2043 10619
rect 1750 10620 1751 10621
rect 1805 10620 1806 10621
rect 1753 10622 1754 10623
rect 1808 10622 1809 10623
rect 1756 10624 1757 10625
rect 1811 10624 1812 10625
rect 1762 10626 1763 10627
rect 1817 10626 1818 10627
rect 1774 10628 1775 10629
rect 1823 10628 1824 10629
rect 1780 10630 1781 10631
rect 2201 10630 2202 10631
rect 1789 10632 1790 10633
rect 1841 10632 1842 10633
rect 1795 10634 1796 10635
rect 1847 10634 1848 10635
rect 1801 10636 1802 10637
rect 1853 10636 1854 10637
rect 1807 10638 1808 10639
rect 1865 10638 1866 10639
rect 1813 10640 1814 10641
rect 1877 10640 1878 10641
rect 1831 10642 1832 10643
rect 2168 10642 2169 10643
rect 1835 10644 1836 10645
rect 1888 10644 1889 10645
rect 1843 10646 1844 10647
rect 1925 10646 1926 10647
rect 1849 10648 1850 10649
rect 1937 10648 1938 10649
rect 1852 10650 1853 10651
rect 1940 10650 1941 10651
rect 1855 10652 1856 10653
rect 1913 10652 1914 10653
rect 1859 10654 1860 10655
rect 2176 10654 2177 10655
rect 1861 10656 1862 10657
rect 1991 10656 1992 10657
rect 1867 10658 1868 10659
rect 2033 10658 2034 10659
rect 1871 10660 1872 10661
rect 2101 10660 2102 10661
rect 1873 10662 1874 10663
rect 1961 10662 1962 10663
rect 1876 10664 1877 10665
rect 2012 10664 2013 10665
rect 1879 10666 1880 10667
rect 1973 10666 1974 10667
rect 1885 10668 1886 10669
rect 1979 10668 1980 10669
rect 1891 10670 1892 10671
rect 1955 10670 1956 10671
rect 1895 10672 1896 10673
rect 2131 10672 2132 10673
rect 1739 10674 1740 10675
rect 1894 10674 1895 10675
rect 1738 10676 1739 10677
rect 1787 10676 1788 10677
rect 1897 10676 1898 10677
rect 2159 10676 2160 10677
rect 1903 10678 1904 10679
rect 1943 10678 1944 10679
rect 1907 10680 1908 10681
rect 2424 10680 2425 10681
rect 1458 10682 1459 10683
rect 1906 10682 1907 10683
rect 1909 10682 1910 10683
rect 2003 10682 2004 10683
rect 1915 10684 1916 10685
rect 1931 10684 1932 10685
rect 1921 10686 1922 10687
rect 1967 10686 1968 10687
rect 1924 10688 1925 10689
rect 2024 10688 2025 10689
rect 1927 10690 1928 10691
rect 2051 10690 2052 10691
rect 1930 10692 1931 10693
rect 2054 10692 2055 10693
rect 1936 10694 1937 10695
rect 2312 10694 2313 10695
rect 1939 10696 1940 10697
rect 2063 10696 2064 10697
rect 1942 10698 1943 10699
rect 2066 10698 2067 10699
rect 1945 10700 1946 10701
rect 2057 10700 2058 10701
rect 1501 10702 1502 10703
rect 2056 10702 2057 10703
rect 1949 10704 1950 10705
rect 2196 10704 2197 10705
rect 1679 10706 1680 10707
rect 1948 10706 1949 10707
rect 1678 10708 1679 10709
rect 1715 10708 1716 10709
rect 1508 10710 1509 10711
rect 1714 10710 1715 10711
rect 1951 10710 1952 10711
rect 2075 10710 2076 10711
rect 1954 10712 1955 10713
rect 2078 10712 2079 10713
rect 1957 10714 1958 10715
rect 2179 10714 2180 10715
rect 1969 10716 1970 10717
rect 2093 10716 2094 10717
rect 1972 10718 1973 10719
rect 2309 10718 2310 10719
rect 1975 10720 1976 10721
rect 2081 10720 2082 10721
rect 1982 10722 1983 10723
rect 2455 10722 2456 10723
rect 1981 10724 1982 10725
rect 2123 10724 2124 10725
rect 1987 10726 1988 10727
rect 2069 10726 2070 10727
rect 1993 10728 1994 10729
rect 2117 10728 2118 10729
rect 1997 10730 1998 10731
rect 2098 10730 2099 10731
rect 1999 10732 2000 10733
rect 2111 10732 2112 10733
rect 2002 10734 2003 10735
rect 2162 10734 2163 10735
rect 2005 10736 2006 10737
rect 2427 10736 2428 10737
rect 2011 10738 2012 10739
rect 2135 10738 2136 10739
rect 2017 10740 2018 10741
rect 2147 10740 2148 10741
rect 2029 10742 2030 10743
rect 2141 10742 2142 10743
rect 2039 10744 2040 10745
rect 2140 10744 2141 10745
rect 2041 10746 2042 10747
rect 2192 10746 2193 10747
rect 2047 10748 2048 10749
rect 2198 10748 2199 10749
rect 2060 10750 2061 10751
rect 2420 10750 2421 10751
rect 2062 10752 2063 10753
rect 2207 10752 2208 10753
rect 2068 10754 2069 10755
rect 2252 10754 2253 10755
rect 2071 10756 2072 10757
rect 2186 10756 2187 10757
rect 1601 10758 1602 10759
rect 2186 10758 2187 10759
rect 1600 10760 1601 10761
rect 1625 10760 1626 10761
rect 1607 10762 1608 10763
rect 1624 10762 1625 10763
rect 1595 10764 1596 10765
rect 1606 10764 1607 10765
rect 1589 10766 1590 10767
rect 1594 10766 1595 10767
rect 1583 10768 1584 10769
rect 1588 10768 1589 10769
rect 1571 10770 1572 10771
rect 1582 10770 1583 10771
rect 2074 10770 2075 10771
rect 2273 10770 2274 10771
rect 2080 10772 2081 10773
rect 2452 10772 2453 10773
rect 2083 10774 2084 10775
rect 2165 10774 2166 10775
rect 2087 10776 2088 10777
rect 2448 10776 2449 10777
rect 2086 10778 2087 10779
rect 2243 10778 2244 10779
rect 2092 10780 2093 10781
rect 2414 10780 2415 10781
rect 2095 10782 2096 10783
rect 2297 10782 2298 10783
rect 2105 10784 2106 10785
rect 2143 10784 2144 10785
rect 2110 10786 2111 10787
rect 2279 10786 2280 10787
rect 2122 10788 2123 10789
rect 2291 10788 2292 10789
rect 2125 10790 2126 10791
rect 2294 10790 2295 10791
rect 2129 10792 2130 10793
rect 2202 10792 2203 10793
rect 2128 10794 2129 10795
rect 2333 10794 2334 10795
rect 2134 10796 2135 10797
rect 2339 10796 2340 10797
rect 2146 10798 2147 10799
rect 2351 10798 2352 10799
rect 2153 10800 2154 10801
rect 2190 10800 2191 10801
rect 2158 10802 2159 10803
rect 2399 10802 2400 10803
rect 2161 10804 2162 10805
rect 2321 10804 2322 10805
rect 2164 10806 2165 10807
rect 2336 10806 2337 10807
rect 2167 10808 2168 10809
rect 2193 10808 2194 10809
rect 2170 10810 2171 10811
rect 2381 10810 2382 10811
rect 2174 10812 2175 10813
rect 2199 10812 2200 10813
rect 2173 10814 2174 10815
rect 2357 10814 2358 10815
rect 2183 10816 2184 10817
rect 2402 10816 2403 10817
rect 2204 10818 2205 10819
rect 2387 10818 2388 10819
rect 2205 10820 2206 10821
rect 2438 10820 2439 10821
rect 2208 10822 2209 10823
rect 2465 10822 2466 10823
rect 2220 10824 2221 10825
rect 2489 10824 2490 10825
rect 2222 10826 2223 10827
rect 2249 10826 2250 10827
rect 2223 10828 2224 10829
rect 2492 10828 2493 10829
rect 2225 10830 2226 10831
rect 2462 10830 2463 10831
rect 2226 10832 2227 10833
rect 2471 10832 2472 10833
rect 2229 10834 2230 10835
rect 2477 10834 2478 10835
rect 2255 10836 2256 10837
rect 2417 10836 2418 10837
rect 2261 10838 2262 10839
rect 2431 10838 2432 10839
rect 2267 10840 2268 10841
rect 2459 10840 2460 10841
rect 2318 10842 2319 10843
rect 2445 10842 2446 10843
rect 2369 10844 2370 10845
rect 2405 10844 2406 10845
rect 2375 10846 2376 10847
rect 2408 10846 2409 10847
rect 2384 10848 2385 10849
rect 2441 10848 2442 10849
rect 1423 10857 1424 10858
rect 1714 10857 1715 10858
rect 1426 10859 1427 10860
rect 1600 10859 1601 10860
rect 1430 10861 1431 10862
rect 1873 10861 1874 10862
rect 1433 10863 1434 10864
rect 1921 10863 1922 10864
rect 1437 10865 1438 10866
rect 1795 10865 1796 10866
rect 1441 10867 1442 10868
rect 1606 10867 1607 10868
rect 1440 10869 1441 10870
rect 1753 10869 1754 10870
rect 1444 10871 1445 10872
rect 1682 10871 1683 10872
rect 1444 10873 1445 10874
rect 1528 10873 1529 10874
rect 1451 10875 1452 10876
rect 1732 10875 1733 10876
rect 1450 10877 1451 10878
rect 1903 10877 1904 10878
rect 1453 10879 1454 10880
rect 2029 10879 2030 10880
rect 1458 10881 1459 10882
rect 1894 10881 1895 10882
rect 1448 10883 1449 10884
rect 1459 10883 1460 10884
rect 1447 10885 1448 10886
rect 1522 10885 1523 10886
rect 1462 10887 1463 10888
rect 1684 10887 1685 10888
rect 1467 10889 1468 10890
rect 1651 10889 1652 10890
rect 1470 10891 1471 10892
rect 1948 10891 1949 10892
rect 1477 10893 1478 10894
rect 2101 10893 2102 10894
rect 1479 10895 1480 10896
rect 1813 10895 1814 10896
rect 1482 10897 1483 10898
rect 1807 10897 1808 10898
rect 1486 10899 1487 10900
rect 1720 10899 1721 10900
rect 1489 10901 1490 10902
rect 1777 10901 1778 10902
rect 1489 10903 1490 10904
rect 1927 10903 1928 10904
rect 1496 10905 1497 10906
rect 1510 10905 1511 10906
rect 1498 10907 1499 10908
rect 1508 10907 1509 10908
rect 1499 10909 1500 10910
rect 1504 10909 1505 10910
rect 1511 10909 1512 10910
rect 1906 10909 1907 10910
rect 1514 10911 1515 10912
rect 1552 10911 1553 10912
rect 1520 10913 1521 10914
rect 1588 10913 1589 10914
rect 1526 10915 1527 10916
rect 1594 10915 1595 10916
rect 1532 10917 1533 10918
rect 1612 10917 1613 10918
rect 1537 10919 1538 10920
rect 1951 10919 1952 10920
rect 1538 10921 1539 10922
rect 1618 10921 1619 10922
rect 1544 10923 1545 10924
rect 1624 10923 1625 10924
rect 1550 10925 1551 10926
rect 1582 10925 1583 10926
rect 1558 10927 1559 10928
rect 1924 10927 1925 10928
rect 1561 10929 1562 10930
rect 1766 10929 1767 10930
rect 1568 10931 1569 10932
rect 1660 10931 1661 10932
rect 1586 10933 1587 10934
rect 1672 10933 1673 10934
rect 1592 10935 1593 10936
rect 1678 10935 1679 10936
rect 1595 10937 1596 10938
rect 1876 10937 1877 10938
rect 1598 10939 1599 10940
rect 1708 10939 1709 10940
rect 1604 10941 1605 10942
rect 1865 10941 1866 10942
rect 1622 10943 1623 10944
rect 1750 10943 1751 10944
rect 1625 10945 1626 10946
rect 1756 10945 1757 10946
rect 1630 10947 1631 10948
rect 2161 10947 2162 10948
rect 1631 10949 1632 10950
rect 1762 10949 1763 10950
rect 1576 10951 1577 10952
rect 1763 10951 1764 10952
rect 1577 10953 1578 10954
rect 1954 10953 1955 10954
rect 1633 10955 1634 10956
rect 2041 10955 2042 10956
rect 1534 10957 1535 10958
rect 1634 10957 1635 10958
rect 1637 10957 1638 10958
rect 1690 10957 1691 10958
rect 1643 10959 1644 10960
rect 1702 10959 1703 10960
rect 1661 10961 1662 10962
rect 1738 10961 1739 10962
rect 1673 10963 1674 10964
rect 1780 10963 1781 10964
rect 1455 10965 1456 10966
rect 1781 10965 1782 10966
rect 1456 10967 1457 10968
rect 1735 10967 1736 10968
rect 1676 10969 1677 10970
rect 2143 10969 2144 10970
rect 1688 10971 1689 10972
rect 1831 10971 1832 10972
rect 1694 10973 1695 10974
rect 1849 10973 1850 10974
rect 1697 10975 1698 10976
rect 1852 10975 1853 10976
rect 1712 10977 1713 10978
rect 1891 10977 1892 10978
rect 1715 10979 1716 10980
rect 1855 10979 1856 10980
rect 1724 10981 1725 10982
rect 1879 10981 1880 10982
rect 1726 10983 1727 10984
rect 1950 10983 1951 10984
rect 1730 10985 1731 10986
rect 1885 10985 1886 10986
rect 1733 10987 1734 10988
rect 1888 10987 1889 10988
rect 1736 10989 1737 10990
rect 1897 10989 1898 10990
rect 1742 10991 1743 10992
rect 1843 10991 1844 10992
rect 1748 10993 1749 10994
rect 1909 10993 1910 10994
rect 1654 10995 1655 10996
rect 1910 10995 1911 10996
rect 1655 10997 1656 10998
rect 1789 10997 1790 10998
rect 1754 10999 1755 11000
rect 1867 10999 1868 11000
rect 1760 11001 1761 11002
rect 1915 11001 1916 11002
rect 1769 11003 1770 11004
rect 1939 11003 1940 11004
rect 1666 11005 1667 11006
rect 1939 11005 1940 11006
rect 1772 11007 1773 11008
rect 1942 11007 1943 11008
rect 1774 11009 1775 11010
rect 2179 11009 2180 11010
rect 1492 11011 1493 11012
rect 1775 11011 1776 11012
rect 1778 11011 1779 11012
rect 1930 11011 1931 11012
rect 1787 11013 1788 11014
rect 1920 11013 1921 11014
rect 1790 11015 1791 11016
rect 2002 11015 2003 11016
rect 1793 11017 1794 11018
rect 1963 11017 1964 11018
rect 1799 11019 1800 11020
rect 1969 11019 1970 11020
rect 1801 11021 1802 11022
rect 1953 11021 1954 11022
rect 1805 11023 1806 11024
rect 2183 11023 2184 11024
rect 1811 11025 1812 11026
rect 1975 11025 1976 11026
rect 1817 11027 1818 11028
rect 1981 11027 1982 11028
rect 1819 11029 1820 11030
rect 2140 11029 2141 11030
rect 1823 11031 1824 11032
rect 1987 11031 1988 11032
rect 1829 11033 1830 11034
rect 2011 11033 2012 11034
rect 1835 11035 1836 11036
rect 2005 11035 2006 11036
rect 1841 11037 1842 11038
rect 2199 11037 2200 11038
rect 1847 11039 1848 11040
rect 2056 11039 2057 11040
rect 1859 11041 1860 11042
rect 2047 11041 2048 11042
rect 1861 11043 1862 11044
rect 1913 11043 1914 11044
rect 1574 11045 1575 11046
rect 1862 11045 1863 11046
rect 1868 11045 1869 11046
rect 2071 11045 2072 11046
rect 1877 11047 1878 11048
rect 2092 11047 2093 11048
rect 1880 11049 1881 11050
rect 2095 11049 2096 11050
rect 1883 11051 1884 11052
rect 1972 11051 1973 11052
rect 1886 11053 1887 11054
rect 1936 11053 1937 11054
rect 1889 11055 1890 11056
rect 2128 11055 2129 11056
rect 1892 11057 1893 11058
rect 2131 11057 2132 11058
rect 1895 11059 1896 11060
rect 2122 11059 2123 11060
rect 1904 11061 1905 11062
rect 2158 11061 2159 11062
rect 1907 11063 1908 11064
rect 2167 11063 2168 11064
rect 1917 11065 1918 11066
rect 1957 11065 1958 11066
rect 1923 11067 1924 11068
rect 2170 11067 2171 11068
rect 1926 11069 1927 11070
rect 2146 11069 2147 11070
rect 1929 11071 1930 11072
rect 2086 11071 2087 11072
rect 1932 11073 1933 11074
rect 2074 11073 2075 11074
rect 1936 11075 1937 11076
rect 1945 11075 1946 11076
rect 1853 11077 1854 11078
rect 1946 11077 1947 11078
rect 1943 11079 1944 11080
rect 2062 11079 2063 11080
rect 1956 11081 1957 11082
rect 2110 11081 2111 11082
rect 1959 11083 1960 11084
rect 2125 11083 2126 11084
rect 1993 11085 1994 11086
rect 2176 11085 2177 11086
rect 1999 11087 2000 11088
rect 2186 11087 2187 11088
rect 2017 11089 2018 11090
rect 2193 11089 2194 11090
rect 2068 11091 2069 11092
rect 2098 11091 2099 11092
rect 2080 11093 2081 11094
rect 2205 11093 2206 11094
rect 2083 11095 2084 11096
rect 2196 11095 2197 11096
rect 2134 11097 2135 11098
rect 2202 11097 2203 11098
rect 2164 11099 2165 11100
rect 2208 11099 2209 11100
rect 2173 11101 2174 11102
rect 2190 11101 2191 11102
rect 2220 11101 2221 11102
rect 2229 11101 2230 11102
rect 2223 11103 2224 11104
rect 2226 11103 2227 11104
rect 1423 11112 1424 11113
rect 1604 11112 1605 11113
rect 1426 11114 1427 11115
rect 1598 11114 1599 11115
rect 1430 11116 1431 11117
rect 1534 11116 1535 11117
rect 1429 11118 1430 11119
rect 1631 11118 1632 11119
rect 1433 11120 1434 11121
rect 1748 11120 1749 11121
rect 1432 11122 1433 11123
rect 1763 11122 1764 11123
rect 1437 11124 1438 11125
rect 1655 11124 1656 11125
rect 1436 11126 1437 11127
rect 1772 11126 1773 11127
rect 1440 11128 1441 11129
rect 1733 11128 1734 11129
rect 1439 11130 1440 11131
rect 1538 11130 1539 11131
rect 1444 11132 1445 11133
rect 1477 11132 1478 11133
rect 1443 11134 1444 11135
rect 1532 11134 1533 11135
rect 1447 11136 1448 11137
rect 1595 11136 1596 11137
rect 1446 11138 1447 11139
rect 1592 11138 1593 11139
rect 1450 11140 1451 11141
rect 1622 11140 1623 11141
rect 1450 11142 1451 11143
rect 1715 11142 1716 11143
rect 1453 11144 1454 11145
rect 1712 11144 1713 11145
rect 1453 11146 1454 11147
rect 1787 11146 1788 11147
rect 1459 11148 1460 11149
rect 1643 11148 1644 11149
rect 1462 11150 1463 11151
rect 1637 11150 1638 11151
rect 1465 11152 1466 11153
rect 1694 11152 1695 11153
rect 1468 11154 1469 11155
rect 1625 11154 1626 11155
rect 1471 11156 1472 11157
rect 1634 11156 1635 11157
rect 1474 11158 1475 11159
rect 1586 11158 1587 11159
rect 1483 11160 1484 11161
rect 1730 11160 1731 11161
rect 1486 11162 1487 11163
rect 1724 11162 1725 11163
rect 1489 11164 1490 11165
rect 1883 11164 1884 11165
rect 1489 11166 1490 11167
rect 1697 11166 1698 11167
rect 1492 11168 1493 11169
rect 1835 11168 1836 11169
rect 1492 11170 1493 11171
rect 1917 11170 1918 11171
rect 1496 11172 1497 11173
rect 1508 11172 1509 11173
rect 1495 11174 1496 11175
rect 1778 11174 1779 11175
rect 1499 11176 1500 11177
rect 1511 11176 1512 11177
rect 1498 11178 1499 11179
rect 1769 11178 1770 11179
rect 1501 11180 1502 11181
rect 1544 11180 1545 11181
rect 1504 11182 1505 11183
rect 1526 11182 1527 11183
rect 1507 11184 1508 11185
rect 1520 11184 1521 11185
rect 1514 11186 1515 11187
rect 1519 11186 1520 11187
rect 1513 11188 1514 11189
rect 1550 11188 1551 11189
rect 1525 11190 1526 11191
rect 1760 11190 1761 11191
rect 1546 11192 1547 11193
rect 1907 11192 1908 11193
rect 1555 11194 1556 11195
rect 1829 11194 1830 11195
rect 1561 11196 1562 11197
rect 1754 11196 1755 11197
rect 1564 11198 1565 11199
rect 1790 11198 1791 11199
rect 1568 11200 1569 11201
rect 1603 11200 1604 11201
rect 1574 11202 1575 11203
rect 1585 11202 1586 11203
rect 1573 11204 1574 11205
rect 1823 11204 1824 11205
rect 1577 11206 1578 11207
rect 1588 11206 1589 11207
rect 1576 11208 1577 11209
rect 1793 11208 1794 11209
rect 1579 11210 1580 11211
rect 1886 11210 1887 11211
rect 1582 11212 1583 11213
rect 1799 11212 1800 11213
rect 1597 11214 1598 11215
rect 1892 11214 1893 11215
rect 1600 11216 1601 11217
rect 1676 11216 1677 11217
rect 1606 11218 1607 11219
rect 1805 11218 1806 11219
rect 1609 11220 1610 11221
rect 1736 11220 1737 11221
rect 1612 11222 1613 11223
rect 1661 11222 1662 11223
rect 1616 11224 1617 11225
rect 1817 11224 1818 11225
rect 1619 11226 1620 11227
rect 1811 11226 1812 11227
rect 1623 11228 1624 11229
rect 1688 11228 1689 11229
rect 1626 11230 1627 11231
rect 1682 11230 1683 11231
rect 1629 11232 1630 11233
rect 1775 11232 1776 11233
rect 1632 11234 1633 11235
rect 1868 11234 1869 11235
rect 1673 11236 1674 11237
rect 1953 11236 1954 11237
rect 1742 11238 1743 11239
rect 1913 11238 1914 11239
rect 1766 11240 1767 11241
rect 1865 11240 1866 11241
rect 1781 11242 1782 11243
rect 1946 11242 1947 11243
rect 1841 11244 1842 11245
rect 1939 11244 1940 11245
rect 1847 11246 1848 11247
rect 1943 11246 1944 11247
rect 1853 11248 1854 11249
rect 1862 11248 1863 11249
rect 1859 11250 1860 11251
rect 1950 11250 1951 11251
rect 1877 11252 1878 11253
rect 1932 11252 1933 11253
rect 1880 11254 1881 11255
rect 1929 11254 1930 11255
rect 1889 11256 1890 11257
rect 1910 11256 1911 11257
rect 1895 11258 1896 11259
rect 1956 11258 1957 11259
rect 1904 11260 1905 11261
rect 1920 11260 1921 11261
rect 1923 11260 1924 11261
rect 1959 11260 1960 11261
rect 1926 11262 1927 11263
rect 1936 11262 1937 11263
rect 1429 11271 1430 11272
rect 1468 11271 1469 11272
rect 1432 11273 1433 11274
rect 1471 11273 1472 11274
rect 1436 11275 1437 11276
rect 1483 11275 1484 11276
rect 1439 11277 1440 11278
rect 1486 11277 1487 11278
rect 1443 11279 1444 11280
rect 1456 11279 1457 11280
rect 1446 11281 1447 11282
rect 1474 11281 1475 11282
rect 1450 11283 1451 11284
rect 1555 11283 1556 11284
rect 1453 11285 1454 11286
rect 1525 11285 1526 11286
rect 1465 11287 1466 11288
rect 1629 11287 1630 11288
rect 1477 11289 1478 11290
rect 1519 11289 1520 11290
rect 1480 11291 1481 11292
rect 1534 11291 1535 11292
rect 1489 11293 1490 11294
rect 1498 11293 1499 11294
rect 1489 11295 1490 11296
rect 1585 11295 1586 11296
rect 1492 11297 1493 11298
rect 1495 11297 1496 11298
rect 1492 11299 1493 11300
rect 1588 11299 1589 11300
rect 1501 11301 1502 11302
rect 1507 11301 1508 11302
rect 1504 11303 1505 11304
rect 1513 11303 1514 11304
rect 1546 11303 1547 11304
rect 1603 11303 1604 11304
rect 1561 11305 1562 11306
rect 1632 11305 1633 11306
rect 1564 11307 1565 11308
rect 1609 11307 1610 11308
rect 1573 11309 1574 11310
rect 1619 11309 1620 11310
rect 1576 11311 1577 11312
rect 1616 11311 1617 11312
rect 1579 11313 1580 11314
rect 1612 11313 1613 11314
rect 1582 11315 1583 11316
rect 1606 11315 1607 11316
rect 1597 11317 1598 11318
rect 1626 11317 1627 11318
rect 1600 11319 1601 11320
rect 1623 11319 1624 11320
rect 1477 11328 1478 11329
rect 1492 11328 1493 11329
rect 1480 11330 1481 11331
rect 1489 11330 1490 11331
<< end >>
