magic
tech scmos
timestamp 1394680307
<< m1p >>
use CELL  1
transform -1 0 1046 0 1 984
box 0 0 6 6
use CELL  2
transform -1 0 1176 0 1 1140
box 0 0 6 6
use CELL  3
transform 1 0 1102 0 -1 1002
box 0 0 6 6
use CELL  4
transform -1 0 1029 0 1 1128
box 0 0 6 6
use CELL  5
transform -1 0 1074 0 1 1092
box 0 0 6 6
use CELL  6
transform -1 0 1015 0 1 1020
box 0 0 6 6
use CELL  7
transform -1 0 1045 0 1 1188
box 0 0 6 6
use CELL  8
transform 1 0 1283 0 -1 1050
box 0 0 6 6
use CELL  9
transform -1 0 1139 0 1 1140
box 0 0 6 6
use CELL  10
transform -1 0 1114 0 -1 990
box 0 0 6 6
use CELL  11
transform 1 0 1231 0 -1 1134
box 0 0 6 6
use CELL  12
transform -1 0 1230 0 1 1056
box 0 0 6 6
use CELL  13
transform 1 0 1095 0 1 984
box 0 0 6 6
use CELL  14
transform 1 0 1111 0 -1 1110
box 0 0 6 6
use CELL  15
transform -1 0 1131 0 1 1176
box 0 0 6 6
use CELL  16
transform -1 0 1088 0 1 1092
box 0 0 6 6
use CELL  17
transform 1 0 1312 0 1 1032
box 0 0 6 6
use CELL  18
transform 1 0 1189 0 -1 1002
box 0 0 6 6
use CELL  19
transform -1 0 1318 0 1 1056
box 0 0 6 6
use CELL  20
transform -1 0 1082 0 1 1032
box 0 0 6 6
use CELL  21
transform 1 0 1305 0 1 1032
box 0 0 6 6
use CELL  22
transform -1 0 1278 0 1 1032
box 0 0 6 6
use CELL  23
transform -1 0 1120 0 -1 1014
box 0 0 6 6
use CELL  24
transform 1 0 1199 0 1 1080
box 0 0 6 6
use CELL  25
transform 1 0 1219 0 1 996
box 0 0 6 6
use CELL  26
transform 1 0 1008 0 -1 1038
box 0 0 6 6
use CELL  27
transform -1 0 1217 0 1 1032
box 0 0 6 6
use CELL  28
transform 1 0 1002 0 1 1128
box 0 0 6 6
use CELL  29
transform -1 0 1065 0 1 1200
box 0 0 6 6
use CELL  30
transform -1 0 1046 0 1 1116
box 0 0 6 6
use CELL  31
transform -1 0 1021 0 1 1116
box 0 0 6 6
use CELL  32
transform 1 0 986 0 1 1044
box 0 0 6 6
use CELL  33
transform -1 0 1173 0 1 1020
box 0 0 6 6
use CELL  34
transform -1 0 1026 0 1 996
box 0 0 6 6
use CELL  35
transform 1 0 1132 0 -1 1086
box 0 0 6 6
use CELL  36
transform -1 0 1034 0 1 1140
box 0 0 6 6
use CELL  37
transform -1 0 1084 0 1 1176
box 0 0 6 6
use CELL  38
transform -1 0 1263 0 1 1116
box 0 0 6 6
use CELL  39
transform -1 0 1267 0 1 1152
box 0 0 6 6
use CELL  40
transform -1 0 1211 0 1 1128
box 0 0 6 6
use CELL  41
transform -1 0 1063 0 1 1164
box 0 0 6 6
use CELL  42
transform 1 0 1077 0 1 1020
box 0 0 6 6
use CELL  43
transform -1 0 1229 0 1 1044
box 0 0 6 6
use CELL  44
transform -1 0 1041 0 1 1044
box 0 0 6 6
use CELL  45
transform 1 0 1207 0 1 1140
box 0 0 6 6
use CELL  46
transform -1 0 1270 0 -1 1122
box 0 0 6 6
use CELL  47
transform -1 0 1295 0 1 1068
box 0 0 6 6
use CELL  48
transform -1 0 1240 0 -1 1110
box 0 0 6 6
use CELL  49
transform -1 0 1038 0 1 1176
box 0 0 6 6
use CELL  50
transform 1 0 1118 0 -1 1182
box 0 0 6 6
use CELL  51
transform 1 0 1008 0 1 996
box 0 0 6 6
use CELL  52
transform -1 0 1205 0 1 1164
box 0 0 6 6
use CELL  53
transform -1 0 1095 0 1 1152
box 0 0 6 6
use CELL  54
transform -1 0 1136 0 1 1164
box 0 0 6 6
use CELL  55
transform -1 0 1290 0 1 1152
box 0 0 6 6
use CELL  56
transform -1 0 1053 0 1 1116
box 0 0 6 6
use CELL  57
transform -1 0 1267 0 1 1068
box 0 0 6 6
use CELL  58
transform 1 0 1267 0 1 1092
box 0 0 6 6
use CELL  59
transform 1 0 1224 0 1 1128
box 0 0 6 6
use CELL  60
transform -1 0 1036 0 1 1128
box 0 0 6 6
use CELL  61
transform 1 0 1061 0 -1 1038
box 0 0 6 6
use CELL  62
transform -1 0 1269 0 1 1080
box 0 0 6 6
use CELL  63
transform 1 0 1205 0 1 996
box 0 0 6 6
use CELL  64
transform 1 0 1147 0 1 996
box 0 0 6 6
use CELL  65
transform -1 0 1023 0 1 1056
box 0 0 6 6
use CELL  66
transform 1 0 1102 0 1 1080
box 0 0 6 6
use CELL  67
transform -1 0 1030 0 1 1056
box 0 0 6 6
use CELL  68
transform -1 0 1064 0 1 1008
box 0 0 6 6
use CELL  69
transform 1 0 1212 0 1 996
box 0 0 6 6
use CELL  70
transform -1 0 1145 0 1 1104
box 0 0 6 6
use CELL  71
transform -1 0 1237 0 1 1056
box 0 0 6 6
use CELL  72
transform -1 0 1023 0 1 1080
box 0 0 6 6
use CELL  73
transform -1 0 1015 0 1 1044
box 0 0 6 6
use CELL  74
transform 1 0 1002 0 -1 1026
box 0 0 6 6
use CELL  75
transform -1 0 1105 0 1 1044
box 0 0 6 6
use CELL  76
transform -1 0 1233 0 1 1152
box 0 0 6 6
use CELL  77
transform -1 0 1044 0 1 1068
box 0 0 6 6
use CELL  78
transform -1 0 1073 0 1 984
box 0 0 6 6
use CELL  79
transform -1 0 1141 0 1 1068
box 0 0 6 6
use CELL  80
transform -1 0 1042 0 1 1104
box 0 0 6 6
use CELL  81
transform 1 0 1079 0 1 996
box 0 0 6 6
use CELL  82
transform 1 0 1319 0 1 1032
box 0 0 6 6
use CELL  83
transform -1 0 1080 0 1 1200
box 0 0 6 6
use CELL  84
transform -1 0 1266 0 1 1044
box 0 0 6 6
use CELL  85
transform -1 0 1125 0 1 1128
box 0 0 6 6
use CELL  86
transform -1 0 1085 0 1 1056
box 0 0 6 6
use CELL  87
transform -1 0 1080 0 1 984
box 0 0 6 6
use CELL  88
transform -1 0 1276 0 1 1056
box 0 0 6 6
use CELL  89
transform 1 0 1191 0 1 1092
box 0 0 6 6
use CELL  90
transform -1 0 1112 0 1 1044
box 0 0 6 6
use CELL  91
transform 1 0 1204 0 -1 1038
box 0 0 6 6
use CELL  92
transform -1 0 1255 0 1 1152
box 0 0 6 6
use CELL  93
transform -1 0 1015 0 1 1128
box 0 0 6 6
use CELL  94
transform -1 0 1108 0 1 984
box 0 0 6 6
use CELL  95
transform 1 0 1075 0 1 1092
box 0 0 6 6
use CELL  96
transform -1 0 1089 0 -1 1038
box 0 0 6 6
use CELL  97
transform -1 0 1002 0 1 1116
box 0 0 6 6
use CELL  98
transform -1 0 1199 0 1 1140
box 0 0 6 6
use CELL  99
transform 1 0 1123 0 1 1116
box 0 0 6 6
use CELL  100
transform 1 0 1219 0 1 1008
box 0 0 6 6
use CELL  101
transform -1 0 1075 0 1 1176
box 0 0 6 6
use CELL  102
transform -1 0 1323 0 1 1068
box 0 0 6 6
use CELL  103
transform -1 0 1022 0 1 1044
box 0 0 6 6
use CELL  104
transform -1 0 1047 0 1 1164
box 0 0 6 6
use CELL  105
transform 1 0 1298 0 1 1032
box 0 0 6 6
use CELL  106
transform -1 0 1058 0 1 1200
box 0 0 6 6
use CELL  107
transform -1 0 1172 0 1 1092
box 0 0 6 6
use CELL  108
transform -1 0 1057 0 1 1188
box 0 0 6 6
use CELL  109
transform 1 0 1059 0 1 1128
box 0 0 6 6
use CELL  110
transform -1 0 1154 0 1 1140
box 0 0 6 6
use CELL  111
transform -1 0 1262 0 1 1080
box 0 0 6 6
use CELL  112
transform -1 0 1253 0 1 1032
box 0 0 6 6
use CELL  113
transform -1 0 1206 0 1 1140
box 0 0 6 6
use CELL  114
transform 1 0 1235 0 1 1008
box 0 0 6 6
use CELL  115
transform 1 0 1132 0 -1 1110
box 0 0 6 6
use CELL  116
transform -1 0 1271 0 1 1032
box 0 0 6 6
use CELL  117
transform 1 0 1003 0 -1 1086
box 0 0 6 6
use CELL  118
transform 1 0 1036 0 -1 1158
box 0 0 6 6
use CELL  119
transform -1 0 1184 0 1 1104
box 0 0 6 6
use CELL  120
transform -1 0 1198 0 1 1164
box 0 0 6 6
use CELL  121
transform -1 0 1219 0 1 1080
box 0 0 6 6
use CELL  122
transform -1 0 1064 0 1 1020
box 0 0 6 6
use CELL  123
transform -1 0 1080 0 1 1008
box 0 0 6 6
use CELL  124
transform -1 0 1036 0 1 1020
box 0 0 6 6
use CELL  125
transform -1 0 1134 0 1 1068
box 0 0 6 6
use CELL  126
transform -1 0 1274 0 1 1152
box 0 0 6 6
use CELL  127
transform -1 0 1041 0 1 1092
box 0 0 6 6
use CELL  128
transform -1 0 1261 0 -1 1110
box 0 0 6 6
use CELL  129
transform -1 0 1142 0 1 1044
box 0 0 6 6
use CELL  130
transform -1 0 1228 0 1 1104
box 0 0 6 6
use CELL  131
transform -1 0 1035 0 1 1152
box 0 0 6 6
use CELL  132
transform 1 0 1038 0 -1 1206
box 0 0 6 6
use CELL  133
transform -1 0 1211 0 1 1056
box 0 0 6 6
use CELL  134
transform -1 0 1230 0 1 1020
box 0 0 6 6
use CELL  135
transform -1 0 1071 0 1 1020
box 0 0 6 6
use CELL  136
transform -1 0 1049 0 1 1152
box 0 0 6 6
use CELL  137
transform -1 0 1056 0 -1 1158
box 0 0 6 6
use CELL  138
transform -1 0 1143 0 1 1020
box 0 0 6 6
use CELL  139
transform -1 0 1040 0 1 1164
box 0 0 6 6
use CELL  140
transform 1 0 1072 0 1 1044
box 0 0 6 6
use CELL  141
transform -1 0 1110 0 1 1176
box 0 0 6 6
use CELL  142
transform -1 0 1050 0 1 1128
box 0 0 6 6
use CELL  143
transform 1 0 1112 0 -1 1194
box 0 0 6 6
use CELL  144
transform -1 0 1009 0 1 1056
box 0 0 6 6
use CELL  145
transform -1 0 1215 0 1 1092
box 0 0 6 6
use CELL  146
transform -1 0 1098 0 1 1176
box 0 0 6 6
use CELL  147
transform -1 0 1023 0 1 1068
box 0 0 6 6
use CELL  148
transform 1 0 1284 0 1 1032
box 0 0 6 6
use CELL  149
transform -1 0 1091 0 1 1176
box 0 0 6 6
use CELL  150
transform -1 0 1099 0 1 996
box 0 0 6 6
use CELL  151
transform -1 0 1154 0 1 1044
box 0 0 6 6
use CELL  152
transform 1 0 1310 0 1 1068
box 0 0 6 6
use CELL  153
transform -1 0 1009 0 1 1068
box 0 0 6 6
use CELL  154
transform 1 0 1305 0 -1 1062
box 0 0 6 6
use CELL  155
transform -1 0 1251 0 1 1128
box 0 0 6 6
use CELL  156
transform 1 0 1296 0 -1 1074
box 0 0 6 6
use CELL  157
transform 1 0 1063 0 1 996
box 0 0 6 6
use CELL  158
transform -1 0 1222 0 1 1140
box 0 0 6 6
use CELL  159
transform -1 0 1089 0 1 1188
box 0 0 6 6
use CELL  160
transform -1 0 1070 0 1 1164
box 0 0 6 6
use CELL  161
transform -1 0 1255 0 1 1020
box 0 0 6 6
use CELL  162
transform -1 0 1029 0 1 1044
box 0 0 6 6
use CELL  163
transform -1 0 1104 0 1 1068
box 0 0 6 6
use CELL  164
transform -1 0 1254 0 1 1104
box 0 0 6 6
use CELL  165
transform -1 0 1082 0 1 1164
box 0 0 6 6
use CELL  166
transform -1 0 1090 0 1 1104
box 0 0 6 6
use CELL  167
transform -1 0 1057 0 1 1008
box 0 0 6 6
use CELL  168
transform -1 0 1304 0 1 1056
box 0 0 6 6
use CELL  169
transform -1 0 1048 0 1 1044
box 0 0 6 6
use CELL  170
transform -1 0 1052 0 -1 990
box 0 0 6 6
use CELL  171
transform -1 0 1071 0 1 1008
box 0 0 6 6
use CELL  172
transform -1 0 1204 0 1 1128
box 0 0 6 6
use CELL  173
transform -1 0 1023 0 -1 1038
box 0 0 6 6
use CELL  174
transform -1 0 1111 0 -1 1194
box 0 0 6 6
use CELL  175
transform -1 0 1037 0 1 1056
box 0 0 6 6
use CELL  176
transform -1 0 1223 0 1 1128
box 0 0 6 6
use CELL  177
transform 1 0 1076 0 1 1188
box 0 0 6 6
use CELL  178
transform -1 0 1246 0 1 1068
box 0 0 6 6
use CELL  179
transform -1 0 1026 0 1 1104
box 0 0 6 6
use CELL  180
transform -1 0 1115 0 1 1164
box 0 0 6 6
use CELL  181
transform -1 0 1064 0 -1 1194
box 0 0 6 6
use CELL  182
transform 1 0 1155 0 -1 1146
box 0 0 6 6
use CELL  183
transform 1 0 1177 0 1 996
box 0 0 6 6
use CELL  184
transform -1 0 1296 0 1 1044
box 0 0 6 6
use CELL  185
transform -1 0 1044 0 1 1056
box 0 0 6 6
use CELL  186
transform -1 0 1167 0 1 1116
box 0 0 6 6
use CELL  187
transform -1 0 1071 0 1 1056
box 0 0 6 6
use CELL  188
transform -1 0 1122 0 1 1116
box 0 0 6 6
use CELL  189
transform -1 0 1062 0 1 996
box 0 0 6 6
use CELL  190
transform 1 0 1065 0 1 1068
box 0 0 6 6
use CELL  191
transform -1 0 1022 0 1 1092
box 0 0 6 6
use CELL  192
transform -1 0 1267 0 1 1092
box 0 0 6 6
use CELL  193
transform -1 0 1027 0 1 1140
box 0 0 6 6
use CELL  194
transform -1 0 985 0 1 1044
box 0 0 6 6
use CELL  195
transform -1 0 1229 0 -1 1146
box 0 0 6 6
use CELL  196
transform -1 0 1050 0 1 1092
box 0 0 6 6
use CELL  197
transform -1 0 1196 0 1 1044
box 0 0 6 6
use CELL  198
transform -1 0 1030 0 -1 1086
box 0 0 6 6
use CELL  199
transform -1 0 1288 0 1 1056
box 0 0 6 6
use CELL  200
transform -1 0 1092 0 1 996
box 0 0 6 6
use CELL  201
transform 1 0 1189 0 1 1008
box 0 0 6 6
use CELL  202
transform 1 0 1060 0 -1 990
box 0 0 6 6
use CELL  203
transform -1 0 1054 0 1 1176
box 0 0 6 6
use CELL  204
transform -1 0 1295 0 1 1056
box 0 0 6 6
use CELL  205
transform -1 0 1299 0 -1 1086
box 0 0 6 6
use CELL  206
transform 1 0 996 0 1 1056
box 0 0 6 6
use CELL  207
transform 1 0 1008 0 1 1152
box 0 0 6 6
use CELL  208
transform -1 0 1255 0 -1 1014
box 0 0 6 6
use CELL  209
transform 1 0 1300 0 1 1080
box 0 0 6 6
use CELL  210
transform -1 0 1033 0 1 1164
box 0 0 6 6
use CELL  211
transform -1 0 1043 0 1 1020
box 0 0 6 6
use CELL  212
transform -1 0 1117 0 1 1176
box 0 0 6 6
use CELL  213
transform -1 0 1002 0 1 1068
box 0 0 6 6
use CELL  214
transform -1 0 1048 0 -1 1146
box 0 0 6 6
use CELL  215
transform -1 0 1016 0 1 1080
box 0 0 6 6
use CELL  216
transform -1 0 1046 0 1 1032
box 0 0 6 6
use CELL  217
transform -1 0 1215 0 1 1116
box 0 0 6 6
use CELL  218
transform -1 0 1038 0 1 1188
box 0 0 6 6
use CELL  219
transform -1 0 1244 0 1 1128
box 0 0 6 6
use CELL  220
transform -1 0 1309 0 1 1068
box 0 0 6 6
use CELL  221
transform 1 0 1242 0 1 1008
box 0 0 6 6
use CELL  222
transform -1 0 1190 0 1 1128
box 0 0 6 6
use CELL  223
transform -1 0 1145 0 1 1080
box 0 0 6 6
use CELL  224
transform -1 0 1224 0 1 1092
box 0 0 6 6
use CELL  225
transform -1 0 1026 0 1 1164
box 0 0 6 6
use CELL  226
transform -1 0 1204 0 -1 1002
box 0 0 6 6
use CELL  227
transform -1 0 1097 0 1 1092
box 0 0 6 6
use CELL  228
transform -1 0 1276 0 1 1068
box 0 0 6 6
use CELL  229
transform -1 0 1092 0 1 1020
box 0 0 6 6
use CELL  230
transform -1 0 1014 0 1 1104
box 0 0 6 6
use CELL  231
transform -1 0 1179 0 1 1092
box 0 0 6 6
use CELL  232
transform -1 0 1220 0 1 1044
box 0 0 6 6
use CELL  233
transform -1 0 1014 0 1 1116
box 0 0 6 6
use CELL  234
transform -1 0 1125 0 1 1188
box 0 0 6 6
use CELL  235
transform -1 0 1032 0 1 984
box 0 0 6 6
use CELL  236
transform -1 0 1022 0 1 1128
box 0 0 6 6
use CELL  237
transform -1 0 1039 0 1 1008
box 0 0 6 6
use CELL  238
transform 1 0 1099 0 1 1188
box 0 0 6 6
use CELL  239
transform -1 0 1212 0 1 1080
box 0 0 6 6
use CELL  240
transform 1 0 1056 0 -1 1122
box 0 0 6 6
use CELL  241
transform -1 0 1179 0 1 1116
box 0 0 6 6
use CELL  242
transform -1 0 1197 0 1 1128
box 0 0 6 6
use CELL  243
transform -1 0 1044 0 1 1080
box 0 0 6 6
use CELL  244
transform -1 0 1015 0 1 1188
box 0 0 6 6
use CELL  245
transform -1 0 1035 0 1 1104
box 0 0 6 6
use CELL  246
transform -1 0 1140 0 1 1176
box 0 0 6 6
use CELL  247
transform -1 0 1240 0 1 1152
box 0 0 6 6
use CELL  248
transform -1 0 1231 0 1 1092
box 0 0 6 6
use CELL  249
transform -1 0 1098 0 1 1008
box 0 0 6 6
use CELL  250
transform -1 0 1160 0 1 1056
box 0 0 6 6
use CELL  251
transform -1 0 1008 0 1 1188
box 0 0 6 6
use CELL  252
transform -1 0 1029 0 1 1020
box 0 0 6 6
use CELL  253
transform 1 0 1256 0 1 1020
box 0 0 6 6
use CELL  254
transform 1 0 1022 0 -1 1158
box 0 0 6 6
use CELL  255
transform -1 0 1297 0 1 1032
box 0 0 6 6
use CELL  256
transform -1 0 1095 0 1 1128
box 0 0 6 6
use CELL  257
transform -1 0 1109 0 1 1140
box 0 0 6 6
use CELL  258
transform -1 0 1285 0 1 1080
box 0 0 6 6
use CELL  259
transform -1 0 1089 0 1 1008
box 0 0 6 6
use CELL  260
transform -1 0 1037 0 1 1080
box 0 0 6 6
use CELL  261
transform -1 0 978 0 1 1044
box 0 0 6 6
use CELL  262
transform -1 0 1030 0 1 1032
box 0 0 6 6
use CELL  263
transform -1 0 1218 0 1 1020
box 0 0 6 6
use CELL  264
transform -1 0 1259 0 1 1044
box 0 0 6 6
use CELL  265
transform -1 0 1283 0 1 1068
box 0 0 6 6
use CELL  266
transform -1 0 1192 0 1 1140
box 0 0 6 6
use CELL  267
transform -1 0 1162 0 1 1128
box 0 0 6 6
use CELL  268
transform -1 0 1028 0 -1 1122
box 0 0 6 6
use CELL  269
transform -1 0 1143 0 1 1116
box 0 0 6 6
use CELL  270
transform -1 0 1237 0 1 1116
box 0 0 6 6
use CELL  271
transform -1 0 1212 0 1 1104
box 0 0 6 6
use CELL  272
transform -1 0 1144 0 1 1008
box 0 0 6 6
use CELL  273
transform 1 0 1213 0 1 1104
box 0 0 6 6
use CELL  274
transform -1 0 1282 0 1 1044
box 0 0 6 6
use CELL  275
transform -1 0 1127 0 1 1164
box 0 0 6 6
use CELL  276
transform 1 0 1173 0 1 1152
box 0 0 6 6
use CELL  277
transform -1 0 1248 0 1 1020
box 0 0 6 6
use CELL  278
transform -1 0 1088 0 1 1152
box 0 0 6 6
use CELL  279
transform 1 0 1164 0 -1 1182
box 0 0 6 6
use CELL  280
transform -1 0 1064 0 1 1140
box 0 0 6 6
use CELL  281
transform -1 0 1231 0 1 1080
box 0 0 6 6
use CELL  282
transform -1 0 1030 0 1 1068
box 0 0 6 6
use CELL  283
transform -1 0 1045 0 1 1176
box 0 0 6 6
use CELL  284
transform -1 0 1087 0 1 984
box 0 0 6 6
use CELL  285
transform -1 0 1258 0 -1 1134
box 0 0 6 6
use CELL  286
transform 1 0 1177 0 1 1140
box 0 0 6 6
use CELL  287
transform -1 0 1098 0 -1 1194
box 0 0 6 6
use CELL  288
transform -1 0 1205 0 1 1044
box 0 0 6 6
use CELL  289
transform 1 0 1185 0 -1 1170
box 0 0 6 6
use CELL  290
transform -1 0 1099 0 -1 1110
box 0 0 6 6
use CELL  291
transform -1 0 1184 0 -1 1170
box 0 0 6 6
use CELL  292
transform 1 0 1205 0 1 1164
box 0 0 6 6
use CELL  293
transform -1 0 1101 0 1 1080
box 0 0 6 6
use CELL  294
transform -1 0 1203 0 1 1032
box 0 0 6 6
use CELL  295
transform -1 0 1154 0 -1 1098
box 0 0 6 6
use CELL  296
transform -1 0 1136 0 1 1056
box 0 0 6 6
use CELL  297
transform -1 0 1269 0 1 1020
box 0 0 6 6
use CELL  298
transform -1 0 1032 0 1 1008
box 0 0 6 6
use CELL  299
transform -1 0 1246 0 1 1092
box 0 0 6 6
use CELL  300
transform 1 0 1053 0 -1 990
box 0 0 6 6
use CELL  301
transform -1 0 1094 0 1 1200
box 0 0 6 6
use CELL  302
transform -1 0 1264 0 1 1056
box 0 0 6 6
use CELL  303
transform 1 0 1010 0 1 1068
box 0 0 6 6
use CELL  304
transform 1 0 1037 0 -1 1134
box 0 0 6 6
use CELL  305
transform -1 0 1222 0 -1 1122
box 0 0 6 6
use CELL  306
transform -1 0 1292 0 1 1080
box 0 0 6 6
use CELL  307
transform -1 0 1244 0 -1 1122
box 0 0 6 6
use CELL  308
transform -1 0 1255 0 1 1068
box 0 0 6 6
use CELL  309
transform -1 0 1054 0 1 1164
box 0 0 6 6
use CELL  310
transform 1 0 1068 0 1 1152
box 0 0 6 6
use CELL  311
transform 1 0 1126 0 1 1188
box 0 0 6 6
use CELL  312
transform -1 0 1278 0 1 1080
box 0 0 6 6
use CELL  313
transform -1 0 1051 0 1 1200
box 0 0 6 6
use CELL  314
transform -1 0 1037 0 1 1068
box 0 0 6 6
use CELL  315
transform -1 0 1283 0 1 1020
box 0 0 6 6
use CELL  316
transform -1 0 1105 0 1 1008
box 0 0 6 6
use CELL  317
transform -1 0 1038 0 1 996
box 0 0 6 6
use CELL  318
transform -1 0 1136 0 1 1116
box 0 0 6 6
use CELL  319
transform -1 0 1169 0 1 1128
box 0 0 6 6
use CELL  320
transform -1 0 1002 0 1 1080
box 0 0 6 6
use CELL  321
transform 1 0 1325 0 1 1032
box 0 0 6 6
use CELL  322
transform -1 0 1008 0 1 1092
box 0 0 6 6
use CELL  323
transform -1 0 1057 0 1 1140
box 0 0 6 6
use CELL  324
transform -1 0 1256 0 1 1116
box 0 0 6 6
use CELL  325
transform 1 0 1269 0 -1 1050
box 0 0 6 6
use CELL  326
transform -1 0 1021 0 1 1152
box 0 0 6 6
use CELL  327
transform -1 0 1087 0 1 1200
box 0 0 6 6
use CELL  328
transform -1 0 1002 0 1 1104
box 0 0 6 6
use CELL  329
transform -1 0 1218 0 1 1056
box 0 0 6 6
use CELL  330
transform -1 0 1020 0 1 1140
box 0 0 6 6
use CELL  331
transform -1 0 1081 0 1 1152
box 0 0 6 6
use CELL  332
transform -1 0 1075 0 1 1104
box 0 0 6 6
use CELL  333
transform -1 0 1094 0 1 984
box 0 0 6 6
use CELL  334
transform -1 0 1029 0 1 1092
box 0 0 6 6
use CELL  335
transform 1 0 1070 0 1 996
box 0 0 6 6
use CELL  336
transform -1 0 1132 0 1 1128
box 0 0 6 6
use CELL  337
transform -1 0 1016 0 1 1056
box 0 0 6 6
use CELL  338
transform 1 0 1016 0 1 1020
box 0 0 6 6
use CELL  339
transform -1 0 1039 0 1 984
box 0 0 6 6
use CELL  340
transform -1 0 1283 0 1 1152
box 0 0 6 6
use CELL  341
transform -1 0 1221 0 1 1152
box 0 0 6 6
use CELL  342
transform -1 0 1148 0 1 1164
box 0 0 6 6
use CELL  343
transform -1 0 1255 0 1 1080
box 0 0 6 6
use CELL  344
transform 1 0 1185 0 1 1104
box 0 0 6 6
use CELL  345
transform -1 0 1234 0 1 1068
box 0 0 6 6
use CELL  346
transform -1 0 1008 0 1 1044
box 0 0 6 6
use CELL  347
transform -1 0 1260 0 1 1092
box 0 0 6 6
use CELL  348
transform -1 0 1128 0 1 1020
box 0 0 6 6
use CELL  349
transform -1 0 1015 0 1 1092
box 0 0 6 6
use CELL  350
transform -1 0 1041 0 1 1140
box 0 0 6 6
use CELL  351
transform 1 0 1233 0 1 1020
box 0 0 6 6
use CELL  352
transform -1 0 1120 0 -1 1002
box 0 0 6 6
use CELL  353
transform -1 0 1094 0 1 1164
box 0 0 6 6
use CELL  354
transform -1 0 1078 0 1 1056
box 0 0 6 6
use CELL  355
transform 1 0 1228 0 1 1008
box 0 0 6 6
use CELL  356
transform -1 0 1247 0 1 1104
box 0 0 6 6
use CELL  357
transform -1 0 1185 0 -1 1026
box 0 0 6 6
use CELL  358
transform -1 0 1276 0 1 1020
box 0 0 6 6
use CELL  359
transform -1 0 1037 0 1 1032
box 0 0 6 6
use CELL  360
transform 1 0 1247 0 -1 1098
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 1050 0 1 996
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 1045 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 1049 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 1055 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 1127 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 1151 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 1125 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 1080 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 1056 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 1066 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 1053 0 1 996
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 1048 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 1052 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 1058 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 1060 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 1050 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 1044 0 1 996
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 1221 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 1037 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 1026 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 1065 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 1034 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 1063 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 1095 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 1050 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 1077 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 1056 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 1056 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 1066 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 1008 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 1014 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 1090 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 1295 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 1161 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 1103 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 1144 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 1141 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 1149 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 1129 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 1106 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 1195 0 1 996
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 1225 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 1239 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 1205 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 1235 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 1173 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 1153 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 1138 0 1 996
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 1171 0 1 996
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 1162 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 1103 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 1175 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 1172 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 1243 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 1126 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 1175 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 1126 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 1195 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 1109 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 1210 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 1296 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 1119 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 1080 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 1076 0 1 996
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 1187 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 1196 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 1209 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 1177 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 1168 0 1 996
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 1225 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 1160 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 1054 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 1051 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 1048 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 1041 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 1044 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 1077 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 1062 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 1217 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 1208 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 1144 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 1141 0 1 996
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 1071 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 1055 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 1104 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 1054 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 1062 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 1086 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 1106 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 1170 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 1130 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 1138 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 1137 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 1109 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 1075 0 1 1176
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 1070 0 1 1188
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 1243 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 1267 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 1237 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 1200 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 1197 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 1225 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 1085 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 1110 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 1276 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 1266 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 1278 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 1230 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-109
transform 1 0 1207 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-110
transform 1 0 1183 0 1 996
box 0 0 3 6
use FEEDTHRU  F-111
transform 1 0 1237 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-112
transform 1 0 1269 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-113
transform 1 0 1045 0 1 1188
box 0 0 3 6
use FEEDTHRU  F-114
transform 1 0 1160 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-115
transform 1 0 1240 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-116
transform 1 0 1183 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-117
transform 1 0 1246 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-118
transform 1 0 1240 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-119
transform 1 0 1261 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-120
transform 1 0 1213 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-121
transform 1 0 1274 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-122
transform 1 0 1110 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-123
transform 1 0 1097 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-124
transform 1 0 1095 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-125
transform 1 0 1231 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-126
transform 1 0 1228 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-127
transform 1 0 1244 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-128
transform 1 0 1211 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-129
transform 1 0 1283 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-130
transform 1 0 1074 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-131
transform 1 0 1096 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-132
transform 1 0 1222 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-133
transform 1 0 1193 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-134
transform 1 0 1175 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-135
transform 1 0 1194 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-136
transform 1 0 1116 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-137
transform 1 0 1191 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-138
transform 1 0 1184 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-139
transform 1 0 1197 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-140
transform 1 0 1234 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-141
transform 1 0 1255 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-142
transform 1 0 1247 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-143
transform 1 0 1259 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-144
transform 1 0 1206 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-145
transform 1 0 1174 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-146
transform 1 0 1165 0 1 996
box 0 0 3 6
use FEEDTHRU  F-147
transform 1 0 1250 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-148
transform 1 0 1262 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-149
transform 1 0 1194 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-150
transform 1 0 1037 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-151
transform 1 0 1078 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-152
transform 1 0 1155 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-153
transform 1 0 1092 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-154
transform 1 0 1187 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-155
transform 1 0 1219 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-156
transform 1 0 1193 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-157
transform 1 0 1136 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-158
transform 1 0 1166 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-159
transform 1 0 1186 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-160
transform 1 0 1196 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-161
transform 1 0 1139 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-162
transform 1 0 1163 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-163
transform 1 0 1136 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-164
transform 1 0 1130 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-165
transform 1 0 1067 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-166
transform 1 0 1126 0 1 996
box 0 0 3 6
use FEEDTHRU  F-167
transform 1 0 1184 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-168
transform 1 0 1181 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-169
transform 1 0 1164 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-170
transform 1 0 1089 0 1 1188
box 0 0 3 6
use FEEDTHRU  F-171
transform 1 0 1098 0 1 1176
box 0 0 3 6
use FEEDTHRU  F-172
transform 1 0 1281 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-173
transform 1 0 1279 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-174
transform 1 0 1192 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-175
transform 1 0 1163 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-176
transform 1 0 1140 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-177
transform 1 0 1107 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-178
transform 1 0 1166 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-179
transform 1 0 1143 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-180
transform 1 0 1110 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-181
transform 1 0 1105 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-182
transform 1 0 1099 0 1 996
box 0 0 3 6
use FEEDTHRU  F-183
transform 1 0 1144 0 1 996
box 0 0 3 6
use FEEDTHRU  F-184
transform 1 0 1053 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-185
transform 1 0 1060 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-186
transform 1 0 1059 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-187
transform 1 0 1089 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-188
transform 1 0 1080 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-189
transform 1 0 1088 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-190
transform 1 0 1087 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-191
transform 1 0 1186 0 1 996
box 0 0 3 6
use FEEDTHRU  F-192
transform 1 0 1180 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-193
transform 1 0 1255 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-194
transform 1 0 1166 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-195
transform 1 0 1123 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-196
transform 1 0 1115 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-197
transform 1 0 1172 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-198
transform 1 0 1174 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-199
transform 1 0 1117 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-200
transform 1 0 1118 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-201
transform 1 0 1163 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-202
transform 1 0 1162 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-203
transform 1 0 1264 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-204
transform 1 0 1241 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-205
transform 1 0 1241 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-206
transform 1 0 1218 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-207
transform 1 0 1213 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-208
transform 1 0 1046 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-209
transform 1 0 1125 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-210
transform 1 0 1073 0 1 1188
box 0 0 3 6
use FEEDTHRU  F-211
transform 1 0 1060 0 1 1176
box 0 0 3 6
use FEEDTHRU  F-212
transform 1 0 1063 0 1 1176
box 0 0 3 6
use FEEDTHRU  F-213
transform 1 0 1121 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-214
transform 1 0 1131 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-215
transform 1 0 1203 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-216
transform 1 0 1206 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-217
transform 1 0 1127 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-218
transform 1 0 1234 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-219
transform 1 0 1179 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-220
transform 1 0 1176 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-221
transform 1 0 1150 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-222
transform 1 0 1149 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-223
transform 1 0 1070 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-224
transform 1 0 1203 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-225
transform 1 0 1206 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-226
transform 1 0 1169 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-227
transform 1 0 1164 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-228
transform 1 0 1197 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-229
transform 1 0 1207 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-230
transform 1 0 1210 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-231
transform 1 0 1199 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-232
transform 1 0 1114 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-233
transform 1 0 1107 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-234
transform 1 0 1215 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-235
transform 1 0 1246 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-236
transform 1 0 1246 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-237
transform 1 0 1267 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-238
transform 1 0 1244 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-239
transform 1 0 1244 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-240
transform 1 0 1221 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-241
transform 1 0 1216 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-242
transform 1 0 1174 0 1 996
box 0 0 3 6
use FEEDTHRU  F-243
transform 1 0 1167 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-244
transform 1 0 1089 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-245
transform 1 0 1104 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-246
transform 1 0 1100 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-247
transform 1 0 1083 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-248
transform 1 0 1113 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-249
transform 1 0 1064 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-250
transform 1 0 1068 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-251
transform 1 0 1068 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-252
transform 1 0 1102 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-253
transform 1 0 1048 0 1 1188
box 0 0 3 6
use FEEDTHRU  F-254
transform 1 0 1045 0 1 1176
box 0 0 3 6
use FEEDTHRU  F-255
transform 1 0 1073 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-256
transform 1 0 1170 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-257
transform 1 0 1148 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-258
transform 1 0 1122 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-259
transform 1 0 1118 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-260
transform 1 0 1200 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-261
transform 1 0 1167 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-262
transform 1 0 1172 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-263
transform 1 0 1092 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-264
transform 1 0 1082 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-265
transform 1 0 1128 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-266
transform 1 0 1101 0 1 1176
box 0 0 3 6
use FEEDTHRU  F-267
transform 1 0 1169 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-268
transform 1 0 1258 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-269
transform 1 0 1161 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-270
transform 1 0 1214 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-271
transform 1 0 1247 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-272
transform 1 0 1231 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-273
transform 1 0 1234 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-274
transform 1 0 1219 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-275
transform 1 0 1286 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-276
transform 1 0 1218 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-277
transform 1 0 1071 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-278
transform 1 0 1068 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-279
transform 1 0 1200 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-280
transform 1 0 1228 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-281
transform 1 0 1100 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-282
transform 1 0 1158 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-283
transform 1 0 1126 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-284
transform 1 0 1101 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-285
transform 1 0 1071 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-286
transform 1 0 1053 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-287
transform 1 0 1056 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-288
transform 1 0 1222 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-289
transform 1 0 1219 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-290
transform 1 0 1206 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-291
transform 1 0 1231 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-292
transform 1 0 1066 0 1 1176
box 0 0 3 6
use FEEDTHRU  F-293
transform 1 0 1094 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-294
transform 1 0 1121 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-295
transform 1 0 1142 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-296
transform 1 0 1142 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-297
transform 1 0 1070 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-298
transform 1 0 1108 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-299
transform 1 0 1097 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-300
transform 1 0 1140 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-301
transform 1 0 1104 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-302
transform 1 0 1107 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-303
transform 1 0 1124 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-304
transform 1 0 1134 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-305
transform 1 0 1107 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-306
transform 1 0 1110 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-307
transform 1 0 1085 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-308
transform 1 0 1220 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-309
transform 1 0 1188 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-310
transform 1 0 1185 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-311
transform 1 0 1186 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-312
transform 1 0 1139 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-313
transform 1 0 1104 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-314
transform 1 0 1092 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-315
transform 1 0 1158 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-316
transform 1 0 1175 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-317
transform 1 0 1093 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-318
transform 1 0 1092 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-319
transform 1 0 1117 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-320
transform 1 0 1062 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-321
transform 1 0 1074 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-322
transform 1 0 1083 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-323
transform 1 0 1106 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-324
transform 1 0 1152 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-325
transform 1 0 1115 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-326
transform 1 0 1165 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-327
transform 1 0 1155 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-328
transform 1 0 1173 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-329
transform 1 0 1182 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-330
transform 1 0 1124 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-331
transform 1 0 1095 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-332
transform 1 0 1181 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-333
transform 1 0 1191 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-334
transform 1 0 1081 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-335
transform 1 0 1077 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-336
transform 1 0 1080 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-337
transform 1 0 1107 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-338
transform 1 0 1113 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-339
transform 1 0 1129 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-340
transform 1 0 1196 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-341
transform 1 0 1152 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-342
transform 1 0 1158 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-343
transform 1 0 1198 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-344
transform 1 0 1062 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-345
transform 1 0 1053 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-346
transform 1 0 1050 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-347
transform 1 0 1048 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-348
transform 1 0 1101 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-349
transform 1 0 1070 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-350
transform 1 0 1074 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-351
transform 1 0 1115 0 1 1164
box 0 0 3 6
use FEEDTHRU  F-352
transform 1 0 1224 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-353
transform 1 0 1127 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-354
transform 1 0 1133 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-355
transform 1 0 1112 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-356
transform 1 0 1083 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-357
transform 1 0 1089 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-358
transform 1 0 1194 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-359
transform 1 0 1203 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-360
transform 1 0 1190 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-361
transform 1 0 1113 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-362
transform 1 0 1169 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-363
transform 1 0 1237 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-364
transform 1 0 1249 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-365
transform 1 0 1153 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-366
transform 1 0 1243 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-367
transform 1 0 1133 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-368
transform 1 0 1151 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-369
transform 1 0 1238 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-370
transform 1 0 1128 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-371
transform 1 0 1258 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-372
transform 1 0 1163 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-373
transform 1 0 1160 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-374
transform 1 0 1104 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-375
transform 1 0 1157 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-376
transform 1 0 1145 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-377
transform 1 0 1160 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-378
transform 1 0 1152 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-379
transform 1 0 1222 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-380
transform 1 0 1180 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-381
transform 1 0 1088 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-382
transform 1 0 1099 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-383
transform 1 0 1086 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-384
transform 1 0 1113 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-385
transform 1 0 1112 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-386
transform 1 0 1146 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-387
transform 1 0 1147 0 1 1128
box 0 0 3 6
use FEEDTHRU  F-388
transform 1 0 1139 0 1 1140
box 0 0 3 6
use FEEDTHRU  F-389
transform 1 0 1246 0 1 1152
box 0 0 3 6
use FEEDTHRU  F-390
transform 1 0 1172 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-391
transform 1 0 1182 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-392
transform 1 0 1203 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-393
transform 1 0 1143 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-394
transform 1 0 1134 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-395
transform 1 0 1161 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-396
transform 1 0 1118 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-397
transform 1 0 1135 0 1 996
box 0 0 3 6
use FEEDTHRU  F-398
transform 1 0 1131 0 1 1176
box 0 0 3 6
use FEEDTHRU  F-399
transform 1 0 1132 0 1 1188
box 0 0 3 6
use FEEDTHRU  F-400
transform 1 0 1143 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-401
transform 1 0 1154 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-402
transform 1 0 1142 0 1 1092
box 0 0 3 6
use FEEDTHRU  F-403
transform 1 0 1157 0 1 1080
box 0 0 3 6
use FEEDTHRU  F-404
transform 1 0 1156 0 1 1068
box 0 0 3 6
use FEEDTHRU  F-405
transform 1 0 1202 0 1 1056
box 0 0 3 6
use FEEDTHRU  F-406
transform 1 0 1211 0 1 1044
box 0 0 3 6
use FEEDTHRU  F-407
transform 1 0 1220 0 1 1032
box 0 0 3 6
use FEEDTHRU  F-408
transform 1 0 1134 0 1 1020
box 0 0 3 6
use FEEDTHRU  F-409
transform 1 0 1147 0 1 1008
box 0 0 3 6
use FEEDTHRU  F-410
transform 1 0 1129 0 1 996
box 0 0 3 6
use FEEDTHRU  F-411
transform 1 0 1090 0 1 1104
box 0 0 3 6
use FEEDTHRU  F-412
transform 1 0 1074 0 1 1116
box 0 0 3 6
use FEEDTHRU  F-413
transform 1 0 1065 0 1 1128
box 0 0 3 6
<< end >>
