magic
tech scmos
timestamp 1395743070
<< m1p >>
use CELL  1
transform 1 0 352 0 1 188
box 0 0 6 6
use CELL  2
transform -1 0 356 0 1 355
box 0 0 6 6
use CELL  3
transform -1 0 265 0 -1 482
box 0 0 6 6
use CELL  4
transform -1 0 253 0 1 188
box 0 0 6 6
use CELL  5
transform -1 0 379 0 1 245
box 0 0 6 6
use CELL  6
transform 1 0 314 0 -1 410
box 0 0 6 6
use CELL  7
transform -1 0 258 0 1 149
box 0 0 6 6
use CELL  8
transform -1 0 339 0 1 298
box 0 0 6 6
use CELL  9
transform 1 0 357 0 1 355
box 0 0 6 6
use CELL  10
transform 1 0 312 0 -1 155
box 0 0 6 6
use CELL  11
transform -1 0 375 0 1 404
box 0 0 6 6
use CELL  12
transform -1 0 229 0 1 298
box 0 0 6 6
use CELL  13
transform -1 0 261 0 -1 130
box 0 0 6 6
use CELL  14
transform -1 0 242 0 1 355
box 0 0 6 6
use CELL  15
transform 1 0 352 0 -1 304
box 0 0 6 6
use CELL  16
transform -1 0 240 0 1 404
box 0 0 6 6
use CELL  17
transform -1 0 309 0 1 476
box 0 0 6 6
use CELL  18
transform 1 0 271 0 1 476
box 0 0 6 6
use CELL  19
transform 1 0 292 0 1 455
box 0 0 6 6
use CELL  20
transform 1 0 285 0 -1 482
box 0 0 6 6
use CELL  21
transform 1 0 364 0 -1 361
box 0 0 6 6
use CELL  22
transform -1 0 258 0 -1 482
box 0 0 6 6
use CELL  23
transform 1 0 245 0 -1 361
box 0 0 6 6
use CELL  24
transform -1 0 368 0 1 404
box 0 0 6 6
use CELL  25
transform -1 0 247 0 1 455
box 0 0 6 6
use CELL  26
transform -1 0 295 0 1 124
box 0 0 6 6
use CELL  27
transform -1 0 337 0 1 455
box 0 0 6 6
use CELL  28
transform -1 0 261 0 1 455
box 0 0 6 6
use CELL  29
transform -1 0 258 0 1 404
box 0 0 6 6
use CELL  30
transform -1 0 228 0 1 355
box 0 0 6 6
use CELL  31
transform -1 0 272 0 1 404
box 0 0 6 6
use CELL  32
transform 1 0 294 0 1 298
box 0 0 6 6
use CELL  33
transform -1 0 243 0 1 245
box 0 0 6 6
use CELL  34
transform -1 0 234 0 1 149
box 0 0 6 6
use CELL  35
transform 1 0 303 0 -1 155
box 0 0 6 6
use CELL  36
transform -1 0 322 0 1 188
box 0 0 6 6
use CELL  37
transform -1 0 325 0 1 355
box 0 0 6 6
use CELL  38
transform -1 0 236 0 1 298
box 0 0 6 6
use CELL  39
transform -1 0 246 0 1 188
box 0 0 6 6
use CELL  40
transform -1 0 310 0 1 188
box 0 0 6 6
use CELL  41
transform 1 0 216 0 -1 304
box 0 0 6 6
use CELL  42
transform -1 0 291 0 1 298
box 0 0 6 6
use CELL  43
transform -1 0 397 0 1 404
box 0 0 6 6
use CELL  44
transform -1 0 252 0 1 124
box 0 0 6 6
use CELL  45
transform -1 0 374 0 1 188
box 0 0 6 6
use CELL  46
transform -1 0 243 0 1 298
box 0 0 6 6
use CELL  47
transform 1 0 229 0 1 355
box 0 0 6 6
use CELL  48
transform -1 0 274 0 1 355
box 0 0 6 6
use CELL  49
transform 1 0 278 0 -1 482
box 0 0 6 6
use CELL  50
transform -1 0 404 0 1 404
box 0 0 6 6
use CELL  51
transform -1 0 288 0 -1 499
box 0 0 6 6
use CELL  52
transform -1 0 332 0 1 355
box 0 0 6 6
use CELL  53
transform -1 0 286 0 1 245
box 0 0 6 6
use CELL  54
transform -1 0 250 0 1 245
box 0 0 6 6
use CELL  55
transform 1 0 361 0 1 188
box 0 0 6 6
use CELL  56
transform -1 0 301 0 1 124
box 0 0 6 6
use CELL  57
transform 1 0 307 0 1 355
box 0 0 6 6
use CELL  58
transform -1 0 337 0 1 245
box 0 0 6 6
use CELL  59
transform -1 0 268 0 1 455
box 0 0 6 6
use CELL  60
transform -1 0 330 0 1 455
box 0 0 6 6
use CELL  61
transform -1 0 279 0 1 493
box 0 0 6 6
use CELL  62
transform -1 0 365 0 1 298
box 0 0 6 6
use CELL  63
transform 1 0 299 0 1 455
box 0 0 6 6
use CELL  64
transform -1 0 264 0 -1 112
box 0 0 6 6
use CELL  65
transform -1 0 268 0 1 124
box 0 0 6 6
use CELL  66
transform -1 0 346 0 1 298
box 0 0 6 6
use CELL  67
transform 1 0 248 0 1 455
box 0 0 6 6
use CELL  68
transform -1 0 390 0 1 404
box 0 0 6 6
use CELL  69
transform -1 0 267 0 1 355
box 0 0 6 6
use CELL  70
transform 1 0 303 0 -1 304
box 0 0 6 6
use CELL  71
transform -1 0 379 0 1 298
box 0 0 6 6
use CELL  72
transform 1 0 310 0 1 245
box 0 0 6 6
use CELL  73
transform -1 0 386 0 1 245
box 0 0 6 6
use CELL  74
transform 1 0 223 0 1 245
box 0 0 6 6
use CELL  75
transform -1 0 372 0 1 298
box 0 0 6 6
use CELL  76
transform -1 0 323 0 1 455
box 0 0 6 6
use CELL  77
transform -1 0 236 0 1 245
box 0 0 6 6
use CELL  78
transform -1 0 286 0 1 188
box 0 0 6 6
use CELL  79
transform -1 0 240 0 1 455
box 0 0 6 6
use CELL  80
transform -1 0 222 0 1 245
box 0 0 6 6
use CELL  81
transform 1 0 273 0 -1 304
box 0 0 6 6
use CELL  82
transform -1 0 273 0 1 149
box 0 0 6 6
use CELL  83
transform -1 0 302 0 1 404
box 0 0 6 6
use CELL  84
transform -1 0 300 0 1 149
box 0 0 6 6
use CELL  85
transform -1 0 258 0 1 355
box 0 0 6 6
use CELL  86
transform -1 0 393 0 1 245
box 0 0 6 6
use CELL  87
transform -1 0 265 0 1 404
box 0 0 6 6
use CELL  88
transform -1 0 381 0 -1 194
box 0 0 6 6
use CELL  89
transform -1 0 349 0 1 245
box 0 0 6 6
use CELL  90
transform -1 0 277 0 1 245
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 344 0 1 355
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 381 0 1 404
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 347 0 1 355
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 268 0 1 476
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 289 0 1 455
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 313 0 1 188
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 274 0 1 188
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 367 0 1 245
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 346 0 1 298
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 370 0 1 245
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 355 0 1 245
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 282 0 1 149
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 331 0 1 188
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 301 0 1 245
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 324 0 1 298
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 301 0 1 355
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 311 0 1 404
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 335 0 1 355
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 375 0 1 404
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 309 0 1 149
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 358 0 1 188
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 349 0 1 245
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 356 0 1 404
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 313 0 1 355
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 359 0 1 404
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 338 0 1 404
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 270 0 1 298
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 249 0 1 404
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 242 0 1 355
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 255 0 1 298
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 268 0 1 245
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 246 0 1 404
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 279 0 1 493
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 297 0 1 476
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 300 0 1 476
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 332 0 1 355
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 277 0 1 455
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 305 0 1 404
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 265 0 1 476
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 283 0 1 124
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 274 0 1 455
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 281 0 1 404
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 272 0 1 404
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 243 0 1 298
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 290 0 1 404
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 267 0 1 298
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 271 0 1 188
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 237 0 1 149
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 268 0 1 188
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 234 0 1 149
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 265 0 1 188
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 265 0 1 245
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 300 0 1 149
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 349 0 1 188
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 346 0 1 188
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 291 0 1 149
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 286 0 1 124
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 322 0 1 245
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 327 0 1 298
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 304 0 1 355
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 288 0 1 149
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 271 0 1 124
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 298 0 1 355
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 315 0 1 298
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 282 0 1 298
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 256 0 1 245
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 262 0 1 245
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 295 0 1 188
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 277 0 1 245
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 292 0 1 188
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 340 0 1 188
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 343 0 1 188
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 307 0 1 245
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 252 0 1 298
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 291 0 1 298
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 286 0 1 245
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 258 0 1 355
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 287 0 1 404
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 378 0 1 404
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 252 0 1 124
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 264 0 1 149
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 310 0 1 188
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 337 0 1 245
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 280 0 1 355
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 283 0 1 355
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 270 0 1 493
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 332 0 1 404
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 300 0 1 298
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 304 0 1 245
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 286 0 1 455
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 308 0 1 404
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 330 0 1 298
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 340 0 1 245
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 268 0 1 124
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 285 0 1 149
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 302 0 1 404
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 311 0 1 455
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 326 0 1 404
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 316 0 1 355
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 349 0 1 298
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 316 0 1 245
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 314 0 1 455
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 320 0 1 404
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 279 0 1 298
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 328 0 1 188
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 279 0 1 149
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 322 0 1 188
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 289 0 1 245
box 0 0 3 6
<< metal1 >>
rect 247 113 254 114
rect 250 115 288 116
rect 262 117 270 118
rect 266 119 285 120
rect 272 121 297 122
rect 229 131 236 132
rect 232 133 239 134
rect 247 133 260 134
rect 250 135 296 136
rect 266 137 270 138
rect 253 139 266 140
rect 284 139 294 140
rect 253 141 284 142
rect 287 141 293 142
rect 263 143 287 144
rect 290 143 299 144
rect 272 145 290 146
rect 271 147 281 148
rect 301 147 305 148
rect 310 147 314 148
rect 238 156 273 157
rect 251 158 276 159
rect 253 160 315 161
rect 256 162 299 163
rect 268 164 287 165
rect 229 166 270 167
rect 280 166 330 167
rect 283 168 333 169
rect 284 170 324 171
rect 289 172 321 173
rect 292 174 348 175
rect 241 176 294 177
rect 295 176 342 177
rect 244 178 297 179
rect 301 178 351 179
rect 308 180 345 181
rect 310 182 360 183
rect 265 184 312 185
rect 235 186 267 187
rect 372 186 377 187
rect 220 195 258 196
rect 234 197 270 198
rect 231 199 270 200
rect 241 201 273 202
rect 245 203 264 204
rect 248 205 294 206
rect 251 207 315 208
rect 272 209 288 210
rect 278 211 297 212
rect 281 213 306 214
rect 284 215 330 216
rect 275 217 285 218
rect 290 217 324 218
rect 302 219 333 220
rect 308 221 342 222
rect 308 223 345 224
rect 317 225 324 226
rect 317 227 345 228
rect 320 229 348 230
rect 332 231 351 232
rect 338 233 370 234
rect 341 235 382 236
rect 350 237 360 238
rect 356 239 375 240
rect 368 241 389 242
rect 371 243 378 244
rect 217 252 245 253
rect 220 254 254 255
rect 231 256 264 257
rect 248 258 306 259
rect 266 260 285 261
rect 257 262 284 263
rect 256 264 270 265
rect 241 266 269 267
rect 272 266 279 267
rect 241 268 272 269
rect 275 268 291 269
rect 287 270 293 271
rect 302 270 336 271
rect 281 272 302 273
rect 234 274 281 275
rect 227 276 235 277
rect 308 276 389 277
rect 323 278 329 279
rect 331 278 364 279
rect 338 280 382 281
rect 325 282 338 283
rect 341 282 361 283
rect 344 284 372 285
rect 347 286 357 287
rect 347 288 375 289
rect 350 290 354 291
rect 317 292 351 293
rect 304 294 317 295
rect 368 294 378 295
rect 370 296 378 297
rect 220 305 254 306
rect 224 307 227 308
rect 223 309 245 310
rect 231 311 284 312
rect 234 313 242 314
rect 238 315 269 316
rect 240 317 272 318
rect 243 319 257 320
rect 256 321 302 322
rect 259 323 287 324
rect 262 325 285 326
rect 272 327 300 328
rect 277 329 281 330
rect 269 331 282 332
rect 289 331 293 332
rect 302 331 326 332
rect 305 333 329 334
rect 314 335 324 336
rect 316 337 321 338
rect 317 339 351 340
rect 331 341 368 342
rect 334 343 342 344
rect 333 345 369 346
rect 345 347 355 348
rect 347 349 361 350
rect 336 351 362 352
rect 348 353 352 354
rect 230 362 238 363
rect 238 364 244 365
rect 246 364 251 365
rect 235 366 248 367
rect 256 366 292 367
rect 259 368 289 369
rect 269 370 285 371
rect 272 372 282 373
rect 260 374 274 375
rect 267 376 283 377
rect 299 376 321 377
rect 265 378 301 379
rect 297 380 322 381
rect 302 382 313 383
rect 262 384 304 385
rect 263 386 310 387
rect 305 388 389 389
rect 270 390 307 391
rect 314 390 358 391
rect 327 392 349 393
rect 317 394 328 395
rect 333 394 396 395
rect 330 396 334 397
rect 336 396 377 397
rect 339 398 374 399
rect 345 400 383 401
rect 360 402 367 403
rect 379 402 386 403
rect 235 411 251 412
rect 235 413 248 414
rect 242 415 257 416
rect 253 417 274 418
rect 260 419 289 420
rect 263 421 304 422
rect 263 423 326 424
rect 267 425 292 426
rect 256 427 291 428
rect 275 429 283 430
rect 278 431 307 432
rect 287 433 310 434
rect 312 433 319 434
rect 312 435 328 436
rect 315 437 367 438
rect 315 439 322 440
rect 321 441 334 442
rect 332 443 400 444
rect 339 445 386 446
rect 357 447 374 448
rect 360 449 371 450
rect 376 449 396 450
rect 379 451 393 452
rect 382 453 389 454
rect 238 462 243 463
rect 256 462 276 463
rect 256 464 279 465
rect 259 466 264 467
rect 266 466 288 467
rect 253 468 267 469
rect 269 468 291 469
rect 282 470 304 471
rect 286 472 299 473
rect 301 472 308 473
rect 312 472 322 473
rect 315 474 319 475
rect 328 474 336 475
rect 256 483 267 484
rect 260 485 270 486
rect 271 485 280 486
rect 274 487 302 488
rect 280 489 308 490
rect 298 491 305 492
rect 271 500 275 501
rect 280 500 284 501
<< metal2 >>
rect 247 113 248 125
rect 253 113 254 125
rect 250 115 251 125
rect 287 115 288 125
rect 262 111 263 118
rect 269 117 270 125
rect 266 119 267 125
rect 284 119 285 125
rect 272 121 273 125
rect 296 121 297 125
rect 229 131 230 150
rect 235 131 236 150
rect 232 133 233 150
rect 238 133 239 150
rect 247 129 248 134
rect 259 129 260 134
rect 250 129 251 136
rect 295 135 296 150
rect 266 129 267 138
rect 269 129 270 138
rect 253 129 254 140
rect 265 139 266 150
rect 284 129 285 140
rect 293 129 294 140
rect 253 141 254 150
rect 283 141 284 150
rect 287 129 288 142
rect 292 141 293 150
rect 263 129 264 144
rect 286 143 287 150
rect 290 129 291 144
rect 298 143 299 150
rect 272 129 273 146
rect 289 145 290 150
rect 271 147 272 150
rect 280 147 281 150
rect 301 147 302 150
rect 304 147 305 150
rect 310 147 311 150
rect 313 147 314 150
rect 238 154 239 157
rect 272 156 273 189
rect 251 158 252 189
rect 275 158 276 189
rect 253 154 254 161
rect 314 160 315 189
rect 256 154 257 163
rect 298 154 299 163
rect 268 154 269 165
rect 286 154 287 165
rect 229 154 230 167
rect 269 166 270 189
rect 280 154 281 167
rect 329 166 330 189
rect 283 154 284 169
rect 332 168 333 189
rect 284 170 285 189
rect 323 170 324 189
rect 289 154 290 173
rect 320 172 321 189
rect 292 154 293 175
rect 347 174 348 189
rect 241 176 242 189
rect 293 176 294 189
rect 295 154 296 177
rect 341 176 342 189
rect 244 178 245 189
rect 296 178 297 189
rect 301 154 302 179
rect 350 178 351 189
rect 308 180 309 189
rect 344 180 345 189
rect 310 154 311 183
rect 359 182 360 189
rect 265 154 266 185
rect 311 184 312 189
rect 235 154 236 187
rect 266 186 267 189
rect 372 186 373 189
rect 376 186 377 189
rect 220 195 221 246
rect 257 195 258 246
rect 234 197 235 246
rect 269 193 270 198
rect 231 199 232 246
rect 269 199 270 246
rect 241 201 242 246
rect 272 193 273 202
rect 245 203 246 246
rect 263 203 264 246
rect 248 205 249 246
rect 293 193 294 206
rect 251 193 252 208
rect 314 193 315 208
rect 266 207 267 246
rect 266 193 267 208
rect 272 209 273 246
rect 287 209 288 246
rect 278 211 279 246
rect 296 193 297 212
rect 281 213 282 246
rect 305 213 306 246
rect 284 193 285 216
rect 329 193 330 216
rect 275 193 276 218
rect 284 217 285 246
rect 290 217 291 246
rect 323 193 324 218
rect 302 219 303 246
rect 332 193 333 220
rect 308 193 309 222
rect 341 193 342 222
rect 308 223 309 246
rect 344 193 345 224
rect 311 223 312 246
rect 311 193 312 224
rect 317 193 318 226
rect 323 225 324 246
rect 317 227 318 246
rect 344 227 345 246
rect 320 193 321 230
rect 347 193 348 230
rect 332 231 333 246
rect 350 193 351 232
rect 338 233 339 246
rect 369 193 370 234
rect 341 235 342 246
rect 381 235 382 246
rect 350 237 351 246
rect 359 193 360 238
rect 356 239 357 246
rect 374 239 375 246
rect 368 241 369 246
rect 388 241 389 246
rect 371 243 372 246
rect 377 243 378 246
rect 217 250 218 253
rect 244 252 245 299
rect 220 250 221 255
rect 253 254 254 299
rect 231 256 232 299
rect 263 250 264 257
rect 248 250 249 259
rect 305 250 306 259
rect 266 250 267 261
rect 284 250 285 261
rect 257 250 258 263
rect 283 262 284 299
rect 256 264 257 299
rect 269 250 270 265
rect 241 250 242 267
rect 268 266 269 299
rect 272 250 273 267
rect 278 250 279 267
rect 241 268 242 299
rect 271 268 272 299
rect 275 250 276 269
rect 290 250 291 269
rect 287 250 288 271
rect 292 270 293 299
rect 302 250 303 271
rect 335 250 336 271
rect 281 250 282 273
rect 301 272 302 299
rect 234 250 235 275
rect 280 274 281 299
rect 227 250 228 277
rect 234 276 235 299
rect 308 250 309 277
rect 388 250 389 277
rect 323 250 324 279
rect 328 278 329 299
rect 331 278 332 299
rect 363 278 364 299
rect 338 250 339 281
rect 381 250 382 281
rect 325 282 326 299
rect 337 282 338 299
rect 341 250 342 283
rect 360 282 361 299
rect 344 250 345 285
rect 371 250 372 285
rect 347 250 348 287
rect 356 250 357 287
rect 347 288 348 299
rect 374 250 375 289
rect 350 250 351 291
rect 353 290 354 299
rect 317 250 318 293
rect 350 292 351 299
rect 304 294 305 299
rect 316 294 317 299
rect 368 250 369 295
rect 377 250 378 295
rect 370 296 371 299
rect 377 296 378 299
rect 220 303 221 306
rect 253 303 254 306
rect 224 303 225 308
rect 226 307 227 356
rect 223 309 224 356
rect 244 303 245 310
rect 231 303 232 312
rect 283 303 284 312
rect 234 303 235 314
rect 241 303 242 314
rect 238 303 239 316
rect 268 303 269 316
rect 240 317 241 356
rect 271 303 272 318
rect 243 319 244 356
rect 256 303 257 320
rect 256 321 257 356
rect 301 303 302 322
rect 259 323 260 356
rect 286 303 287 324
rect 262 325 263 356
rect 284 325 285 356
rect 272 327 273 356
rect 299 327 300 356
rect 277 303 278 330
rect 280 303 281 330
rect 269 331 270 356
rect 281 331 282 356
rect 289 303 290 332
rect 292 303 293 332
rect 302 331 303 356
rect 325 303 326 332
rect 305 333 306 356
rect 328 303 329 334
rect 314 335 315 356
rect 323 335 324 356
rect 316 303 317 338
rect 320 337 321 356
rect 317 339 318 356
rect 350 303 351 340
rect 331 303 332 342
rect 367 303 368 342
rect 334 303 335 344
rect 341 303 342 344
rect 333 345 334 356
rect 368 345 369 356
rect 345 347 346 356
rect 354 347 355 356
rect 347 303 348 350
rect 360 303 361 350
rect 336 351 337 356
rect 361 351 362 356
rect 348 353 349 356
rect 351 353 352 356
rect 230 360 231 363
rect 237 360 238 363
rect 238 364 239 405
rect 243 360 244 365
rect 246 360 247 365
rect 250 364 251 405
rect 235 366 236 405
rect 247 366 248 405
rect 256 360 257 367
rect 291 366 292 405
rect 259 360 260 369
rect 288 368 289 405
rect 269 360 270 371
rect 284 360 285 371
rect 272 360 273 373
rect 281 360 282 373
rect 260 374 261 405
rect 273 374 274 405
rect 267 376 268 405
rect 282 376 283 405
rect 299 360 300 377
rect 320 360 321 377
rect 265 360 266 379
rect 300 378 301 405
rect 297 380 298 405
rect 321 380 322 405
rect 302 360 303 383
rect 312 382 313 405
rect 262 360 263 385
rect 303 384 304 405
rect 263 386 264 405
rect 309 386 310 405
rect 305 360 306 389
rect 388 388 389 405
rect 270 390 271 405
rect 306 390 307 405
rect 314 360 315 391
rect 357 390 358 405
rect 327 360 328 393
rect 348 360 349 393
rect 317 360 318 395
rect 327 394 328 405
rect 333 360 334 395
rect 395 394 396 405
rect 330 360 331 397
rect 333 396 334 405
rect 336 360 337 397
rect 376 396 377 405
rect 339 398 340 405
rect 373 398 374 405
rect 345 360 346 401
rect 382 400 383 405
rect 360 402 361 405
rect 366 402 367 405
rect 379 402 380 405
rect 385 402 386 405
rect 235 409 236 412
rect 250 409 251 412
rect 235 413 236 456
rect 247 409 248 414
rect 242 415 243 456
rect 256 409 257 416
rect 253 409 254 418
rect 273 409 274 418
rect 260 409 261 420
rect 288 409 289 420
rect 263 409 264 422
rect 303 409 304 422
rect 263 423 264 456
rect 325 423 326 456
rect 267 409 268 426
rect 291 409 292 426
rect 256 427 257 456
rect 290 427 291 456
rect 275 429 276 456
rect 282 409 283 430
rect 278 431 279 456
rect 306 409 307 432
rect 287 433 288 456
rect 309 409 310 434
rect 312 409 313 434
rect 318 433 319 456
rect 312 435 313 456
rect 327 409 328 436
rect 315 409 316 438
rect 366 409 367 438
rect 315 439 316 456
rect 321 409 322 440
rect 321 441 322 456
rect 333 409 334 442
rect 332 443 333 456
rect 399 409 400 444
rect 339 409 340 446
rect 385 409 386 446
rect 357 409 358 448
rect 373 409 374 448
rect 360 409 361 450
rect 370 409 371 450
rect 376 409 377 450
rect 395 409 396 450
rect 379 409 380 452
rect 392 409 393 452
rect 382 409 383 454
rect 388 409 389 454
rect 238 460 239 463
rect 242 460 243 463
rect 256 460 257 463
rect 275 460 276 463
rect 256 464 257 477
rect 278 460 279 465
rect 259 460 260 467
rect 263 460 264 467
rect 266 460 267 467
rect 287 460 288 467
rect 253 468 254 477
rect 266 468 267 477
rect 269 468 270 477
rect 290 460 291 469
rect 282 470 283 477
rect 303 460 304 471
rect 286 472 287 477
rect 298 472 299 477
rect 301 472 302 477
rect 307 472 308 477
rect 312 460 313 473
rect 321 460 322 473
rect 315 460 316 475
rect 318 460 319 475
rect 328 460 329 475
rect 335 460 336 475
rect 256 481 257 484
rect 266 481 267 484
rect 260 481 261 486
rect 269 481 270 486
rect 271 485 272 494
rect 279 481 280 486
rect 274 487 275 494
rect 301 481 302 488
rect 280 489 281 494
rect 307 481 308 490
rect 298 481 299 492
rect 304 481 305 492
rect 271 498 272 501
rect 274 498 275 501
rect 280 498 281 501
rect 283 498 284 501
<< via >>
rect 247 113 248 114
rect 253 113 254 114
rect 250 115 251 116
rect 287 115 288 116
rect 262 117 263 118
rect 269 117 270 118
rect 266 119 267 120
rect 284 119 285 120
rect 272 121 273 122
rect 296 121 297 122
rect 229 131 230 132
rect 235 131 236 132
rect 232 133 233 134
rect 238 133 239 134
rect 247 133 248 134
rect 259 133 260 134
rect 250 135 251 136
rect 295 135 296 136
rect 266 137 267 138
rect 269 137 270 138
rect 253 139 254 140
rect 265 139 266 140
rect 284 139 285 140
rect 293 139 294 140
rect 253 141 254 142
rect 283 141 284 142
rect 287 141 288 142
rect 292 141 293 142
rect 263 143 264 144
rect 286 143 287 144
rect 290 143 291 144
rect 298 143 299 144
rect 272 145 273 146
rect 289 145 290 146
rect 271 147 272 148
rect 280 147 281 148
rect 301 147 302 148
rect 304 147 305 148
rect 310 147 311 148
rect 313 147 314 148
rect 238 156 239 157
rect 272 156 273 157
rect 251 158 252 159
rect 275 158 276 159
rect 253 160 254 161
rect 314 160 315 161
rect 256 162 257 163
rect 298 162 299 163
rect 268 164 269 165
rect 286 164 287 165
rect 229 166 230 167
rect 269 166 270 167
rect 280 166 281 167
rect 329 166 330 167
rect 283 168 284 169
rect 332 168 333 169
rect 284 170 285 171
rect 323 170 324 171
rect 289 172 290 173
rect 320 172 321 173
rect 292 174 293 175
rect 347 174 348 175
rect 241 176 242 177
rect 293 176 294 177
rect 295 176 296 177
rect 341 176 342 177
rect 244 178 245 179
rect 296 178 297 179
rect 301 178 302 179
rect 350 178 351 179
rect 308 180 309 181
rect 344 180 345 181
rect 310 182 311 183
rect 359 182 360 183
rect 265 184 266 185
rect 311 184 312 185
rect 235 186 236 187
rect 266 186 267 187
rect 372 186 373 187
rect 376 186 377 187
rect 220 195 221 196
rect 257 195 258 196
rect 234 197 235 198
rect 269 197 270 198
rect 231 199 232 200
rect 269 199 270 200
rect 241 201 242 202
rect 272 201 273 202
rect 245 203 246 204
rect 263 203 264 204
rect 248 205 249 206
rect 293 205 294 206
rect 251 207 252 208
rect 314 207 315 208
rect 272 209 273 210
rect 287 209 288 210
rect 278 211 279 212
rect 296 211 297 212
rect 281 213 282 214
rect 305 213 306 214
rect 284 215 285 216
rect 329 215 330 216
rect 275 217 276 218
rect 284 217 285 218
rect 290 217 291 218
rect 323 217 324 218
rect 302 219 303 220
rect 332 219 333 220
rect 308 221 309 222
rect 341 221 342 222
rect 308 223 309 224
rect 344 223 345 224
rect 317 225 318 226
rect 323 225 324 226
rect 317 227 318 228
rect 344 227 345 228
rect 320 229 321 230
rect 347 229 348 230
rect 332 231 333 232
rect 350 231 351 232
rect 338 233 339 234
rect 369 233 370 234
rect 341 235 342 236
rect 381 235 382 236
rect 350 237 351 238
rect 359 237 360 238
rect 356 239 357 240
rect 374 239 375 240
rect 368 241 369 242
rect 388 241 389 242
rect 371 243 372 244
rect 377 243 378 244
rect 217 252 218 253
rect 244 252 245 253
rect 220 254 221 255
rect 253 254 254 255
rect 231 256 232 257
rect 263 256 264 257
rect 248 258 249 259
rect 305 258 306 259
rect 266 260 267 261
rect 284 260 285 261
rect 257 262 258 263
rect 283 262 284 263
rect 256 264 257 265
rect 269 264 270 265
rect 241 266 242 267
rect 268 266 269 267
rect 272 266 273 267
rect 278 266 279 267
rect 241 268 242 269
rect 271 268 272 269
rect 275 268 276 269
rect 290 268 291 269
rect 287 270 288 271
rect 292 270 293 271
rect 302 270 303 271
rect 335 270 336 271
rect 281 272 282 273
rect 301 272 302 273
rect 234 274 235 275
rect 280 274 281 275
rect 227 276 228 277
rect 234 276 235 277
rect 308 276 309 277
rect 388 276 389 277
rect 323 278 324 279
rect 328 278 329 279
rect 331 278 332 279
rect 363 278 364 279
rect 338 280 339 281
rect 381 280 382 281
rect 325 282 326 283
rect 337 282 338 283
rect 341 282 342 283
rect 360 282 361 283
rect 344 284 345 285
rect 371 284 372 285
rect 347 286 348 287
rect 356 286 357 287
rect 347 288 348 289
rect 374 288 375 289
rect 350 290 351 291
rect 353 290 354 291
rect 317 292 318 293
rect 350 292 351 293
rect 304 294 305 295
rect 316 294 317 295
rect 368 294 369 295
rect 377 294 378 295
rect 370 296 371 297
rect 377 296 378 297
rect 220 305 221 306
rect 253 305 254 306
rect 224 307 225 308
rect 226 307 227 308
rect 223 309 224 310
rect 244 309 245 310
rect 231 311 232 312
rect 283 311 284 312
rect 234 313 235 314
rect 241 313 242 314
rect 238 315 239 316
rect 268 315 269 316
rect 240 317 241 318
rect 271 317 272 318
rect 243 319 244 320
rect 256 319 257 320
rect 256 321 257 322
rect 301 321 302 322
rect 259 323 260 324
rect 286 323 287 324
rect 262 325 263 326
rect 284 325 285 326
rect 272 327 273 328
rect 299 327 300 328
rect 277 329 278 330
rect 280 329 281 330
rect 269 331 270 332
rect 281 331 282 332
rect 289 331 290 332
rect 292 331 293 332
rect 302 331 303 332
rect 325 331 326 332
rect 305 333 306 334
rect 328 333 329 334
rect 314 335 315 336
rect 323 335 324 336
rect 316 337 317 338
rect 320 337 321 338
rect 317 339 318 340
rect 350 339 351 340
rect 331 341 332 342
rect 367 341 368 342
rect 334 343 335 344
rect 341 343 342 344
rect 333 345 334 346
rect 368 345 369 346
rect 345 347 346 348
rect 354 347 355 348
rect 347 349 348 350
rect 360 349 361 350
rect 336 351 337 352
rect 361 351 362 352
rect 348 353 349 354
rect 351 353 352 354
rect 230 362 231 363
rect 237 362 238 363
rect 238 364 239 365
rect 243 364 244 365
rect 246 364 247 365
rect 250 364 251 365
rect 235 366 236 367
rect 247 366 248 367
rect 256 366 257 367
rect 291 366 292 367
rect 259 368 260 369
rect 288 368 289 369
rect 269 370 270 371
rect 284 370 285 371
rect 272 372 273 373
rect 281 372 282 373
rect 260 374 261 375
rect 273 374 274 375
rect 267 376 268 377
rect 282 376 283 377
rect 299 376 300 377
rect 320 376 321 377
rect 265 378 266 379
rect 300 378 301 379
rect 297 380 298 381
rect 321 380 322 381
rect 302 382 303 383
rect 312 382 313 383
rect 262 384 263 385
rect 303 384 304 385
rect 263 386 264 387
rect 309 386 310 387
rect 305 388 306 389
rect 388 388 389 389
rect 270 390 271 391
rect 306 390 307 391
rect 314 390 315 391
rect 357 390 358 391
rect 327 392 328 393
rect 348 392 349 393
rect 317 394 318 395
rect 327 394 328 395
rect 333 394 334 395
rect 395 394 396 395
rect 330 396 331 397
rect 333 396 334 397
rect 336 396 337 397
rect 376 396 377 397
rect 339 398 340 399
rect 373 398 374 399
rect 345 400 346 401
rect 382 400 383 401
rect 360 402 361 403
rect 366 402 367 403
rect 379 402 380 403
rect 385 402 386 403
rect 235 411 236 412
rect 250 411 251 412
rect 235 413 236 414
rect 247 413 248 414
rect 242 415 243 416
rect 256 415 257 416
rect 253 417 254 418
rect 273 417 274 418
rect 260 419 261 420
rect 288 419 289 420
rect 263 421 264 422
rect 303 421 304 422
rect 263 423 264 424
rect 325 423 326 424
rect 267 425 268 426
rect 291 425 292 426
rect 256 427 257 428
rect 290 427 291 428
rect 275 429 276 430
rect 282 429 283 430
rect 278 431 279 432
rect 306 431 307 432
rect 287 433 288 434
rect 309 433 310 434
rect 312 433 313 434
rect 318 433 319 434
rect 312 435 313 436
rect 327 435 328 436
rect 315 437 316 438
rect 366 437 367 438
rect 315 439 316 440
rect 321 439 322 440
rect 321 441 322 442
rect 333 441 334 442
rect 332 443 333 444
rect 399 443 400 444
rect 339 445 340 446
rect 385 445 386 446
rect 357 447 358 448
rect 373 447 374 448
rect 360 449 361 450
rect 370 449 371 450
rect 376 449 377 450
rect 395 449 396 450
rect 379 451 380 452
rect 392 451 393 452
rect 382 453 383 454
rect 388 453 389 454
rect 238 462 239 463
rect 242 462 243 463
rect 256 462 257 463
rect 275 462 276 463
rect 256 464 257 465
rect 278 464 279 465
rect 259 466 260 467
rect 263 466 264 467
rect 266 466 267 467
rect 287 466 288 467
rect 253 468 254 469
rect 266 468 267 469
rect 269 468 270 469
rect 290 468 291 469
rect 282 470 283 471
rect 303 470 304 471
rect 286 472 287 473
rect 298 472 299 473
rect 301 472 302 473
rect 307 472 308 473
rect 312 472 313 473
rect 321 472 322 473
rect 315 474 316 475
rect 318 474 319 475
rect 328 474 329 475
rect 335 474 336 475
rect 256 483 257 484
rect 266 483 267 484
rect 260 485 261 486
rect 269 485 270 486
rect 271 485 272 486
rect 279 485 280 486
rect 274 487 275 488
rect 301 487 302 488
rect 280 489 281 490
rect 307 489 308 490
rect 298 491 299 492
rect 304 491 305 492
rect 271 500 272 501
rect 274 500 275 501
rect 280 500 281 501
rect 283 500 284 501
<< end >>
