magic
tech scmos
timestamp 1394680307
<< m1p >>
use CELL  1
transform -1 0 511 0 1 516
box 0 0 6 6
use CELL  2
transform -1 0 487 0 -1 594
box 0 0 6 6
use CELL  3
transform 1 0 509 0 1 552
box 0 0 6 6
use CELL  4
transform -1 0 494 0 1 588
box 0 0 6 6
use CELL  5
transform -1 0 521 0 1 624
box 0 0 6 6
use CELL  6
transform 1 0 521 0 1 612
box 0 0 6 6
use CELL  7
transform -1 0 606 0 1 516
box 0 0 6 6
use CELL  8
transform -1 0 523 0 1 504
box 0 0 6 6
use CELL  9
transform -1 0 513 0 1 588
box 0 0 6 6
use CELL  10
transform 1 0 644 0 1 588
box 0 0 6 6
use CELL  11
transform -1 0 634 0 1 564
box 0 0 6 6
use CELL  12
transform -1 0 609 0 1 504
box 0 0 6 6
use CELL  13
transform 1 0 532 0 -1 582
box 0 0 6 6
use CELL  14
transform -1 0 498 0 1 540
box 0 0 6 6
use CELL  15
transform -1 0 504 0 1 516
box 0 0 6 6
use CELL  16
transform -1 0 589 0 1 504
box 0 0 6 6
use CELL  17
transform -1 0 529 0 1 480
box 0 0 6 6
use CELL  18
transform -1 0 516 0 -1 510
box 0 0 6 6
use CELL  19
transform -1 0 494 0 1 600
box 0 0 6 6
use CELL  20
transform -1 0 535 0 1 480
box 0 0 6 6
use CELL  21
transform -1 0 576 0 -1 546
box 0 0 6 6
use CELL  22
transform -1 0 542 0 -1 486
box 0 0 6 6
use CELL  23
transform 1 0 480 0 1 504
box 0 0 6 6
use CELL  24
transform 1 0 489 0 1 516
box 0 0 6 6
use CELL  25
transform -1 0 577 0 -1 534
box 0 0 6 6
use CELL  26
transform 1 0 522 0 -1 630
box 0 0 6 6
use CELL  27
transform -1 0 613 0 1 516
box 0 0 6 6
use CELL  28
transform -1 0 495 0 1 576
box 0 0 6 6
use CELL  29
transform 1 0 544 0 -1 510
box 0 0 6 6
use CELL  30
transform -1 0 584 0 1 528
box 0 0 6 6
use CELL  31
transform -1 0 628 0 1 540
box 0 0 6 6
use CELL  32
transform 1 0 492 0 -1 486
box 0 0 6 6
use CELL  33
transform -1 0 493 0 1 504
box 0 0 6 6
use CELL  34
transform -1 0 523 0 1 492
box 0 0 6 6
use CELL  35
transform 1 0 641 0 1 528
box 0 0 6 6
use CELL  36
transform -1 0 556 0 1 564
box 0 0 6 6
use CELL  37
transform -1 0 510 0 1 540
box 0 0 6 6
use CELL  38
transform -1 0 592 0 1 588
box 0 0 6 6
use CELL  39
transform -1 0 487 0 1 600
box 0 0 6 6
use CELL  40
transform -1 0 506 0 1 612
box 0 0 6 6
use CELL  41
transform 1 0 583 0 -1 606
box 0 0 6 6
use CELL  42
transform -1 0 486 0 1 540
box 0 0 6 6
use CELL  43
transform -1 0 501 0 1 600
box 0 0 6 6
use CELL  44
transform -1 0 494 0 1 564
box 0 0 6 6
use CELL  45
transform -1 0 518 0 1 612
box 0 0 6 6
use CELL  46
transform 1 0 474 0 1 528
box 0 0 6 6
use CELL  47
transform -1 0 629 0 1 576
box 0 0 6 6
use CELL  48
transform 1 0 615 0 1 552
box 0 0 6 6
use CELL  49
transform -1 0 690 0 1 576
box 0 0 6 6
use CELL  50
transform -1 0 511 0 1 528
box 0 0 6 6
use CELL  51
transform -1 0 534 0 1 612
box 0 0 6 6
use CELL  52
transform 1 0 653 0 1 564
box 0 0 6 6
use CELL  53
transform -1 0 541 0 1 504
box 0 0 6 6
use CELL  54
transform -1 0 480 0 1 600
box 0 0 6 6
use CELL  55
transform -1 0 564 0 1 504
box 0 0 6 6
use CELL  56
transform -1 0 633 0 1 528
box 0 0 6 6
use CELL  57
transform -1 0 522 0 1 480
box 0 0 6 6
use CELL  58
transform 1 0 699 0 -1 582
box 0 0 6 6
use CELL  59
transform -1 0 664 0 1 588
box 0 0 6 6
use CELL  60
transform -1 0 515 0 1 600
box 0 0 6 6
use CELL  61
transform -1 0 656 0 -1 558
box 0 0 6 6
use CELL  62
transform 1 0 572 0 1 492
box 0 0 6 6
use CELL  63
transform -1 0 480 0 1 564
box 0 0 6 6
use CELL  64
transform 1 0 651 0 1 540
box 0 0 6 6
use CELL  65
transform -1 0 583 0 1 588
box 0 0 6 6
use CELL  66
transform -1 0 699 0 1 576
box 0 0 6 6
use CELL  67
transform 1 0 576 0 1 504
box 0 0 6 6
use CELL  68
transform -1 0 643 0 1 588
box 0 0 6 6
use CELL  69
transform -1 0 492 0 1 528
box 0 0 6 6
use CELL  70
transform -1 0 480 0 1 492
box 0 0 6 6
use CELL  71
transform -1 0 532 0 1 492
box 0 0 6 6
use CELL  72
transform 1 0 634 0 1 552
box 0 0 6 6
use CELL  73
transform 1 0 576 0 1 612
box 0 0 6 6
use CELL  74
transform 1 0 492 0 1 624
box 0 0 6 6
use CELL  75
transform -1 0 573 0 1 504
box 0 0 6 6
use CELL  76
transform -1 0 493 0 1 492
box 0 0 6 6
use CELL  77
transform -1 0 557 0 1 504
box 0 0 6 6
use CELL  78
transform -1 0 522 0 1 540
box 0 0 6 6
use CELL  79
transform -1 0 508 0 1 552
box 0 0 6 6
use CELL  80
transform -1 0 583 0 1 516
box 0 0 6 6
use CELL  81
transform 1 0 488 0 -1 558
box 0 0 6 6
use CELL  82
transform -1 0 558 0 1 552
box 0 0 6 6
use CELL  83
transform -1 0 488 0 -1 582
box 0 0 6 6
use CELL  84
transform -1 0 553 0 1 588
box 0 0 6 6
use CELL  85
transform -1 0 481 0 1 576
box 0 0 6 6
use CELL  86
transform -1 0 564 0 1 540
box 0 0 6 6
use CELL  87
transform -1 0 487 0 1 552
box 0 0 6 6
use CELL  88
transform -1 0 474 0 1 576
box 0 0 6 6
use CELL  89
transform -1 0 535 0 1 516
box 0 0 6 6
use CELL  90
transform -1 0 545 0 1 576
box 0 0 6 6
use CELL  91
transform 1 0 651 0 1 588
box 0 0 6 6
use CELL  92
transform -1 0 649 0 1 552
box 0 0 6 6
use CELL  93
transform -1 0 507 0 1 576
box 0 0 6 6
use CELL  94
transform -1 0 590 0 1 516
box 0 0 6 6
use CELL  95
transform -1 0 574 0 1 516
box 0 0 6 6
use CELL  96
transform -1 0 636 0 -1 522
box 0 0 6 6
use CELL  97
transform -1 0 591 0 1 528
box 0 0 6 6
use CELL  98
transform -1 0 661 0 1 576
box 0 0 6 6
use CELL  99
transform -1 0 514 0 -1 630
box 0 0 6 6
use CELL  100
transform -1 0 509 0 1 504
box 0 0 6 6
use CELL  101
transform -1 0 500 0 1 504
box 0 0 6 6
use CELL  102
transform 1 0 495 0 1 564
box 0 0 6 6
use CELL  103
transform -1 0 622 0 1 564
box 0 0 6 6
use CELL  104
transform -1 0 515 0 1 564
box 0 0 6 6
use CELL  105
transform -1 0 588 0 1 612
box 0 0 6 6
use CELL  106
transform 1 0 623 0 1 516
box 0 0 6 6
use CELL  107
transform -1 0 505 0 1 624
box 0 0 6 6
use CELL  108
transform 1 0 593 0 1 516
box 0 0 6 6
use CELL  109
transform 1 0 670 0 1 576
box 0 0 6 6
use CELL  110
transform 1 0 517 0 1 636
box 0 0 6 6
use CELL  111
transform -1 0 617 0 1 576
box 0 0 6 6
use CELL  112
transform -1 0 564 0 1 492
box 0 0 6 6
use CELL  113
transform -1 0 596 0 1 504
box 0 0 6 6
use CELL  114
transform -1 0 645 0 1 516
box 0 0 6 6
use CELL  115
transform -1 0 666 0 1 540
box 0 0 6 6
use CELL  116
transform -1 0 568 0 1 612
box 0 0 6 6
use CELL  117
transform 1 0 585 0 1 492
box 0 0 6 6
use CELL  118
transform -1 0 650 0 1 540
box 0 0 6 6
use CELL  119
transform -1 0 552 0 1 540
box 0 0 6 6
use CELL  120
transform -1 0 616 0 1 504
box 0 0 6 6
use CELL  121
transform -1 0 550 0 1 492
box 0 0 6 6
use CELL  122
transform -1 0 487 0 1 564
box 0 0 6 6
use CELL  123
transform -1 0 549 0 1 564
box 0 0 6 6
use CELL  124
transform -1 0 609 0 1 540
box 0 0 6 6
use CELL  125
transform -1 0 712 0 1 576
box 0 0 6 6
use CELL  126
transform -1 0 582 0 1 552
box 0 0 6 6
use CELL  127
transform -1 0 487 0 1 492
box 0 0 6 6
use CELL  128
transform 1 0 659 0 -1 558
box 0 0 6 6
use CELL  129
transform -1 0 566 0 1 600
box 0 0 6 6
use CELL  130
transform -1 0 531 0 1 564
box 0 0 6 6
use CELL  131
transform -1 0 516 0 1 636
box 0 0 6 6
use CELL  132
transform -1 0 621 0 1 540
box 0 0 6 6
use CELL  133
transform -1 0 596 0 1 600
box 0 0 6 6
use CELL  134
transform -1 0 546 0 1 588
box 0 0 6 6
use CELL  135
transform -1 0 603 0 1 600
box 0 0 6 6
use CELL  136
transform -1 0 486 0 1 516
box 0 0 6 6
use CELL  137
transform -1 0 531 0 1 588
box 0 0 6 6
use CELL  138
transform -1 0 504 0 1 528
box 0 0 6 6
use CELL  139
transform -1 0 527 0 1 552
box 0 0 6 6
use CELL  140
transform -1 0 603 0 1 504
box 0 0 6 6
use CELL  141
transform -1 0 508 0 1 564
box 0 0 6 6
use CELL  142
transform -1 0 647 0 1 576
box 0 0 6 6
use CELL  143
transform -1 0 480 0 1 588
box 0 0 6 6
use CELL  144
transform -1 0 480 0 1 552
box 0 0 6 6
use CELL  145
transform -1 0 561 0 1 612
box 0 0 6 6
use CELL  146
transform -1 0 508 0 1 600
box 0 0 6 6
use CELL  147
transform 1 0 622 0 1 552
box 0 0 6 6
use CELL  148
transform -1 0 613 0 1 564
box 0 0 6 6
use CELL  149
transform -1 0 643 0 1 540
box 0 0 6 6
use CELL  150
transform 1 0 620 0 -1 534
box 0 0 6 6
use CELL  151
transform -1 0 619 0 1 528
box 0 0 6 6
use CELL  152
transform -1 0 598 0 1 528
box 0 0 6 6
use CELL  153
transform -1 0 550 0 1 528
box 0 0 6 6
use CELL  154
transform -1 0 575 0 1 612
box 0 0 6 6
use CELL  155
transform -1 0 622 0 -1 522
box 0 0 6 6
use CELL  156
transform 1 0 510 0 1 492
box 0 0 6 6
use CELL  157
transform 1 0 667 0 1 540
box 0 0 6 6
use CELL  158
transform -1 0 573 0 1 600
box 0 0 6 6
use CELL  159
transform -1 0 501 0 1 588
box 0 0 6 6
use CELL  160
transform -1 0 589 0 1 564
box 0 0 6 6
use CELL  161
transform -1 0 519 0 1 576
box 0 0 6 6
use CELL  162
transform -1 0 527 0 1 600
box 0 0 6 6
use CELL  163
transform -1 0 683 0 1 576
box 0 0 6 6
use CELL  164
transform -1 0 619 0 -1 594
box 0 0 6 6
use CELL  165
transform -1 0 501 0 1 552
box 0 0 6 6
use CELL  166
transform -1 0 654 0 1 576
box 0 0 6 6
use CELL  167
transform -1 0 492 0 1 612
box 0 0 6 6
use CELL  168
transform -1 0 610 0 1 588
box 0 0 6 6
use CELL  169
transform -1 0 640 0 1 528
box 0 0 6 6
use CELL  170
transform -1 0 526 0 1 576
box 0 0 6 6
use CELL  171
transform -1 0 522 0 1 564
box 0 0 6 6
use CELL  172
transform -1 0 580 0 1 600
box 0 0 6 6
use CELL  173
transform -1 0 652 0 1 564
box 0 0 6 6
use CELL  174
transform 1 0 565 0 1 492
box 0 0 6 6
use CELL  175
transform 1 0 551 0 1 492
box 0 0 6 6
use CELL  176
transform 1 0 493 0 -1 618
box 0 0 6 6
use CELL  177
transform 1 0 578 0 -1 498
box 0 0 6 6
use CELL  178
transform 1 0 625 0 1 588
box 0 0 6 6
use CELL  179
transform -1 0 609 0 1 552
box 0 0 6 6
use CELL  180
transform -1 0 534 0 1 552
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 540 0 1 540
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 529 0 1 528
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 575 0 1 576
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 552 0 1 612
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 542 0 1 600
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 574 0 1 588
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 569 0 1 576
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 559 0 1 564
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 549 0 1 552
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 540 0 1 612
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 539 0 1 600
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 571 0 1 588
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 554 0 1 576
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 537 0 1 564
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 549 0 1 612
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 564 0 1 504
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 607 0 1 528
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 610 0 1 528
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 609 0 1 540
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 565 0 1 516
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 603 0 1 600
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 628 0 1 552
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 628 0 1 540
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 661 0 1 576
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 631 0 1 588
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 636 0 1 516
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 647 0 1 528
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 657 0 1 540
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 656 0 1 552
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 665 0 1 564
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 690 0 1 576
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 500 0 1 504
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 613 0 1 516
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 523 0 1 492
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 541 0 1 504
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 574 0 1 516
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 511 0 1 516
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 526 0 1 528
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 543 0 1 540
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 543 0 1 552
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 562 0 1 588
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 507 0 1 576
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 506 0 1 612
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 538 0 1 492
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 541 0 1 492
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 553 0 1 528
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 544 0 1 516
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 529 0 1 504
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 546 0 1 612
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 551 0 1 600
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 547 0 1 516
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 486 0 1 516
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 492 0 1 528
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 501 0 1 540
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 532 0 1 504
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 517 0 1 516
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 556 0 1 528
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 608 0 1 576
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 596 0 1 576
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 495 0 1 528
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 495 0 1 516
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 578 0 1 576
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 598 0 1 564
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 591 0 1 552
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 579 0 1 540
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 587 0 1 576
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 568 0 1 564
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 515 0 1 600
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 534 0 1 588
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 526 0 1 576
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 513 0 1 588
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 505 0 1 624
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 659 0 1 564
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 523 0 1 516
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 550 0 1 516
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 559 0 1 528
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 612 0 1 540
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 597 0 1 552
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 667 0 1 576
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 662 0 1 564
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 640 0 1 552
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 634 0 1 540
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 604 0 1 528
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 590 0 1 516
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 573 0 1 504
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 537 0 1 588
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 554 0 1 600
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 584 0 1 576
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 574 0 1 564
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 664 0 1 576
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 640 0 1 564
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 498 0 1 540
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 643 0 1 564
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 509 0 1 612
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 559 0 1 516
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 562 0 1 516
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 565 0 1 528
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 588 0 1 540
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 600 0 1 552
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 541 0 1 516
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 550 0 1 528
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 525 0 1 540
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 532 0 1 528
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 522 0 1 564
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 566 0 1 576
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 533 0 1 600
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 553 0 1 588
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 556 0 1 564
box 0 0 3 6
use FEEDTHRU  F-109
transform 1 0 546 0 1 552
box 0 0 3 6
use FEEDTHRU  F-110
transform 1 0 555 0 1 540
box 0 0 3 6
use FEEDTHRU  F-111
transform 1 0 573 0 1 552
box 0 0 3 6
use FEEDTHRU  F-112
transform 1 0 514 0 1 516
box 0 0 3 6
use FEEDTHRU  F-113
transform 1 0 511 0 1 528
box 0 0 3 6
use FEEDTHRU  F-114
transform 1 0 522 0 1 540
box 0 0 3 6
use FEEDTHRU  F-115
transform 1 0 545 0 1 576
box 0 0 3 6
use FEEDTHRU  F-116
transform 1 0 531 0 1 588
box 0 0 3 6
use FEEDTHRU  F-117
transform 1 0 620 0 1 576
box 0 0 3 6
use FEEDTHRU  F-118
transform 1 0 610 0 1 588
box 0 0 3 6
use FEEDTHRU  F-119
transform 1 0 540 0 1 552
box 0 0 3 6
use FEEDTHRU  F-120
transform 1 0 534 0 1 540
box 0 0 3 6
use FEEDTHRU  F-121
transform 1 0 520 0 1 528
box 0 0 3 6
use FEEDTHRU  F-122
transform 1 0 580 0 1 600
box 0 0 3 6
use FEEDTHRU  F-123
transform 1 0 634 0 1 588
box 0 0 3 6
use FEEDTHRU  F-124
transform 1 0 629 0 1 576
box 0 0 3 6
use FEEDTHRU  F-125
transform 1 0 622 0 1 564
box 0 0 3 6
use FEEDTHRU  F-126
transform 1 0 631 0 1 552
box 0 0 3 6
use FEEDTHRU  F-127
transform 1 0 631 0 1 540
box 0 0 3 6
use FEEDTHRU  F-128
transform 1 0 568 0 1 528
box 0 0 3 6
use FEEDTHRU  F-129
transform 1 0 518 0 1 612
box 0 0 3 6
use FEEDTHRU  F-130
transform 1 0 583 0 1 588
box 0 0 3 6
use FEEDTHRU  F-131
transform 1 0 557 0 1 600
box 0 0 3 6
use FEEDTHRU  F-132
transform 1 0 601 0 1 588
box 0 0 3 6
use FEEDTHRU  F-133
transform 1 0 599 0 1 576
box 0 0 3 6
use FEEDTHRU  F-134
transform 1 0 570 0 1 552
box 0 0 3 6
use FEEDTHRU  F-135
transform 1 0 577 0 1 564
box 0 0 3 6
use FEEDTHRU  F-136
transform 1 0 605 0 1 576
box 0 0 3 6
use FEEDTHRU  F-137
transform 1 0 598 0 1 588
box 0 0 3 6
use FEEDTHRU  F-138
transform 1 0 552 0 1 540
box 0 0 3 6
use FEEDTHRU  F-139
transform 1 0 604 0 1 564
box 0 0 3 6
use FEEDTHRU  F-140
transform 1 0 582 0 1 540
box 0 0 3 6
use FEEDTHRU  F-141
transform 1 0 594 0 1 552
box 0 0 3 6
use FEEDTHRU  F-142
transform 1 0 601 0 1 564
box 0 0 3 6
use FEEDTHRU  F-143
transform 1 0 617 0 1 576
box 0 0 3 6
use FEEDTHRU  F-144
transform 1 0 576 0 1 540
box 0 0 3 6
use FEEDTHRU  F-145
transform 1 0 588 0 1 552
box 0 0 3 6
use FEEDTHRU  F-146
transform 1 0 595 0 1 564
box 0 0 3 6
use FEEDTHRU  F-147
transform 1 0 613 0 1 564
box 0 0 3 6
use FEEDTHRU  F-148
transform 1 0 518 0 1 600
box 0 0 3 6
use FEEDTHRU  F-149
transform 1 0 559 0 1 588
box 0 0 3 6
use FEEDTHRU  F-150
transform 1 0 572 0 1 576
box 0 0 3 6
<< end >>
