magic
tech scmos
timestamp 1394680308
<< m1p >>
use CELL  1
transform -1 0 2240 0 1 2076
box 0 0 6 6
use CELL  2
transform 1 0 2060 0 1 2172
box 0 0 6 6
use CELL  3
transform 1 0 2707 0 1 2232
box 0 0 6 6
use CELL  4
transform 1 0 2124 0 -1 2034
box 0 0 6 6
use CELL  5
transform -1 0 2077 0 1 2112
box 0 0 6 6
use CELL  6
transform -1 0 2638 0 1 2256
box 0 0 6 6
use CELL  7
transform 1 0 2101 0 1 2028
box 0 0 6 6
use CELL  8
transform -1 0 2631 0 1 2148
box 0 0 6 6
use CELL  9
transform -1 0 2243 0 1 2304
box 0 0 6 6
use CELL  10
transform 1 0 2082 0 1 2040
box 0 0 6 6
use CELL  11
transform -1 0 2695 0 1 2268
box 0 0 6 6
use CELL  12
transform -1 0 2132 0 1 2184
box 0 0 6 6
use CELL  13
transform -1 0 2344 0 1 2100
box 0 0 6 6
use CELL  14
transform -1 0 2647 0 1 2268
box 0 0 6 6
use CELL  15
transform -1 0 2073 0 1 2148
box 0 0 6 6
use CELL  16
transform -1 0 2099 0 1 2172
box 0 0 6 6
use CELL  17
transform -1 0 2372 0 -1 2226
box 0 0 6 6
use CELL  18
transform 1 0 2132 0 -1 2082
box 0 0 6 6
use CELL  19
transform -1 0 2593 0 1 2196
box 0 0 6 6
use CELL  20
transform -1 0 2678 0 1 2160
box 0 0 6 6
use CELL  21
transform 1 0 2278 0 1 2040
box 0 0 6 6
use CELL  22
transform -1 0 2691 0 -1 2262
box 0 0 6 6
use CELL  23
transform -1 0 2086 0 1 2232
box 0 0 6 6
use CELL  24
transform -1 0 2116 0 1 2304
box 0 0 6 6
use CELL  25
transform 1 0 2271 0 1 2040
box 0 0 6 6
use CELL  26
transform -1 0 2598 0 1 2112
box 0 0 6 6
use CELL  27
transform -1 0 2186 0 1 2088
box 0 0 6 6
use CELL  28
transform -1 0 2384 0 1 2148
box 0 0 6 6
use CELL  29
transform -1 0 2126 0 1 2256
box 0 0 6 6
use CELL  30
transform -1 0 2098 0 1 2196
box 0 0 6 6
use CELL  31
transform -1 0 2098 0 1 2136
box 0 0 6 6
use CELL  32
transform -1 0 2441 0 1 2076
box 0 0 6 6
use CELL  33
transform -1 0 2606 0 1 2220
box 0 0 6 6
use CELL  34
transform -1 0 2206 0 1 2292
box 0 0 6 6
use CELL  35
transform -1 0 2479 0 1 2172
box 0 0 6 6
use CELL  36
transform -1 0 2059 0 1 2172
box 0 0 6 6
use CELL  37
transform 1 0 2644 0 -1 2250
box 0 0 6 6
use CELL  38
transform -1 0 2052 0 1 2172
box 0 0 6 6
use CELL  39
transform -1 0 2454 0 1 2172
box 0 0 6 6
use CELL  40
transform -1 0 2148 0 1 2208
box 0 0 6 6
use CELL  41
transform -1 0 2095 0 1 2304
box 0 0 6 6
use CELL  42
transform 1 0 2608 0 1 2196
box 0 0 6 6
use CELL  43
transform -1 0 2236 0 1 2220
box 0 0 6 6
use CELL  44
transform -1 0 2034 0 -1 2286
box 0 0 6 6
use CELL  45
transform -1 0 2132 0 1 2064
box 0 0 6 6
use CELL  46
transform 1 0 2347 0 -1 2070
box 0 0 6 6
use CELL  47
transform -1 0 2112 0 1 2196
box 0 0 6 6
use CELL  48
transform -1 0 2077 0 1 2088
box 0 0 6 6
use CELL  49
transform -1 0 2157 0 1 2328
box 0 0 6 6
use CELL  50
transform -1 0 2190 0 1 2028
box 0 0 6 6
use CELL  51
transform -1 0 2362 0 1 2304
box 0 0 6 6
use CELL  52
transform -1 0 2209 0 1 2196
box 0 0 6 6
use CELL  53
transform 1 0 2450 0 1 2292
box 0 0 6 6
use CELL  54
transform -1 0 2066 0 1 2160
box 0 0 6 6
use CELL  55
transform -1 0 2733 0 1 2232
box 0 0 6 6
use CELL  56
transform -1 0 2671 0 -1 2166
box 0 0 6 6
use CELL  57
transform 1 0 2064 0 -1 2094
box 0 0 6 6
use CELL  58
transform 1 0 2403 0 1 2076
box 0 0 6 6
use CELL  59
transform -1 0 2688 0 1 2244
box 0 0 6 6
use CELL  60
transform -1 0 2113 0 1 2328
box 0 0 6 6
use CELL  61
transform -1 0 2248 0 1 2244
box 0 0 6 6
use CELL  62
transform -1 0 2598 0 1 2136
box 0 0 6 6
use CELL  63
transform 1 0 2052 0 -1 2226
box 0 0 6 6
use CELL  64
transform -1 0 2304 0 -1 2046
box 0 0 6 6
use CELL  65
transform -1 0 2229 0 1 2280
box 0 0 6 6
use CELL  66
transform 1 0 2111 0 1 2088
box 0 0 6 6
use CELL  67
transform -1 0 2684 0 1 2256
box 0 0 6 6
use CELL  68
transform -1 0 2100 0 1 2232
box 0 0 6 6
use CELL  69
transform -1 0 2518 0 1 2184
box 0 0 6 6
use CELL  70
transform 1 0 2659 0 -1 2226
box 0 0 6 6
use CELL  71
transform -1 0 2620 0 1 2244
box 0 0 6 6
use CELL  72
transform -1 0 2432 0 1 2292
box 0 0 6 6
use CELL  73
transform -1 0 2273 0 -1 2310
box 0 0 6 6
use CELL  74
transform 1 0 2382 0 1 2076
box 0 0 6 6
use CELL  75
transform -1 0 2547 0 1 2112
box 0 0 6 6
use CELL  76
transform -1 0 2564 0 1 2232
box 0 0 6 6
use CELL  77
transform -1 0 2686 0 1 2196
box 0 0 6 6
use CELL  78
transform -1 0 2237 0 1 2064
box 0 0 6 6
use CELL  79
transform -1 0 2610 0 1 2268
box 0 0 6 6
use CELL  80
transform -1 0 2065 0 1 2220
box 0 0 6 6
use CELL  81
transform 1 0 2054 0 1 2124
box 0 0 6 6
use CELL  82
transform -1 0 2143 0 -1 2334
box 0 0 6 6
use CELL  83
transform -1 0 2176 0 1 2064
box 0 0 6 6
use CELL  84
transform -1 0 2708 0 1 2124
box 0 0 6 6
use CELL  85
transform -1 0 2611 0 1 2124
box 0 0 6 6
use CELL  86
transform 1 0 2446 0 -1 2094
box 0 0 6 6
use CELL  87
transform -1 0 2503 0 1 2172
box 0 0 6 6
use CELL  88
transform 1 0 2264 0 1 2040
box 0 0 6 6
use CELL  89
transform -1 0 2106 0 1 2244
box 0 0 6 6
use CELL  90
transform -1 0 2131 0 1 2268
box 0 0 6 6
use CELL  91
transform -1 0 2554 0 -1 2286
box 0 0 6 6
use CELL  92
transform 1 0 2721 0 1 2232
box 0 0 6 6
use CELL  93
transform -1 0 2598 0 1 2232
box 0 0 6 6
use CELL  94
transform -1 0 2657 0 1 2244
box 0 0 6 6
use CELL  95
transform -1 0 2502 0 1 2292
box 0 0 6 6
use CELL  96
transform -1 0 2619 0 -1 2118
box 0 0 6 6
use CELL  97
transform -1 0 2099 0 1 2124
box 0 0 6 6
use CELL  98
transform -1 0 2521 0 1 2172
box 0 0 6 6
use CELL  99
transform 1 0 2250 0 1 2040
box 0 0 6 6
use CELL  100
transform 1 0 2257 0 1 2040
box 0 0 6 6
use CELL  101
transform -1 0 2507 0 1 2280
box 0 0 6 6
use CELL  102
transform -1 0 2155 0 1 2304
box 0 0 6 6
use CELL  103
transform -1 0 2632 0 1 2124
box 0 0 6 6
use CELL  104
transform -1 0 2644 0 1 2112
box 0 0 6 6
use CELL  105
transform 1 0 2213 0 1 2040
box 0 0 6 6
use CELL  106
transform -1 0 2218 0 1 2244
box 0 0 6 6
use CELL  107
transform -1 0 2092 0 -1 2250
box 0 0 6 6
use CELL  108
transform -1 0 2071 0 1 2256
box 0 0 6 6
use CELL  109
transform -1 0 2625 0 1 2124
box 0 0 6 6
use CELL  110
transform -1 0 2270 0 1 2268
box 0 0 6 6
use CELL  111
transform -1 0 2102 0 1 2292
box 0 0 6 6
use CELL  112
transform -1 0 2548 0 1 2184
box 0 0 6 6
use CELL  113
transform 1 0 2106 0 -1 2022
box 0 0 6 6
use CELL  114
transform 1 0 2657 0 1 2196
box 0 0 6 6
use CELL  115
transform -1 0 2178 0 1 2124
box 0 0 6 6
use CELL  116
transform -1 0 2510 0 1 2100
box 0 0 6 6
use CELL  117
transform -1 0 2402 0 1 2076
box 0 0 6 6
use CELL  118
transform -1 0 2509 0 1 2160
box 0 0 6 6
use CELL  119
transform -1 0 2416 0 1 2160
box 0 0 6 6
use CELL  120
transform 1 0 2644 0 -1 2166
box 0 0 6 6
use CELL  121
transform -1 0 2221 0 1 2208
box 0 0 6 6
use CELL  122
transform -1 0 2585 0 1 2160
box 0 0 6 6
use CELL  123
transform -1 0 2668 0 1 2112
box 0 0 6 6
use CELL  124
transform -1 0 2084 0 1 2220
box 0 0 6 6
use CELL  125
transform -1 0 2641 0 1 2160
box 0 0 6 6
use CELL  126
transform 1 0 2734 0 1 2232
box 0 0 6 6
use CELL  127
transform -1 0 2284 0 1 2064
box 0 0 6 6
use CELL  128
transform -1 0 2102 0 1 2304
box 0 0 6 6
use CELL  129
transform -1 0 2080 0 1 2268
box 0 0 6 6
use CELL  130
transform 1 0 2251 0 1 2052
box 0 0 6 6
use CELL  131
transform -1 0 2498 0 1 2100
box 0 0 6 6
use CELL  132
transform -1 0 2657 0 1 2124
box 0 0 6 6
use CELL  133
transform -1 0 2083 0 1 2184
box 0 0 6 6
use CELL  134
transform -1 0 2353 0 1 2076
box 0 0 6 6
use CELL  135
transform -1 0 2173 0 1 2148
box 0 0 6 6
use CELL  136
transform -1 0 2278 0 1 2256
box 0 0 6 6
use CELL  137
transform -1 0 2376 0 1 2304
box 0 0 6 6
use CELL  138
transform -1 0 2240 0 1 2040
box 0 0 6 6
use CELL  139
transform 1 0 2100 0 -1 2334
box 0 0 6 6
use CELL  140
transform 1 0 2669 0 1 2268
box 0 0 6 6
use CELL  141
transform -1 0 2264 0 1 2232
box 0 0 6 6
use CELL  142
transform -1 0 2205 0 1 2220
box 0 0 6 6
use CELL  143
transform -1 0 2394 0 1 2088
box 0 0 6 6
use CELL  144
transform -1 0 2461 0 1 2100
box 0 0 6 6
use CELL  145
transform -1 0 2547 0 1 2196
box 0 0 6 6
use CELL  146
transform -1 0 2103 0 1 2100
box 0 0 6 6
use CELL  147
transform -1 0 2580 0 1 2148
box 0 0 6 6
use CELL  148
transform -1 0 2677 0 1 2196
box 0 0 6 6
use CELL  149
transform -1 0 2346 0 1 2304
box 0 0 6 6
use CELL  150
transform -1 0 2078 0 -1 2166
box 0 0 6 6
use CELL  151
transform -1 0 2155 0 1 2196
box 0 0 6 6
use CELL  152
transform -1 0 2174 0 1 2088
box 0 0 6 6
use CELL  153
transform -1 0 2248 0 1 2052
box 0 0 6 6
use CELL  154
transform -1 0 2299 0 1 2160
box 0 0 6 6
use CELL  155
transform -1 0 2089 0 1 2064
box 0 0 6 6
use CELL  156
transform -1 0 2620 0 1 2100
box 0 0 6 6
use CELL  157
transform -1 0 2632 0 1 2244
box 0 0 6 6
use CELL  158
transform -1 0 2595 0 -1 2286
box 0 0 6 6
use CELL  159
transform -1 0 2094 0 1 2268
box 0 0 6 6
use CELL  160
transform -1 0 2641 0 1 2184
box 0 0 6 6
use CELL  161
transform -1 0 2625 0 1 2184
box 0 0 6 6
use CELL  162
transform -1 0 2287 0 1 2100
box 0 0 6 6
use CELL  163
transform -1 0 2201 0 1 2184
box 0 0 6 6
use CELL  164
transform -1 0 2059 0 1 2160
box 0 0 6 6
use CELL  165
transform -1 0 2126 0 1 2136
box 0 0 6 6
use CELL  166
transform -1 0 2178 0 1 2292
box 0 0 6 6
use CELL  167
transform -1 0 2098 0 1 2112
box 0 0 6 6
use CELL  168
transform 1 0 2261 0 1 2316
box 0 0 6 6
use CELL  169
transform -1 0 2167 0 1 2028
box 0 0 6 6
use CELL  170
transform 1 0 2581 0 -1 2250
box 0 0 6 6
use CELL  171
transform -1 0 2143 0 -1 2250
box 0 0 6 6
use CELL  172
transform -1 0 2153 0 1 2316
box 0 0 6 6
use CELL  173
transform -1 0 2483 0 1 2148
box 0 0 6 6
use CELL  174
transform 1 0 2612 0 1 2184
box 0 0 6 6
use CELL  175
transform 1 0 2133 0 -1 2070
box 0 0 6 6
use CELL  176
transform 1 0 2133 0 -1 2166
box 0 0 6 6
use CELL  177
transform 1 0 2300 0 1 2052
box 0 0 6 6
use CELL  178
transform -1 0 2584 0 1 2136
box 0 0 6 6
use CELL  179
transform -1 0 2584 0 1 2112
box 0 0 6 6
use CELL  180
transform 1 0 2307 0 1 2052
box 0 0 6 6
use CELL  181
transform -1 0 2117 0 1 2280
box 0 0 6 6
use CELL  182
transform -1 0 2568 0 1 2148
box 0 0 6 6
use CELL  183
transform -1 0 2241 0 1 2052
box 0 0 6 6
use CELL  184
transform -1 0 2591 0 1 2112
box 0 0 6 6
use CELL  185
transform -1 0 2644 0 1 2232
box 0 0 6 6
use CELL  186
transform -1 0 2263 0 1 2148
box 0 0 6 6
use CELL  187
transform -1 0 2706 0 1 2232
box 0 0 6 6
use CELL  188
transform -1 0 2133 0 1 2136
box 0 0 6 6
use CELL  189
transform -1 0 2614 0 1 2172
box 0 0 6 6
use CELL  190
transform -1 0 2605 0 -1 2118
box 0 0 6 6
use CELL  191
transform -1 0 2064 0 -1 2238
box 0 0 6 6
use CELL  192
transform -1 0 2046 0 -1 2130
box 0 0 6 6
use CELL  193
transform 1 0 2479 0 1 2088
box 0 0 6 6
use CELL  194
transform -1 0 2720 0 1 2124
box 0 0 6 6
use CELL  195
transform -1 0 2124 0 1 2148
box 0 0 6 6
use CELL  196
transform -1 0 2626 0 1 2112
box 0 0 6 6
use CELL  197
transform -1 0 2558 0 1 2268
box 0 0 6 6
use CELL  198
transform 1 0 2291 0 1 2040
box 0 0 6 6
use CELL  199
transform 1 0 2114 0 1 2160
box 0 0 6 6
use CELL  200
transform -1 0 2085 0 1 2172
box 0 0 6 6
use CELL  201
transform 1 0 2657 0 1 2256
box 0 0 6 6
use CELL  202
transform 1 0 2308 0 -1 2070
box 0 0 6 6
use CELL  203
transform -1 0 2122 0 1 2268
box 0 0 6 6
use CELL  204
transform -1 0 2728 0 -1 2226
box 0 0 6 6
use CELL  205
transform -1 0 2091 0 1 2112
box 0 0 6 6
use CELL  206
transform -1 0 2247 0 1 2088
box 0 0 6 6
use CELL  207
transform -1 0 2092 0 1 2172
box 0 0 6 6
use CELL  208
transform 1 0 2606 0 -1 2118
box 0 0 6 6
use CELL  209
transform -1 0 2070 0 1 2112
box 0 0 6 6
use CELL  210
transform -1 0 2679 0 1 2220
box 0 0 6 6
use CELL  211
transform -1 0 2127 0 1 2160
box 0 0 6 6
use CELL  212
transform -1 0 2614 0 1 2208
box 0 0 6 6
use CELL  213
transform -1 0 2759 0 -1 2130
box 0 0 6 6
use CELL  214
transform -1 0 2298 0 1 2064
box 0 0 6 6
use CELL  215
transform 1 0 2611 0 1 2268
box 0 0 6 6
use CELL  216
transform -1 0 2445 0 1 2088
box 0 0 6 6
use CELL  217
transform -1 0 2064 0 -1 2250
box 0 0 6 6
use CELL  218
transform -1 0 2118 0 1 2040
box 0 0 6 6
use CELL  219
transform -1 0 2656 0 1 2196
box 0 0 6 6
use CELL  220
transform -1 0 2082 0 1 2280
box 0 0 6 6
use CELL  221
transform 1 0 2314 0 1 2052
box 0 0 6 6
use CELL  222
transform -1 0 2568 0 -1 2286
box 0 0 6 6
use CELL  223
transform -1 0 2360 0 1 2076
box 0 0 6 6
use CELL  224
transform -1 0 2171 0 1 2328
box 0 0 6 6
use CELL  225
transform -1 0 2100 0 1 2316
box 0 0 6 6
use CELL  226
transform -1 0 2096 0 1 2280
box 0 0 6 6
use CELL  227
transform -1 0 2648 0 1 2136
box 0 0 6 6
use CELL  228
transform 1 0 2220 0 1 2052
box 0 0 6 6
use CELL  229
transform -1 0 2079 0 1 2076
box 0 0 6 6
use CELL  230
transform -1 0 2272 0 1 2244
box 0 0 6 6
use CELL  231
transform -1 0 2085 0 1 2244
box 0 0 6 6
use CELL  232
transform -1 0 2113 0 1 2244
box 0 0 6 6
use CELL  233
transform -1 0 2074 0 1 2124
box 0 0 6 6
use CELL  234
transform -1 0 2126 0 1 2292
box 0 0 6 6
use CELL  235
transform 1 0 2206 0 1 2040
box 0 0 6 6
use CELL  236
transform -1 0 2228 0 1 2268
box 0 0 6 6
use CELL  237
transform 1 0 2185 0 1 2040
box 0 0 6 6
use CELL  238
transform 1 0 2306 0 -1 2226
box 0 0 6 6
use CELL  239
transform 1 0 2053 0 -1 2154
box 0 0 6 6
use CELL  240
transform 1 0 2188 0 -1 2250
box 0 0 6 6
use CELL  241
transform 1 0 2265 0 -1 2262
box 0 0 6 6
use CELL  242
transform -1 0 2104 0 1 2184
box 0 0 6 6
use CELL  243
transform -1 0 2250 0 1 2184
box 0 0 6 6
use CELL  244
transform 1 0 2622 0 1 2208
box 0 0 6 6
use CELL  245
transform 1 0 2347 0 1 2304
box 0 0 6 6
use CELL  246
transform 1 0 2198 0 1 2076
box 0 0 6 6
use CELL  247
transform 1 0 2128 0 1 2040
box 0 0 6 6
use CELL  248
transform -1 0 2084 0 1 2112
box 0 0 6 6
use CELL  249
transform -1 0 2575 0 1 2244
box 0 0 6 6
use CELL  250
transform -1 0 2148 0 1 2304
box 0 0 6 6
use CELL  251
transform 1 0 2109 0 1 2268
box 0 0 6 6
use CELL  252
transform -1 0 2520 0 -1 2118
box 0 0 6 6
use CELL  253
transform 1 0 2158 0 1 2040
box 0 0 6 6
use CELL  254
transform -1 0 2110 0 1 2148
box 0 0 6 6
use CELL  255
transform -1 0 2553 0 1 2136
box 0 0 6 6
use CELL  256
transform -1 0 2305 0 1 2220
box 0 0 6 6
use CELL  257
transform 1 0 2413 0 -1 2094
box 0 0 6 6
use CELL  258
transform -1 0 2096 0 1 2100
box 0 0 6 6
use CELL  259
transform -1 0 2105 0 1 2088
box 0 0 6 6
use CELL  260
transform -1 0 2144 0 1 2184
box 0 0 6 6
use CELL  261
transform -1 0 2150 0 -1 2334
box 0 0 6 6
use CELL  262
transform -1 0 2126 0 1 2076
box 0 0 6 6
use CELL  263
transform -1 0 2488 0 1 2292
box 0 0 6 6
use CELL  264
transform -1 0 2119 0 1 2052
box 0 0 6 6
use CELL  265
transform -1 0 2192 0 1 2232
box 0 0 6 6
use CELL  266
transform -1 0 2128 0 1 2100
box 0 0 6 6
use CELL  267
transform -1 0 2547 0 1 2124
box 0 0 6 6
use CELL  268
transform -1 0 2567 0 1 2160
box 0 0 6 6
use CELL  269
transform -1 0 2639 0 1 2124
box 0 0 6 6
use CELL  270
transform -1 0 2250 0 1 2112
box 0 0 6 6
use CELL  271
transform -1 0 2241 0 1 2196
box 0 0 6 6
use CELL  272
transform -1 0 2213 0 1 2292
box 0 0 6 6
use CELL  273
transform -1 0 2431 0 -1 2262
box 0 0 6 6
use CELL  274
transform -1 0 2112 0 1 2136
box 0 0 6 6
use CELL  275
transform -1 0 2643 0 1 2148
box 0 0 6 6
use CELL  276
transform 1 0 2220 0 1 2040
box 0 0 6 6
use CELL  277
transform 1 0 2692 0 -1 2262
box 0 0 6 6
use CELL  278
transform -1 0 2114 0 1 2316
box 0 0 6 6
use CELL  279
transform -1 0 2306 0 -1 2178
box 0 0 6 6
use CELL  280
transform 1 0 2133 0 1 2316
box 0 0 6 6
use CELL  281
transform -1 0 2046 0 1 2208
box 0 0 6 6
use CELL  282
transform -1 0 2753 0 1 2124
box 0 0 6 6
use CELL  283
transform -1 0 2105 0 -1 2202
box 0 0 6 6
use CELL  284
transform -1 0 2054 0 1 2184
box 0 0 6 6
use CELL  285
transform -1 0 2696 0 1 2112
box 0 0 6 6
use CELL  286
transform -1 0 2520 0 1 2148
box 0 0 6 6
use CELL  287
transform -1 0 2276 0 1 2232
box 0 0 6 6
use CELL  288
transform -1 0 2321 0 1 2172
box 0 0 6 6
use CELL  289
transform 1 0 2185 0 1 2196
box 0 0 6 6
use CELL  290
transform -1 0 2187 0 1 2112
box 0 0 6 6
use CELL  291
transform 1 0 2293 0 1 2052
box 0 0 6 6
use CELL  292
transform 1 0 2133 0 1 2112
box 0 0 6 6
use CELL  293
transform -1 0 2672 0 1 2220
box 0 0 6 6
use CELL  294
transform -1 0 2248 0 1 2220
box 0 0 6 6
use CELL  295
transform -1 0 2145 0 1 2292
box 0 0 6 6
use CELL  296
transform 1 0 2285 0 -1 2070
box 0 0 6 6
use CELL  297
transform -1 0 2611 0 1 2160
box 0 0 6 6
use CELL  298
transform -1 0 2219 0 1 2172
box 0 0 6 6
use CELL  299
transform -1 0 2076 0 -1 2310
box 0 0 6 6
use CELL  300
transform -1 0 2093 0 1 2256
box 0 0 6 6
use CELL  301
transform 1 0 2062 0 -1 2190
box 0 0 6 6
use CELL  302
transform -1 0 2550 0 1 2148
box 0 0 6 6
use CELL  303
transform -1 0 2495 0 1 2292
box 0 0 6 6
use CELL  304
transform -1 0 2185 0 1 2292
box 0 0 6 6
use CELL  305
transform -1 0 2138 0 1 2232
box 0 0 6 6
use CELL  306
transform -1 0 2449 0 1 2160
box 0 0 6 6
use CELL  307
transform -1 0 2093 0 1 2208
box 0 0 6 6
use CELL  308
transform -1 0 2221 0 1 2268
box 0 0 6 6
use CELL  309
transform -1 0 2654 0 1 2268
box 0 0 6 6
use CELL  310
transform 1 0 2272 0 1 2052
box 0 0 6 6
use CELL  311
transform -1 0 2100 0 1 2256
box 0 0 6 6
use CELL  312
transform -1 0 2078 0 1 2172
box 0 0 6 6
use CELL  313
transform -1 0 2110 0 1 2280
box 0 0 6 6
use CELL  314
transform -1 0 2123 0 1 2208
box 0 0 6 6
use CELL  315
transform 1 0 2655 0 -1 2274
box 0 0 6 6
use CELL  316
transform -1 0 2412 0 1 2088
box 0 0 6 6
use CELL  317
transform -1 0 2595 0 1 2172
box 0 0 6 6
use CELL  318
transform -1 0 2133 0 1 2292
box 0 0 6 6
use CELL  319
transform -1 0 2474 0 1 2292
box 0 0 6 6
use CELL  320
transform -1 0 2432 0 -1 2082
box 0 0 6 6
use CELL  321
transform -1 0 2712 0 1 2256
box 0 0 6 6
use CELL  322
transform -1 0 2136 0 1 2016
box 0 0 6 6
use CELL  323
transform -1 0 2150 0 1 2076
box 0 0 6 6
use CELL  324
transform -1 0 2086 0 -1 2262
box 0 0 6 6
use CELL  325
transform 1 0 2321 0 1 2052
box 0 0 6 6
use CELL  326
transform -1 0 2346 0 1 2076
box 0 0 6 6
use CELL  327
transform -1 0 2376 0 1 2136
box 0 0 6 6
use CELL  328
transform -1 0 2085 0 1 2160
box 0 0 6 6
use CELL  329
transform -1 0 2081 0 -1 2130
box 0 0 6 6
use CELL  330
transform 1 0 2639 0 -1 2262
box 0 0 6 6
use CELL  331
transform 1 0 2453 0 1 2088
box 0 0 6 6
use CELL  332
transform -1 0 2358 0 1 2088
box 0 0 6 6
use CELL  333
transform -1 0 2086 0 1 2076
box 0 0 6 6
use CELL  334
transform -1 0 2447 0 1 2292
box 0 0 6 6
use CELL  335
transform -1 0 2546 0 1 2220
box 0 0 6 6
use CELL  336
transform 1 0 2669 0 -1 2118
box 0 0 6 6
use CELL  337
transform -1 0 2107 0 1 2316
box 0 0 6 6
use CELL  338
transform -1 0 2242 0 1 2208
box 0 0 6 6
use CELL  339
transform 1 0 2595 0 1 2148
box 0 0 6 6
use CELL  340
transform -1 0 2560 0 1 2136
box 0 0 6 6
use CELL  341
transform -1 0 2513 0 1 2148
box 0 0 6 6
use CELL  342
transform 1 0 2059 0 -1 2202
box 0 0 6 6
use CELL  343
transform -1 0 2114 0 1 2256
box 0 0 6 6
use CELL  344
transform -1 0 2641 0 1 2136
box 0 0 6 6
use CELL  345
transform -1 0 2631 0 1 2256
box 0 0 6 6
use CELL  346
transform 1 0 2531 0 -1 2166
box 0 0 6 6
use CELL  347
transform -1 0 2635 0 1 2208
box 0 0 6 6
use CELL  348
transform -1 0 2523 0 1 2136
box 0 0 6 6
use CELL  349
transform -1 0 2662 0 1 2136
box 0 0 6 6
use CELL  350
transform -1 0 2590 0 1 2100
box 0 0 6 6
use CELL  351
transform -1 0 2142 0 1 2136
box 0 0 6 6
use CELL  352
transform -1 0 2574 0 1 2172
box 0 0 6 6
use CELL  353
transform 1 0 2284 0 1 2148
box 0 0 6 6
use CELL  354
transform -1 0 2565 0 1 2112
box 0 0 6 6
use CELL  355
transform 1 0 2158 0 1 2064
box 0 0 6 6
use CELL  356
transform -1 0 2072 0 1 2136
box 0 0 6 6
use CELL  357
transform 1 0 2061 0 -1 2130
box 0 0 6 6
use CELL  358
transform -1 0 2705 0 1 2256
box 0 0 6 6
use CELL  359
transform -1 0 2181 0 1 2280
box 0 0 6 6
use CELL  360
transform -1 0 2089 0 1 2100
box 0 0 6 6
use CELL  361
transform -1 0 2369 0 1 2076
box 0 0 6 6
use CELL  362
transform -1 0 2582 0 -1 2286
box 0 0 6 6
use CELL  363
transform -1 0 2082 0 1 2100
box 0 0 6 6
use CELL  364
transform -1 0 2511 0 1 2184
box 0 0 6 6
use CELL  365
transform -1 0 2668 0 1 2268
box 0 0 6 6
use CELL  366
transform -1 0 2084 0 1 2136
box 0 0 6 6
use CELL  367
transform -1 0 2657 0 1 2160
box 0 0 6 6
use CELL  368
transform -1 0 2098 0 1 2088
box 0 0 6 6
use CELL  369
transform -1 0 2480 0 1 2100
box 0 0 6 6
use CELL  370
transform 1 0 2140 0 -1 2322
box 0 0 6 6
use CELL  371
transform -1 0 2052 0 1 2112
box 0 0 6 6
use CELL  372
transform -1 0 2507 0 1 2088
box 0 0 6 6
use CELL  373
transform -1 0 2052 0 1 2160
box 0 0 6 6
use CELL  374
transform 1 0 2551 0 -1 2106
box 0 0 6 6
use CELL  375
transform -1 0 2121 0 1 2220
box 0 0 6 6
use CELL  376
transform -1 0 2238 0 1 2136
box 0 0 6 6
use CELL  377
transform -1 0 2465 0 1 2280
box 0 0 6 6
use CELL  378
transform -1 0 2343 0 1 2124
box 0 0 6 6
use CELL  379
transform -1 0 2236 0 1 2316
box 0 0 6 6
use CELL  380
transform -1 0 2089 0 1 2280
box 0 0 6 6
use CELL  381
transform 1 0 2243 0 1 2040
box 0 0 6 6
use CELL  382
transform -1 0 2101 0 1 2052
box 0 0 6 6
use CELL  383
transform -1 0 2481 0 1 2292
box 0 0 6 6
use CELL  384
transform 1 0 2645 0 1 2232
box 0 0 6 6
use CELL  385
transform -1 0 2103 0 1 2280
box 0 0 6 6
use CELL  386
transform -1 0 2365 0 1 2208
box 0 0 6 6
use CELL  387
transform -1 0 2575 0 1 2280
box 0 0 6 6
use CELL  388
transform -1 0 2077 0 1 2196
box 0 0 6 6
use CELL  389
transform -1 0 2369 0 1 2304
box 0 0 6 6
use CELL  390
transform -1 0 2071 0 1 2232
box 0 0 6 6
use CELL  391
transform -1 0 2600 0 1 2196
box 0 0 6 6
use CELL  392
transform 1 0 2103 0 1 2304
box 0 0 6 6
use CELL  393
transform -1 0 2285 0 1 2052
box 0 0 6 6
use CELL  394
transform 1 0 2583 0 -1 2286
box 0 0 6 6
use CELL  395
transform -1 0 2485 0 1 2160
box 0 0 6 6
use CELL  396
transform -1 0 2531 0 1 2100
box 0 0 6 6
use CELL  397
transform -1 0 2420 0 -1 2298
box 0 0 6 6
use CELL  398
transform -1 0 2119 0 1 2076
box 0 0 6 6
use CELL  399
transform -1 0 2458 0 1 2280
box 0 0 6 6
use CELL  400
transform -1 0 2496 0 1 2136
box 0 0 6 6
use CELL  401
transform -1 0 2087 0 1 2148
box 0 0 6 6
use CELL  402
transform 1 0 2611 0 1 2136
box 0 0 6 6
use CELL  403
transform -1 0 2105 0 1 2136
box 0 0 6 6
use CELL  404
transform -1 0 2367 0 -1 2070
box 0 0 6 6
use CELL  405
transform -1 0 2082 0 1 2064
box 0 0 6 6
use CELL  406
transform -1 0 2110 0 1 2100
box 0 0 6 6
use CELL  407
transform -1 0 2047 0 1 2184
box 0 0 6 6
use CELL  408
transform -1 0 2070 0 1 2100
box 0 0 6 6
use CELL  409
transform -1 0 2716 0 1 2112
box 0 0 6 6
use CELL  410
transform 1 0 2104 0 1 2052
box 0 0 6 6
use CELL  411
transform 1 0 2094 0 1 2028
box 0 0 6 6
use CELL  412
transform 1 0 2683 0 1 2268
box 0 0 6 6
use CELL  413
transform -1 0 2560 0 1 2184
box 0 0 6 6
use CELL  414
transform 1 0 2172 0 1 2328
box 0 0 6 6
use CELL  415
transform -1 0 2212 0 1 2220
box 0 0 6 6
use CELL  416
transform -1 0 2519 0 1 2100
box 0 0 6 6
use CELL  417
transform -1 0 2166 0 1 2292
box 0 0 6 6
use CELL  418
transform -1 0 2171 0 1 2184
box 0 0 6 6
use CELL  419
transform 1 0 2082 0 -1 2034
box 0 0 6 6
use CELL  420
transform -1 0 2339 0 1 2064
box 0 0 6 6
use CELL  421
transform -1 0 2584 0 1 2124
box 0 0 6 6
use CELL  422
transform -1 0 2451 0 1 2280
box 0 0 6 6
use CELL  423
transform 1 0 2721 0 1 2124
box 0 0 6 6
use CELL  424
transform 1 0 2034 0 -1 2190
box 0 0 6 6
use CELL  425
transform -1 0 2734 0 1 2124
box 0 0 6 6
use CELL  426
transform -1 0 2093 0 -1 2226
box 0 0 6 6
use CELL  427
transform -1 0 2101 0 1 2268
box 0 0 6 6
use CELL  428
transform -1 0 2471 0 1 2088
box 0 0 6 6
use CELL  429
transform 1 0 2047 0 1 2208
box 0 0 6 6
use CELL  430
transform -1 0 2332 0 1 2256
box 0 0 6 6
use CELL  431
transform -1 0 2602 0 1 2244
box 0 0 6 6
use CELL  432
transform -1 0 2408 0 1 2292
box 0 0 6 6
use CELL  433
transform -1 0 2671 0 1 2124
box 0 0 6 6
use CELL  434
transform -1 0 2227 0 1 2160
box 0 0 6 6
use CELL  435
transform -1 0 2554 0 1 2124
box 0 0 6 6
use CELL  436
transform -1 0 2108 0 1 2268
box 0 0 6 6
use CELL  437
transform -1 0 2119 0 1 2136
box 0 0 6 6
use CELL  438
transform -1 0 2091 0 1 2196
box 0 0 6 6
use CELL  439
transform 1 0 2671 0 1 2208
box 0 0 6 6
use CELL  440
transform -1 0 2091 0 1 2136
box 0 0 6 6
use CELL  441
transform 1 0 2120 0 1 2052
box 0 0 6 6
use CELL  442
transform 1 0 2131 0 -1 2034
box 0 0 6 6
use CELL  443
transform 1 0 2298 0 -1 2082
box 0 0 6 6
use CELL  444
transform -1 0 2388 0 1 2304
box 0 0 6 6
use CELL  445
transform -1 0 2160 0 -1 2322
box 0 0 6 6
use CELL  446
transform -1 0 2130 0 1 2112
box 0 0 6 6
use CELL  447
transform -1 0 2605 0 1 2208
box 0 0 6 6
use CELL  448
transform -1 0 2164 0 1 2328
box 0 0 6 6
use CELL  449
transform 1 0 2340 0 -1 2070
box 0 0 6 6
use CELL  450
transform 1 0 2139 0 -1 2130
box 0 0 6 6
use CELL  451
transform -1 0 2323 0 1 2064
box 0 0 6 6
use CELL  452
transform 1 0 2220 0 1 2028
box 0 0 6 6
use CELL  453
transform -1 0 2099 0 1 2244
box 0 0 6 6
use CELL  454
transform -1 0 2536 0 1 2208
box 0 0 6 6
use CELL  455
transform 1 0 2258 0 1 2052
box 0 0 6 6
use CELL  456
transform 1 0 2177 0 -1 2178
box 0 0 6 6
use CELL  457
transform -1 0 2092 0 1 2160
box 0 0 6 6
use CELL  458
transform -1 0 2125 0 1 2184
box 0 0 6 6
use CELL  459
transform -1 0 2172 0 1 2256
box 0 0 6 6
use CELL  460
transform 1 0 2340 0 1 2136
box 0 0 6 6
use CELL  461
transform -1 0 2186 0 1 2304
box 0 0 6 6
use CELL  462
transform -1 0 2127 0 1 2124
box 0 0 6 6
use CELL  463
transform -1 0 2550 0 1 2100
box 0 0 6 6
use CELL  464
transform -1 0 2718 0 1 2244
box 0 0 6 6
use CELL  465
transform -1 0 2094 0 1 2052
box 0 0 6 6
use CELL  466
transform -1 0 2061 0 1 2184
box 0 0 6 6
use CELL  467
transform -1 0 2666 0 1 2148
box 0 0 6 6
use CELL  468
transform -1 0 2514 0 1 2280
box 0 0 6 6
use CELL  469
transform 1 0 2140 0 1 2028
box 0 0 6 6
use CELL  470
transform 1 0 2146 0 1 2040
box 0 0 6 6
use CELL  471
transform -1 0 2123 0 1 2316
box 0 0 6 6
use CELL  472
transform 1 0 2522 0 -1 2178
box 0 0 6 6
use CELL  473
transform -1 0 2114 0 1 2220
box 0 0 6 6
use CELL  474
transform 1 0 2208 0 1 2052
box 0 0 6 6
use CELL  475
transform -1 0 2607 0 1 2196
box 0 0 6 6
use CELL  476
transform -1 0 2528 0 1 2088
box 0 0 6 6
use CELL  477
transform -1 0 2073 0 1 2268
box 0 0 6 6
use CELL  478
transform -1 0 2090 0 1 2184
box 0 0 6 6
use CELL  479
transform -1 0 2572 0 1 2100
box 0 0 6 6
use CELL  480
transform 1 0 2672 0 -1 2130
box 0 0 6 6
use CELL  481
transform -1 0 2107 0 1 2256
box 0 0 6 6
use CELL  482
transform -1 0 2605 0 1 2232
box 0 0 6 6
use CELL  483
transform -1 0 2072 0 1 2220
box 0 0 6 6
use CELL  484
transform -1 0 2106 0 1 2124
box 0 0 6 6
use CELL  485
transform -1 0 2364 0 1 2184
box 0 0 6 6
use CELL  486
transform -1 0 2602 0 1 2280
box 0 0 6 6
use CELL  487
transform -1 0 2565 0 1 2268
box 0 0 6 6
use CELL  488
transform -1 0 2116 0 1 2208
box 0 0 6 6
use CELL  489
transform -1 0 2084 0 1 2088
box 0 0 6 6
use CELL  490
transform -1 0 2130 0 1 2316
box 0 0 6 6
use CELL  491
transform -1 0 2605 0 1 2136
box 0 0 6 6
use CELL  492
transform -1 0 2133 0 1 2256
box 0 0 6 6
use CELL  493
transform -1 0 2663 0 1 2232
box 0 0 6 6
use CELL  494
transform -1 0 2192 0 1 2076
box 0 0 6 6
use CELL  495
transform -1 0 2307 0 1 2064
box 0 0 6 6
use CELL  496
transform 1 0 2715 0 1 2220
box 0 0 6 6
use CELL  497
transform 1 0 2389 0 -1 2310
box 0 0 6 6
use CELL  498
transform -1 0 2591 0 1 2232
box 0 0 6 6
use CELL  499
transform 1 0 2118 0 -1 2286
box 0 0 6 6
use CELL  500
transform -1 0 2088 0 1 2292
box 0 0 6 6
use CELL  501
transform -1 0 2235 0 1 2208
box 0 0 6 6
use CELL  502
transform -1 0 2330 0 1 2292
box 0 0 6 6
use CELL  503
transform -1 0 2709 0 1 2220
box 0 0 6 6
use CELL  504
transform -1 0 2592 0 1 2160
box 0 0 6 6
use CELL  505
transform -1 0 2093 0 1 2232
box 0 0 6 6
use CELL  506
transform -1 0 2162 0 1 2232
box 0 0 6 6
use CELL  507
transform 1 0 2760 0 1 2124
box 0 0 6 6
use CELL  508
transform -1 0 2439 0 1 2172
box 0 0 6 6
use CELL  509
transform -1 0 2066 0 1 2148
box 0 0 6 6
use CELL  510
transform -1 0 2283 0 1 2316
box 0 0 6 6
use CELL  511
transform 1 0 2703 0 1 2244
box 0 0 6 6
use CELL  512
transform -1 0 2611 0 1 2100
box 0 0 6 6
use CELL  513
transform -1 0 2664 0 1 2244
box 0 0 6 6
use CELL  514
transform -1 0 2241 0 1 2280
box 0 0 6 6
use CELL  515
transform -1 0 2145 0 1 2220
box 0 0 6 6
use CELL  516
transform -1 0 2344 0 1 2160
box 0 0 6 6
use CELL  517
transform 1 0 2198 0 -1 2034
box 0 0 6 6
use CELL  518
transform -1 0 2709 0 1 2268
box 0 0 6 6
use CELL  519
transform -1 0 2289 0 1 2088
box 0 0 6 6
use CELL  520
transform 1 0 2040 0 -1 2142
box 0 0 6 6
use CELL  521
transform -1 0 2593 0 1 2184
box 0 0 6 6
use CELL  522
transform -1 0 2360 0 1 2064
box 0 0 6 6
use CELL  523
transform -1 0 2114 0 1 2064
box 0 0 6 6
use CELL  524
transform -1 0 2129 0 1 2328
box 0 0 6 6
use CELL  525
transform 1 0 2059 0 1 2136
box 0 0 6 6
use CELL  526
transform -1 0 2183 0 1 2064
box 0 0 6 6
use CELL  527
transform -1 0 2607 0 1 2172
box 0 0 6 6
use CELL  528
transform -1 0 2587 0 1 2148
box 0 0 6 6
use CELL  529
transform -1 0 2369 0 1 2172
box 0 0 6 6
use CELL  530
transform 1 0 2074 0 -1 2154
box 0 0 6 6
use CELL  531
transform -1 0 2530 0 1 2160
box 0 0 6 6
use CELL  532
transform -1 0 2618 0 1 2124
box 0 0 6 6
use CELL  533
transform -1 0 2272 0 1 2064
box 0 0 6 6
use CELL  534
transform -1 0 2114 0 1 2232
box 0 0 6 6
use CELL  535
transform -1 0 2597 0 1 2100
box 0 0 6 6
use CELL  536
transform -1 0 2567 0 1 2172
box 0 0 6 6
use CELL  537
transform -1 0 2107 0 1 2232
box 0 0 6 6
use CELL  538
transform -1 0 2137 0 1 2196
box 0 0 6 6
use CELL  539
transform -1 0 2122 0 1 2328
box 0 0 6 6
use CELL  540
transform -1 0 2243 0 1 2316
box 0 0 6 6
use CELL  541
transform -1 0 2185 0 1 2328
box 0 0 6 6
use CELL  542
transform -1 0 2190 0 1 2256
box 0 0 6 6
use CELL  543
transform -1 0 2282 0 1 2268
box 0 0 6 6
use CELL  544
transform -1 0 2203 0 1 2100
box 0 0 6 6
use CELL  545
transform -1 0 2367 0 1 2124
box 0 0 6 6
use CELL  546
transform -1 0 2175 0 1 2052
box 0 0 6 6
use CELL  547
transform -1 0 2216 0 1 2196
box 0 0 6 6
use CELL  548
transform -1 0 2086 0 1 2208
box 0 0 6 6
use CELL  549
transform -1 0 2064 0 1 2268
box 0 0 6 6
use CELL  550
transform 1 0 2191 0 1 2028
box 0 0 6 6
use CELL  551
transform 1 0 2644 0 1 2148
box 0 0 6 6
use CELL  552
transform -1 0 2687 0 1 2232
box 0 0 6 6
use CELL  553
transform -1 0 2290 0 1 2316
box 0 0 6 6
use CELL  554
transform 1 0 2265 0 1 2052
box 0 0 6 6
use CELL  555
transform -1 0 2432 0 1 2172
box 0 0 6 6
use CELL  556
transform -1 0 2297 0 1 2076
box 0 0 6 6
use CELL  557
transform -1 0 2167 0 1 2208
box 0 0 6 6
use CELL  558
transform 1 0 2676 0 1 2268
box 0 0 6 6
use CELL  559
transform 1 0 2566 0 1 2184
box 0 0 6 6
use CELL  560
transform 1 0 2623 0 -1 2274
box 0 0 6 6
use CELL  561
transform -1 0 2554 0 1 2208
box 0 0 6 6
use CELL  562
transform -1 0 2058 0 1 2196
box 0 0 6 6
use CELL  563
transform -1 0 2720 0 1 2232
box 0 0 6 6
use CELL  564
transform -1 0 2052 0 1 2148
box 0 0 6 6
use CELL  565
transform 1 0 2117 0 -1 2034
box 0 0 6 6
use CELL  566
transform -1 0 2699 0 -1 2238
box 0 0 6 6
use CELL  567
transform -1 0 2613 0 1 2220
box 0 0 6 6
use CELL  568
transform -1 0 2118 0 -1 2346
box 0 0 6 6
use CELL  569
transform -1 0 2060 0 1 2208
box 0 0 6 6
use CELL  570
transform -1 0 2113 0 1 2160
box 0 0 6 6
use CELL  571
transform -1 0 2294 0 1 2232
box 0 0 6 6
use CELL  572
transform -1 0 2526 0 1 2196
box 0 0 6 6
use CELL  573
transform 1 0 2729 0 -1 2226
box 0 0 6 6
use CELL  574
transform 1 0 2678 0 1 2112
box 0 0 6 6
use CELL  575
transform -1 0 2334 0 1 2076
box 0 0 6 6
use CELL  576
transform 1 0 2324 0 1 2064
box 0 0 6 6
use CELL  577
transform -1 0 2094 0 -1 2154
box 0 0 6 6
use CELL  578
transform -1 0 2594 0 1 2256
box 0 0 6 6
use CELL  579
transform -1 0 2274 0 1 2316
box 0 0 6 6
use CELL  580
transform 1 0 2529 0 -1 2202
box 0 0 6 6
use CELL  581
transform 1 0 2419 0 1 2076
box 0 0 6 6
use CELL  582
transform -1 0 2076 0 1 2244
box 0 0 6 6
use CELL  583
transform -1 0 2160 0 1 2280
box 0 0 6 6
use CELL  584
transform 1 0 2540 0 1 2268
box 0 0 6 6
use CELL  585
transform -1 0 2424 0 1 2136
box 0 0 6 6
use CELL  586
transform -1 0 2058 0 1 2136
box 0 0 6 6
use CELL  587
transform 1 0 2494 0 1 2088
box 0 0 6 6
use CELL  588
transform 1 0 2531 0 1 2172
box 0 0 6 6
use CELL  589
transform 1 0 2371 0 1 2148
box 0 0 6 6
use CELL  590
transform -1 0 2203 0 1 2040
box 0 0 6 6
use CELL  591
transform 1 0 2100 0 1 2040
box 0 0 6 6
use CELL  592
transform -1 0 2376 0 1 2076
box 0 0 6 6
use CELL  593
transform -1 0 2064 0 1 2256
box 0 0 6 6
use CELL  594
transform 1 0 2685 0 -1 2214
box 0 0 6 6
use CELL  595
transform -1 0 2664 0 1 2160
box 0 0 6 6
use CELL  596
transform -1 0 2554 0 1 2196
box 0 0 6 6
use CELL  597
transform -1 0 2307 0 1 2136
box 0 0 6 6
use CELL  598
transform -1 0 2102 0 1 2208
box 0 0 6 6
use CELL  599
transform -1 0 2703 0 1 2112
box 0 0 6 6
use CELL  600
transform -1 0 2674 0 -1 2142
box 0 0 6 6
use CELL  601
transform -1 0 2160 0 1 2208
box 0 0 6 6
use CELL  602
transform -1 0 2228 0 1 2208
box 0 0 6 6
use CELL  603
transform -1 0 2487 0 1 2112
box 0 0 6 6
use CELL  604
transform 1 0 2286 0 1 2052
box 0 0 6 6
use CELL  605
transform -1 0 2118 0 1 2184
box 0 0 6 6
use CELL  606
transform -1 0 2262 0 1 2184
box 0 0 6 6
use CELL  607
transform -1 0 2702 0 1 2244
box 0 0 6 6
use CELL  608
transform -1 0 2632 0 1 2184
box 0 0 6 6
use CELL  609
transform -1 0 2157 0 1 2064
box 0 0 6 6
use CELL  610
transform -1 0 2174 0 1 2028
box 0 0 6 6
use CELL  611
transform 1 0 2684 0 1 2124
box 0 0 6 6
use CELL  612
transform -1 0 2635 0 1 2172
box 0 0 6 6
use CELL  613
transform -1 0 2594 0 1 2220
box 0 0 6 6
use CELL  614
transform 1 0 2618 0 -1 2262
box 0 0 6 6
use CELL  615
transform 1 0 2651 0 1 2148
box 0 0 6 6
use CELL  616
transform 1 0 2563 0 -1 2262
box 0 0 6 6
use CELL  617
transform -1 0 2231 0 1 2184
box 0 0 6 6
use CELL  618
transform -1 0 2105 0 1 2112
box 0 0 6 6
use CELL  619
transform -1 0 2473 0 1 2100
box 0 0 6 6
use CELL  620
transform 1 0 2227 0 1 2040
box 0 0 6 6
use CELL  621
transform -1 0 2655 0 1 2136
box 0 0 6 6
use CELL  622
transform 1 0 2704 0 1 2112
box 0 0 6 6
use CELL  623
transform -1 0 2180 0 1 2076
box 0 0 6 6
use CELL  624
transform -1 0 2438 0 1 2088
box 0 0 6 6
use CELL  625
transform -1 0 2109 0 1 2208
box 0 0 6 6
use CELL  626
transform -1 0 2244 0 1 2064
box 0 0 6 6
use CELL  627
transform -1 0 2084 0 1 2196
box 0 0 6 6
use CELL  628
transform -1 0 2621 0 1 2208
box 0 0 6 6
use CELL  629
transform 1 0 2137 0 1 2040
box 0 0 6 6
use CELL  630
transform -1 0 2572 0 1 2112
box 0 0 6 6
use CELL  631
transform -1 0 2133 0 1 2220
box 0 0 6 6
use CELL  632
transform -1 0 2395 0 1 2076
box 0 0 6 6
use CELL  633
transform -1 0 2130 0 1 2304
box 0 0 6 6
use CELL  634
transform -1 0 2088 0 1 2304
box 0 0 6 6
use CELL  635
transform 1 0 2621 0 1 2100
box 0 0 6 6
use CELL  636
transform -1 0 2210 0 1 2028
box 0 0 6 6
use CELL  637
transform -1 0 2530 0 1 2184
box 0 0 6 6
use CELL  638
transform -1 0 2234 0 1 2196
box 0 0 6 6
use CELL  639
transform -1 0 2095 0 1 2292
box 0 0 6 6
use CELL  640
transform -1 0 2111 0 1 2184
box 0 0 6 6
use CELL  641
transform -1 0 2097 0 1 2184
box 0 0 6 6
use CELL  642
transform -1 0 2576 0 1 2256
box 0 0 6 6
use CELL  643
transform -1 0 2604 0 1 2100
box 0 0 6 6
use CELL  644
transform -1 0 2147 0 1 2052
box 0 0 6 6
use CELL  645
transform -1 0 2098 0 1 2064
box 0 0 6 6
use CELL  646
transform -1 0 2634 0 1 2100
box 0 0 6 6
use CELL  647
transform -1 0 2120 0 1 2124
box 0 0 6 6
use CELL  648
transform -1 0 2394 0 1 2196
box 0 0 6 6
use CELL  649
transform -1 0 2628 0 1 2172
box 0 0 6 6
use CELL  650
transform -1 0 2101 0 1 2148
box 0 0 6 6
use CELL  651
transform -1 0 2211 0 1 2280
box 0 0 6 6
use CELL  652
transform 1 0 2068 0 1 2208
box 0 0 6 6
use CELL  653
transform -1 0 2117 0 1 2148
box 0 0 6 6
use CELL  654
transform -1 0 2718 0 1 2256
box 0 0 6 6
use CELL  655
transform -1 0 2416 0 -1 2082
box 0 0 6 6
use CELL  656
transform -1 0 2561 0 1 2280
box 0 0 6 6
use CELL  657
transform -1 0 2104 0 1 2160
box 0 0 6 6
use CELL  658
transform -1 0 2555 0 1 2172
box 0 0 6 6
use CELL  659
transform -1 0 2113 0 1 2124
box 0 0 6 6
use CELL  660
transform 1 0 2626 0 -1 2238
box 0 0 6 6
use CELL  661
transform -1 0 2176 0 1 2268
box 0 0 6 6
use CELL  662
transform -1 0 2136 0 1 2328
box 0 0 6 6
use CELL  663
transform 1 0 2148 0 1 2052
box 0 0 6 6
use CELL  664
transform -1 0 2141 0 1 2208
box 0 0 6 6
use CELL  665
transform -1 0 2461 0 1 2172
box 0 0 6 6
use CELL  666
transform -1 0 2136 0 1 2148
box 0 0 6 6
use CELL  667
transform 1 0 2186 0 -1 2334
box 0 0 6 6
use CELL  668
transform -1 0 2160 0 1 2028
box 0 0 6 6
use CELL  669
transform -1 0 2116 0 1 2028
box 0 0 6 6
use CELL  670
transform -1 0 2123 0 1 2304
box 0 0 6 6
use CELL  671
transform -1 0 2221 0 -1 2106
box 0 0 6 6
use CELL  672
transform -1 0 2259 0 1 2136
box 0 0 6 6
use CELL  673
transform -1 0 2294 0 1 2304
box 0 0 6 6
use CELL  674
transform -1 0 2664 0 1 2124
box 0 0 6 6
use CELL  675
transform -1 0 2591 0 1 2136
box 0 0 6 6
use CELL  676
transform -1 0 2070 0 1 2076
box 0 0 6 6
use CELL  677
transform -1 0 2335 0 1 2148
box 0 0 6 6
use CELL  678
transform -1 0 2126 0 1 2232
box 0 0 6 6
use CELL  679
transform -1 0 2091 0 1 2088
box 0 0 6 6
use CELL  680
transform -1 0 2746 0 1 2124
box 0 0 6 6
use CELL  681
transform -1 0 2229 0 1 2316
box 0 0 6 6
use CELL  682
transform -1 0 2105 0 1 2064
box 0 0 6 6
use CELL  683
transform -1 0 2670 0 -1 2262
box 0 0 6 6
use CELL  684
transform -1 0 2155 0 1 2100
box 0 0 6 6
use CELL  685
transform -1 0 2112 0 1 2112
box 0 0 6 6
use CELL  686
transform -1 0 2529 0 -1 2286
box 0 0 6 6
use CELL  687
transform -1 0 2067 0 1 2208
box 0 0 6 6
use CELL  688
transform 1 0 2696 0 1 2268
box 0 0 6 6
use CELL  689
transform 1 0 2605 0 -1 2190
box 0 0 6 6
use CELL  690
transform -1 0 2301 0 1 2304
box 0 0 6 6
use CELL  691
transform -1 0 2287 0 1 2244
box 0 0 6 6
use CELL  692
transform -1 0 2431 0 1 2088
box 0 0 6 6
use CELL  693
transform -1 0 2125 0 1 2040
box 0 0 6 6
use CELL  694
transform -1 0 2238 0 1 2184
box 0 0 6 6
use CELL  695
transform 1 0 2137 0 1 2148
box 0 0 6 6
use CELL  696
transform -1 0 2478 0 1 2088
box 0 0 6 6
use CELL  697
transform -1 0 2265 0 1 2064
box 0 0 6 6
use CELL  698
transform -1 0 2538 0 1 2100
box 0 0 6 6
use CELL  699
transform -1 0 2621 0 1 2172
box 0 0 6 6
use CELL  700
transform -1 0 2131 0 1 2244
box 0 0 6 6
use CELL  701
transform 1 0 2652 0 -1 2226
box 0 0 6 6
use CELL  702
transform -1 0 2695 0 1 2244
box 0 0 6 6
use CELL  703
transform -1 0 2163 0 1 2220
box 0 0 6 6
use CELL  704
transform -1 0 2547 0 1 2280
box 0 0 6 6
use CELL  705
transform -1 0 2114 0 1 2172
box 0 0 6 6
use CELL  706
transform -1 0 2162 0 1 2304
box 0 0 6 6
use CELL  707
transform -1 0 2087 0 1 2268
box 0 0 6 6
use CELL  708
transform -1 0 2119 0 1 2196
box 0 0 6 6
use CELL  709
transform -1 0 2146 0 1 2160
box 0 0 6 6
use CELL  710
transform -1 0 2204 0 1 2232
box 0 0 6 6
use CELL  711
transform -1 0 2443 0 1 2208
box 0 0 6 6
use CELL  712
transform -1 0 2594 0 1 2148
box 0 0 6 6
use CELL  713
transform -1 0 2382 0 1 2088
box 0 0 6 6
use CELL  714
transform -1 0 2684 0 1 2208
box 0 0 6 6
use CELL  715
transform -1 0 2670 0 -1 2202
box 0 0 6 6
use CELL  716
transform -1 0 2053 0 1 2124
box 0 0 6 6
use CELL  717
transform 1 0 2285 0 1 2040
box 0 0 6 6
use CELL  718
transform -1 0 2604 0 1 2160
box 0 0 6 6
use CELL  719
transform -1 0 2677 0 1 2256
box 0 0 6 6
use CELL  720
transform 1 0 2187 0 1 2088
box 0 0 6 6
use FEEDTHRU  F-1
transform 1 0 2361 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-2
transform 1 0 2464 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-3
transform 1 0 2523 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-4
transform 1 0 2125 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-5
transform 1 0 2132 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-6
transform 1 0 2170 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-7
transform 1 0 2259 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-8
transform 1 0 2632 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-9
transform 1 0 2632 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-10
transform 1 0 2640 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-11
transform 1 0 2581 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-12
transform 1 0 2581 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-13
transform 1 0 2536 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-14
transform 1 0 2543 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-15
transform 1 0 2617 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-16
transform 1 0 2517 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-17
transform 1 0 2447 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-18
transform 1 0 2629 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-19
transform 1 0 2708 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-20
transform 1 0 2656 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-21
transform 1 0 2321 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-22
transform 1 0 2388 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-23
transform 1 0 2537 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-24
transform 1 0 2554 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-25
transform 1 0 2578 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-26
transform 1 0 2582 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-27
transform 1 0 2309 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-28
transform 1 0 2391 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-29
transform 1 0 2531 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-30
transform 1 0 2545 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-31
transform 1 0 2308 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-32
transform 1 0 2255 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-33
transform 1 0 2259 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-34
transform 1 0 2324 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-35
transform 1 0 2524 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-36
transform 1 0 2125 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-37
transform 1 0 2269 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-38
transform 1 0 2239 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-39
transform 1 0 2231 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-40
transform 1 0 2233 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-41
transform 1 0 2448 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-42
transform 1 0 2575 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-43
transform 1 0 2268 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-44
transform 1 0 2173 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-45
transform 1 0 2135 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-46
transform 1 0 2204 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-47
transform 1 0 2065 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-48
transform 1 0 2311 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-49
transform 1 0 2333 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-50
transform 1 0 2339 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-51
transform 1 0 2326 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-52
transform 1 0 2299 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-53
transform 1 0 2166 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-54
transform 1 0 2169 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-55
transform 1 0 2308 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-56
transform 1 0 2256 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-57
transform 1 0 2278 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-58
transform 1 0 2322 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-59
transform 1 0 2358 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-60
transform 1 0 2584 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-61
transform 1 0 2643 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-62
transform 1 0 2635 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-63
transform 1 0 2635 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-64
transform 1 0 2615 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-65
transform 1 0 2620 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-66
transform 1 0 2520 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-67
transform 1 0 2575 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-68
transform 1 0 2539 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-69
transform 1 0 2546 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-70
transform 1 0 2567 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-71
transform 1 0 2550 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-72
transform 1 0 2566 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-73
transform 1 0 2657 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-74
transform 1 0 2676 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-75
transform 1 0 2687 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-76
transform 1 0 2709 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-77
transform 1 0 2665 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-78
transform 1 0 2644 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-79
transform 1 0 2599 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-80
transform 1 0 2402 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-81
transform 1 0 2102 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-82
transform 1 0 2114 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-83
transform 1 0 2113 0 1 2328
box 0 0 3 6
use FEEDTHRU  F-84
transform 1 0 2188 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-85
transform 1 0 2214 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-86
transform 1 0 2231 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-87
transform 1 0 2229 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-88
transform 1 0 2510 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-89
transform 1 0 2272 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-90
transform 1 0 2310 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-91
transform 1 0 2346 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-92
transform 1 0 2292 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-93
transform 1 0 2320 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-94
transform 1 0 2335 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-95
transform 1 0 2209 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-96
transform 1 0 2169 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-97
transform 1 0 2250 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-98
transform 1 0 2214 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-99
transform 1 0 2194 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-100
transform 1 0 2215 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-101
transform 1 0 2518 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-102
transform 1 0 2503 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-103
transform 1 0 2521 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-104
transform 1 0 2538 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-105
transform 1 0 2514 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-106
transform 1 0 2249 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-107
transform 1 0 2263 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-108
transform 1 0 2158 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-109
transform 1 0 2232 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-110
transform 1 0 2410 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-111
transform 1 0 2420 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-112
transform 1 0 2408 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-113
transform 1 0 2389 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-114
transform 1 0 2347 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-115
transform 1 0 2176 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-116
transform 1 0 2127 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-117
transform 1 0 2181 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-118
transform 1 0 2160 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-119
transform 1 0 2194 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-120
transform 1 0 2519 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-121
transform 1 0 2611 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-122
transform 1 0 2675 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-123
transform 1 0 2516 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-124
transform 1 0 2195 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-125
transform 1 0 2418 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-126
transform 1 0 2460 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-127
transform 1 0 2470 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-128
transform 1 0 2576 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-129
transform 1 0 2579 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-130
transform 1 0 2557 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-131
transform 1 0 2509 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-132
transform 1 0 2495 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-133
transform 1 0 2502 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-134
transform 1 0 2584 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-135
transform 1 0 2547 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-136
transform 1 0 2486 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-137
transform 1 0 2104 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-138
transform 1 0 2101 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-139
transform 1 0 2074 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-140
transform 1 0 2068 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-141
transform 1 0 2093 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-142
transform 1 0 2093 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-143
transform 1 0 2475 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-144
transform 1 0 2481 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-145
transform 1 0 2343 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-146
transform 1 0 2376 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-147
transform 1 0 2455 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-148
transform 1 0 2485 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-149
transform 1 0 2492 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-150
transform 1 0 2499 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-151
transform 1 0 2566 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-152
transform 1 0 2535 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-153
transform 1 0 2373 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-154
transform 1 0 2432 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-155
transform 1 0 2396 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-156
transform 1 0 2377 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-157
transform 1 0 2359 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-158
transform 1 0 2378 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-159
transform 1 0 2331 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-160
transform 1 0 2117 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-161
transform 1 0 2108 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-162
transform 1 0 2124 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-163
transform 1 0 2114 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-164
transform 1 0 2581 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-165
transform 1 0 2428 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-166
transform 1 0 2303 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-167
transform 1 0 2272 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-168
transform 1 0 2335 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-169
transform 1 0 2064 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-170
transform 1 0 2071 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-171
transform 1 0 2076 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-172
transform 1 0 2077 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-173
transform 1 0 2084 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-174
transform 1 0 2171 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-175
transform 1 0 2250 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-176
transform 1 0 2266 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-177
transform 1 0 2316 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-178
transform 1 0 2436 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-179
transform 1 0 2283 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-180
transform 1 0 2278 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-181
transform 1 0 2311 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-182
transform 1 0 2432 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-183
transform 1 0 2507 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-184
transform 1 0 2206 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-185
transform 1 0 2196 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-186
transform 1 0 2192 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-187
transform 1 0 2194 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-188
transform 1 0 2185 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-189
transform 1 0 2304 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-190
transform 1 0 2294 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-191
transform 1 0 2320 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-192
transform 1 0 2293 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-193
transform 1 0 2310 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-194
transform 1 0 2310 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-195
transform 1 0 2286 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-196
transform 1 0 2131 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-197
transform 1 0 2235 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-198
transform 1 0 2145 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-199
transform 1 0 2223 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-200
transform 1 0 2254 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-201
transform 1 0 2284 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-202
transform 1 0 2234 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-203
transform 1 0 2210 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-204
transform 1 0 2331 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-205
transform 1 0 2386 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-206
transform 1 0 2133 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-207
transform 1 0 2193 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-208
transform 1 0 2246 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-209
transform 1 0 2315 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-210
transform 1 0 2172 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-211
transform 1 0 2184 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-212
transform 1 0 2204 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-213
transform 1 0 2190 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-214
transform 1 0 2231 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-215
transform 1 0 2432 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-216
transform 1 0 2331 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-217
transform 1 0 2442 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-218
transform 1 0 2495 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-219
transform 1 0 2592 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-220
transform 1 0 2612 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-221
transform 1 0 2620 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-222
transform 1 0 2099 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-223
transform 1 0 2735 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-224
transform 1 0 2691 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-225
transform 1 0 2677 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-226
transform 1 0 2632 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-227
transform 1 0 2635 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-228
transform 1 0 2678 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-229
transform 1 0 2666 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-230
transform 1 0 2662 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-231
transform 1 0 2734 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-232
transform 1 0 2684 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-233
transform 1 0 2709 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-234
transform 1 0 2485 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-235
transform 1 0 2578 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-236
transform 1 0 2650 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-237
transform 1 0 2696 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-238
transform 1 0 2623 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-239
transform 1 0 2631 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-240
transform 1 0 2641 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-241
transform 1 0 2595 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-242
transform 1 0 2593 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-243
transform 1 0 2638 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-244
transform 1 0 2659 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-245
transform 1 0 2697 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-246
transform 1 0 2675 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-247
transform 1 0 2670 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-248
transform 1 0 2651 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-249
transform 1 0 2635 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-250
transform 1 0 2535 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-251
transform 1 0 2462 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-252
transform 1 0 2645 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-253
transform 1 0 2629 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-254
transform 1 0 2529 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-255
transform 1 0 2456 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-256
transform 1 0 2376 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-257
transform 1 0 2663 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-258
transform 1 0 2691 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-259
transform 1 0 2647 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-260
transform 1 0 2626 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-261
transform 1 0 2578 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-262
transform 1 0 2580 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-263
transform 1 0 2629 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-264
transform 1 0 2619 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-265
transform 1 0 2605 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-266
transform 1 0 2678 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-267
transform 1 0 2632 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-268
transform 1 0 2563 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-269
transform 1 0 2622 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-270
transform 1 0 2632 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-271
transform 1 0 2601 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-272
transform 1 0 2611 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-273
transform 1 0 2583 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-274
transform 1 0 2572 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-275
transform 1 0 2629 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-276
transform 1 0 2650 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-277
transform 1 0 2694 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-278
transform 1 0 2522 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-279
transform 1 0 2536 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-280
transform 1 0 2563 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-281
transform 1 0 2573 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-282
transform 1 0 2498 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-283
transform 1 0 2664 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-284
transform 1 0 2669 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-285
transform 1 0 2685 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-286
transform 1 0 2653 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-287
transform 1 0 2632 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-288
transform 1 0 2584 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-289
transform 1 0 2586 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-290
transform 1 0 2623 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-291
transform 1 0 2613 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-292
transform 1 0 2617 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-293
transform 1 0 2690 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-294
transform 1 0 2644 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-295
transform 1 0 2572 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-296
transform 1 0 2491 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-297
transform 1 0 2416 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-298
transform 1 0 2330 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-299
transform 1 0 2554 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-300
transform 1 0 2593 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-301
transform 1 0 2628 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-302
transform 1 0 2614 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-303
transform 1 0 2631 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-304
transform 1 0 2594 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-305
transform 1 0 2580 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-306
transform 1 0 2483 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-307
transform 1 0 2420 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-308
transform 1 0 2334 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-309
transform 1 0 2255 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-310
transform 1 0 2617 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-311
transform 1 0 2613 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-312
transform 1 0 2486 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-313
transform 1 0 2583 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-314
transform 1 0 2471 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-315
transform 1 0 2337 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-316
transform 1 0 2258 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-317
transform 1 0 2360 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-318
transform 1 0 2480 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-319
transform 1 0 2593 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-320
transform 1 0 2508 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-321
transform 1 0 2501 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-322
transform 1 0 2573 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-323
transform 1 0 2575 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-324
transform 1 0 2551 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-325
transform 1 0 2534 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-326
transform 1 0 2193 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-327
transform 1 0 2307 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-328
transform 1 0 2394 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-329
transform 1 0 2196 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-330
transform 1 0 2167 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-331
transform 1 0 2597 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-332
transform 1 0 2602 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-333
transform 1 0 2130 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-334
transform 1 0 2285 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-335
transform 1 0 2288 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-336
transform 1 0 2358 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-337
transform 1 0 2461 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-338
transform 1 0 2520 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-339
transform 1 0 2572 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-340
transform 1 0 2647 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-341
transform 1 0 2575 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-342
transform 1 0 2518 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-343
transform 1 0 2535 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-344
transform 1 0 2253 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-345
transform 1 0 2435 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-346
transform 1 0 2353 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-347
transform 1 0 2274 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-348
transform 1 0 2594 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-349
transform 1 0 2590 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-350
transform 1 0 2557 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-351
transform 1 0 2546 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-352
transform 1 0 2582 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-353
transform 1 0 2574 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-354
transform 1 0 2489 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-355
transform 1 0 2514 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-356
transform 1 0 2598 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-357
transform 1 0 2606 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-358
transform 1 0 2667 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-359
transform 1 0 2672 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-360
transform 1 0 2688 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-361
transform 1 0 2656 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-362
transform 1 0 2635 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-363
transform 1 0 2549 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-364
transform 1 0 2538 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-365
transform 1 0 2423 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-366
transform 1 0 2301 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-367
transform 1 0 2243 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-368
transform 1 0 2249 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-369
transform 1 0 2304 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-370
transform 1 0 2411 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-371
transform 1 0 2518 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-372
transform 1 0 2536 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-373
transform 1 0 2252 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-374
transform 1 0 2307 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-375
transform 1 0 2414 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-376
transform 1 0 2521 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-377
transform 1 0 2539 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-378
transform 1 0 2489 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-379
transform 1 0 2572 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-380
transform 1 0 2498 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-381
transform 1 0 2419 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-382
transform 1 0 2334 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-383
transform 1 0 2272 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-384
transform 1 0 2229 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-385
transform 1 0 2581 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-386
transform 1 0 2488 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-387
transform 1 0 2376 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-388
transform 1 0 2314 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-389
transform 1 0 2332 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-390
transform 1 0 2282 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-391
transform 1 0 2247 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-392
transform 1 0 2300 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-393
transform 1 0 2312 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-394
transform 1 0 2425 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-395
transform 1 0 2122 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-396
transform 1 0 2541 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-397
transform 1 0 2539 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-398
transform 1 0 2566 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-399
transform 1 0 2482 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-400
transform 1 0 2455 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-401
transform 1 0 2136 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-402
transform 1 0 2584 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-403
transform 1 0 2566 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-404
transform 1 0 2107 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-405
transform 1 0 2109 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-406
transform 1 0 2110 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-407
transform 1 0 2123 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-408
transform 1 0 2168 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-409
transform 1 0 2247 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-410
transform 1 0 2263 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-411
transform 1 0 2313 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-412
transform 1 0 2433 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-413
transform 1 0 2553 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-414
transform 1 0 2599 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-415
transform 1 0 2544 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-416
transform 1 0 2541 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-417
transform 1 0 2552 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-418
transform 1 0 2397 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-419
transform 1 0 2489 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-420
transform 1 0 2496 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-421
transform 1 0 2491 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-422
transform 1 0 2472 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-423
transform 1 0 2478 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-424
transform 1 0 2452 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-425
transform 1 0 2501 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-426
transform 1 0 2576 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-427
transform 1 0 2419 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-428
transform 1 0 2431 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-429
transform 1 0 2525 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-430
transform 1 0 2265 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-431
transform 1 0 2442 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-432
transform 1 0 2382 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-433
transform 1 0 2467 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-434
transform 1 0 2497 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-435
transform 1 0 2465 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-436
transform 1 0 2478 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-437
transform 1 0 2560 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-438
transform 1 0 2508 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-439
transform 1 0 2449 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-440
transform 1 0 2343 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-441
transform 1 0 2219 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-442
transform 1 0 2445 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-443
transform 1 0 2385 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-444
transform 1 0 2470 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-445
transform 1 0 2500 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-446
transform 1 0 2468 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-447
transform 1 0 2481 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-448
transform 1 0 2554 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-449
transform 1 0 2502 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-450
transform 1 0 2386 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-451
transform 1 0 2519 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-452
transform 1 0 2693 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-453
transform 1 0 2620 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-454
transform 1 0 2616 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-455
transform 1 0 2626 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-456
transform 1 0 2639 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-457
transform 1 0 2598 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-458
transform 1 0 2634 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-459
transform 1 0 2626 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-460
transform 1 0 2232 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-461
transform 1 0 2191 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-462
transform 1 0 2154 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-463
transform 1 0 2181 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-464
transform 1 0 2185 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-465
transform 1 0 2384 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-466
transform 1 0 2151 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-467
transform 1 0 2167 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-468
transform 1 0 2137 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-469
transform 1 0 2171 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-470
transform 1 0 2189 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-471
transform 1 0 2145 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-472
transform 1 0 2155 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-473
transform 1 0 2147 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-474
transform 1 0 2382 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-475
transform 1 0 2526 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-476
transform 1 0 2569 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-477
transform 1 0 2553 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-478
transform 1 0 2570 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-479
transform 1 0 2523 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-480
transform 1 0 2520 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-481
transform 1 0 2132 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-482
transform 1 0 2170 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-483
transform 1 0 2161 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-484
transform 1 0 2163 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-485
transform 1 0 2166 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-486
transform 1 0 2145 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-487
transform 1 0 2120 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-488
transform 1 0 2152 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-489
transform 1 0 2164 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-490
transform 1 0 2157 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-491
transform 1 0 2157 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-492
transform 1 0 2148 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-493
transform 1 0 2128 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-494
transform 1 0 2208 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-495
transform 1 0 2070 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-496
transform 1 0 2358 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-497
transform 1 0 2517 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-498
transform 1 0 2364 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-499
transform 1 0 2314 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-500
transform 1 0 2226 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-501
transform 1 0 2130 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-502
transform 1 0 2210 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-503
transform 1 0 2489 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-504
transform 1 0 2425 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-505
transform 1 0 2550 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-506
transform 1 0 2538 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-507
transform 1 0 2569 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-508
transform 1 0 2388 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-509
transform 1 0 2384 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-510
transform 1 0 2334 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-511
transform 1 0 2596 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-512
transform 1 0 2567 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-513
transform 1 0 2531 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-514
transform 1 0 2605 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-515
transform 1 0 2494 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-516
transform 1 0 2504 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-517
transform 1 0 2436 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-518
transform 1 0 2499 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-519
transform 1 0 2485 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-520
transform 1 0 2515 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-521
transform 1 0 2486 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-522
transform 1 0 2484 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-523
transform 1 0 2502 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-524
transform 1 0 2488 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-525
transform 1 0 2505 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-526
transform 1 0 2590 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-527
transform 1 0 2532 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-528
transform 1 0 2548 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-529
transform 1 0 2357 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-530
transform 1 0 2442 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-531
transform 1 0 2510 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-532
transform 1 0 2506 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-533
transform 1 0 2530 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-534
transform 1 0 2552 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-535
transform 1 0 2114 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-536
transform 1 0 2147 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-537
transform 1 0 2416 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-538
transform 1 0 2350 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-539
transform 1 0 2445 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-540
transform 1 0 2107 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-541
transform 1 0 2177 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-542
transform 1 0 2179 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-543
transform 1 0 2157 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-544
transform 1 0 2178 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-545
transform 1 0 2175 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-546
transform 1 0 2173 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-547
transform 1 0 2188 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-548
transform 1 0 2258 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-549
transform 1 0 2292 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-550
transform 1 0 2301 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-551
transform 1 0 2179 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-552
transform 1 0 2163 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-553
transform 1 0 2150 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-554
transform 1 0 2170 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-555
transform 1 0 2160 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-556
transform 1 0 2366 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-557
transform 1 0 2110 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-558
transform 1 0 2159 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-559
transform 1 0 2092 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-560
transform 1 0 2132 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-561
transform 1 0 2161 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-562
transform 1 0 2555 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-563
transform 1 0 2555 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-564
transform 1 0 2497 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-565
transform 1 0 2514 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-566
transform 1 0 2478 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-567
transform 1 0 2148 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-568
transform 1 0 2158 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-569
transform 1 0 2313 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-570
transform 1 0 2528 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-571
transform 1 0 2573 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-572
transform 1 0 2578 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-573
transform 1 0 2605 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-574
transform 1 0 2625 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-575
transform 1 0 2605 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-576
transform 1 0 2587 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-577
transform 1 0 2548 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-578
transform 1 0 2565 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-579
transform 1 0 2647 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-580
transform 1 0 2668 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-581
transform 1 0 2509 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-582
transform 1 0 2555 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-583
transform 1 0 2328 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-584
transform 1 0 2277 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-585
transform 1 0 2520 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-586
transform 1 0 2361 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-587
transform 1 0 2356 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-588
transform 1 0 2386 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-589
transform 1 0 2357 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-590
transform 1 0 2345 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-591
transform 1 0 2389 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-592
transform 1 0 2322 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-593
transform 1 0 2314 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-594
transform 1 0 2315 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-595
transform 1 0 2216 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-596
transform 1 0 2325 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-597
transform 1 0 2321 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-598
transform 1 0 2350 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-599
transform 1 0 2311 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-600
transform 1 0 2319 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-601
transform 1 0 2379 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-602
transform 1 0 2271 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-603
transform 1 0 2302 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-604
transform 1 0 2301 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-605
transform 1 0 2193 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-606
transform 1 0 2281 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-607
transform 1 0 2314 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-608
transform 1 0 2237 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-609
transform 1 0 2174 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-610
transform 1 0 2196 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-611
transform 1 0 2316 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-612
transform 1 0 2199 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-613
transform 1 0 2211 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-614
transform 1 0 2179 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-615
transform 1 0 2206 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-616
transform 1 0 2150 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-617
transform 1 0 2176 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-618
transform 1 0 2232 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-619
transform 1 0 2176 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-620
transform 1 0 2205 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-621
transform 1 0 2256 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-622
transform 1 0 2392 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-623
transform 1 0 2330 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-624
transform 1 0 2301 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-625
transform 1 0 2235 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-626
transform 1 0 2208 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-627
transform 1 0 2209 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-628
transform 1 0 2192 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-629
transform 1 0 2225 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-630
transform 1 0 2268 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-631
transform 1 0 2270 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-632
transform 1 0 2259 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-633
transform 1 0 2275 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-634
transform 1 0 2425 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-635
transform 1 0 2381 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-636
transform 1 0 2409 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-637
transform 1 0 2439 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-638
transform 1 0 2485 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-639
transform 1 0 2597 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-640
transform 1 0 2486 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-641
transform 1 0 2593 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-642
transform 1 0 2560 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-643
transform 1 0 2549 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-644
transform 1 0 2364 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-645
transform 1 0 2602 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-646
transform 1 0 2556 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-647
transform 1 0 2200 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-648
transform 1 0 2335 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-649
transform 1 0 2400 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-650
transform 1 0 2457 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-651
transform 1 0 2535 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-652
transform 1 0 2475 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-653
transform 1 0 2431 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-654
transform 1 0 2508 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-655
transform 1 0 2504 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-656
transform 1 0 2323 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-657
transform 1 0 2306 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-658
transform 1 0 2313 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-659
transform 1 0 2310 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-660
transform 1 0 2582 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-661
transform 1 0 2551 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-662
transform 1 0 2277 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-663
transform 1 0 2223 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-664
transform 1 0 2271 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-665
transform 1 0 2217 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-666
transform 1 0 2496 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-667
transform 1 0 2245 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-668
transform 1 0 2240 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-669
transform 1 0 2286 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-670
transform 1 0 2244 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-671
transform 1 0 2297 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-672
transform 1 0 2222 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-673
transform 1 0 2319 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-674
transform 1 0 2203 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-675
transform 1 0 2193 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-676
transform 1 0 2195 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-677
transform 1 0 2197 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-678
transform 1 0 2164 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-679
transform 1 0 2153 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-680
transform 1 0 2435 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-681
transform 1 0 2169 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-682
transform 1 0 2166 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-683
transform 1 0 2690 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-684
transform 1 0 2679 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-685
transform 1 0 2500 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-686
transform 1 0 2516 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-687
transform 1 0 2155 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-688
transform 1 0 2126 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-689
transform 1 0 2086 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-690
transform 1 0 2249 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-691
transform 1 0 2201 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-692
transform 1 0 2157 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-693
transform 1 0 2265 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-694
transform 1 0 2307 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-695
transform 1 0 2538 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-696
transform 1 0 2460 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-697
transform 1 0 2426 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-698
transform 1 0 2437 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-699
transform 1 0 2399 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-700
transform 1 0 2151 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-701
transform 1 0 2506 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-702
transform 1 0 2466 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-703
transform 1 0 2442 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-704
transform 1 0 2417 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-705
transform 1 0 2455 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-706
transform 1 0 2441 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-707
transform 1 0 2608 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-708
transform 1 0 2681 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-709
transform 1 0 2451 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-710
transform 1 0 2427 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-711
transform 1 0 2402 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-712
transform 1 0 2440 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-713
transform 1 0 2429 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-714
transform 1 0 2394 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-715
transform 1 0 2439 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-716
transform 1 0 2478 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-717
transform 1 0 2434 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-718
transform 1 0 2264 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-719
transform 1 0 2340 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-720
transform 1 0 2374 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-721
transform 1 0 2397 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-722
transform 1 0 2499 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-723
transform 1 0 2382 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-724
transform 1 0 2408 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-725
transform 1 0 2416 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-726
transform 1 0 2369 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-727
transform 1 0 2377 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-728
transform 1 0 2400 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-729
transform 1 0 2421 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-730
transform 1 0 2362 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-731
transform 1 0 2373 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-732
transform 1 0 2350 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-733
transform 1 0 2355 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-734
transform 1 0 2415 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-735
transform 1 0 2376 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-736
transform 1 0 2596 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-737
transform 1 0 2131 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-738
transform 1 0 2139 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-739
transform 1 0 2149 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-740
transform 1 0 2638 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-741
transform 1 0 2654 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-742
transform 1 0 2673 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-743
transform 1 0 2678 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-744
transform 1 0 2700 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-745
transform 1 0 2422 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-746
transform 1 0 2275 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-747
transform 1 0 2199 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-748
transform 1 0 2194 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-749
transform 1 0 2214 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-750
transform 1 0 2217 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-751
transform 1 0 2228 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-752
transform 1 0 2363 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-753
transform 1 0 2139 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-754
transform 1 0 2157 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-755
transform 1 0 2145 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-756
transform 1 0 2255 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-757
transform 1 0 2256 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-758
transform 1 0 2164 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-759
transform 1 0 2162 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-760
transform 1 0 2175 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-761
transform 1 0 2191 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-762
transform 1 0 2200 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-763
transform 1 0 2177 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-764
transform 1 0 2159 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-765
transform 1 0 2254 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-766
transform 1 0 2242 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-767
transform 1 0 2459 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-768
transform 1 0 2473 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-769
transform 1 0 2423 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-770
transform 1 0 2551 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-771
transform 1 0 2502 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-772
transform 1 0 2554 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-773
transform 1 0 2117 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-774
transform 1 0 2143 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-775
transform 1 0 2267 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-776
transform 1 0 2275 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-777
transform 1 0 2398 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-778
transform 1 0 2148 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-779
transform 1 0 2149 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-780
transform 1 0 2148 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-781
transform 1 0 2152 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-782
transform 1 0 2187 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-783
transform 1 0 2214 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-784
transform 1 0 2218 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-785
transform 1 0 2133 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-786
transform 1 0 2147 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-787
transform 1 0 2176 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-788
transform 1 0 2261 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-789
transform 1 0 2377 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-790
transform 1 0 2504 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-791
transform 1 0 2511 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-792
transform 1 0 2596 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-793
transform 1 0 2268 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-794
transform 1 0 2483 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-795
transform 1 0 2283 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-796
transform 1 0 2305 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-797
transform 1 0 2456 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-798
transform 1 0 2468 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-799
transform 1 0 2666 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-800
transform 1 0 2410 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-801
transform 1 0 2648 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-802
transform 1 0 2148 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-803
transform 1 0 2163 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-804
transform 1 0 2154 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-805
transform 1 0 2146 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-806
transform 1 0 2222 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-807
transform 1 0 2284 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-808
transform 1 0 2252 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-809
transform 1 0 2160 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-810
transform 1 0 2191 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-811
transform 1 0 2250 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-812
transform 1 0 2285 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-813
transform 1 0 2332 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-814
transform 1 0 2337 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-815
transform 1 0 2255 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-816
transform 1 0 2194 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-817
transform 1 0 2153 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-818
transform 1 0 2183 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-819
transform 1 0 2167 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-820
transform 1 0 2362 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-821
transform 1 0 2383 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-822
transform 1 0 2248 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-823
transform 1 0 2241 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-824
transform 1 0 2250 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-825
transform 1 0 2494 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-826
transform 1 0 2173 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-827
transform 1 0 2241 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-828
transform 1 0 2292 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-829
transform 1 0 2291 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-830
transform 1 0 2239 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-831
transform 1 0 2224 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-832
transform 1 0 2225 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-833
transform 1 0 2181 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-834
transform 1 0 2186 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-835
transform 1 0 2228 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-836
transform 1 0 2217 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-837
transform 1 0 2105 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-838
transform 1 0 2532 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-839
transform 1 0 2379 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-840
transform 1 0 2120 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-841
transform 1 0 2126 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-842
transform 1 0 2162 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-843
transform 1 0 2185 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-844
transform 1 0 2211 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-845
transform 1 0 2226 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-846
transform 1 0 2196 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-847
transform 1 0 2218 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-848
transform 1 0 2233 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-849
transform 1 0 2195 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-850
transform 1 0 2314 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-851
transform 1 0 2317 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-852
transform 1 0 2315 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-853
transform 1 0 2280 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-854
transform 1 0 2197 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-855
transform 1 0 2177 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-856
transform 1 0 2163 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-857
transform 1 0 2345 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-858
transform 1 0 2206 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-859
transform 1 0 2196 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-860
transform 1 0 2191 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-861
transform 1 0 2199 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-862
transform 1 0 2202 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-863
transform 1 0 2298 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-864
transform 1 0 2250 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-865
transform 1 0 2221 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-866
transform 1 0 2211 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-867
transform 1 0 2156 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-868
transform 1 0 2336 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-869
transform 1 0 2481 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-870
transform 1 0 2359 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-871
transform 1 0 2331 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-872
transform 1 0 2262 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-873
transform 1 0 2272 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-874
transform 1 0 2266 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-875
transform 1 0 2438 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-876
transform 1 0 2440 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-877
transform 1 0 2404 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-878
transform 1 0 2402 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-879
transform 1 0 2355 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-880
transform 1 0 2240 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-881
transform 1 0 2247 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-882
transform 1 0 2254 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-883
transform 1 0 2246 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-884
transform 1 0 2278 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-885
transform 1 0 2302 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-886
transform 1 0 2258 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-887
transform 1 0 2212 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-888
transform 1 0 2214 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-889
transform 1 0 2220 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-890
transform 1 0 2205 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-891
transform 1 0 2168 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-892
transform 1 0 2185 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-893
transform 1 0 2193 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-894
transform 1 0 2203 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-895
transform 1 0 2202 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-896
transform 1 0 2128 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-897
transform 1 0 2144 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-898
transform 1 0 2186 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-899
transform 1 0 2230 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-900
transform 1 0 2665 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-901
transform 1 0 2669 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-902
transform 1 0 2687 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-903
transform 1 0 2437 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-904
transform 1 0 2403 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-905
transform 1 0 2360 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-906
transform 1 0 2487 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-907
transform 1 0 2436 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-908
transform 1 0 2462 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-909
transform 1 0 2576 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-910
transform 1 0 2380 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-911
transform 1 0 2333 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-912
transform 1 0 2370 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-913
transform 1 0 2517 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-914
transform 1 0 2491 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-915
transform 1 0 2558 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-916
transform 1 0 2294 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-917
transform 1 0 2533 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-918
transform 1 0 2509 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-919
transform 1 0 2513 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-920
transform 1 0 2257 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-921
transform 1 0 2263 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-922
transform 1 0 2238 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-923
transform 1 0 2268 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-924
transform 1 0 2250 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-925
transform 1 0 2366 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-926
transform 1 0 2335 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-927
transform 1 0 2422 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-928
transform 1 0 2438 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-929
transform 1 0 2335 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-930
transform 1 0 2247 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-931
transform 1 0 2274 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-932
transform 1 0 2296 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-933
transform 1 0 2265 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-934
transform 1 0 2283 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-935
transform 1 0 2270 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-936
transform 1 0 2328 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-937
transform 1 0 2151 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-938
transform 1 0 2160 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-939
transform 1 0 2182 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-940
transform 1 0 2178 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-941
transform 1 0 2182 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-942
transform 1 0 2174 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-943
transform 1 0 2181 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-944
transform 1 0 2209 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-945
transform 1 0 2191 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-946
transform 1 0 2207 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-947
transform 1 0 2171 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-948
transform 1 0 2209 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-949
transform 1 0 2206 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-950
transform 1 0 2190 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-951
transform 1 0 2208 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-952
transform 1 0 2187 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-953
transform 1 0 2167 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-954
transform 1 0 2196 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-955
transform 1 0 2104 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-956
transform 1 0 2089 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-957
transform 1 0 2070 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-958
transform 1 0 2070 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-959
transform 1 0 2182 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-960
transform 1 0 2179 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-961
transform 1 0 2538 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-962
transform 1 0 2417 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-963
transform 1 0 2395 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-964
transform 1 0 2431 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-965
transform 1 0 2471 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-966
transform 1 0 2224 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-967
transform 1 0 2323 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-968
transform 1 0 2397 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-969
transform 1 0 2438 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-970
transform 1 0 2201 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-971
transform 1 0 2276 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-972
transform 1 0 2222 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-973
transform 1 0 2213 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-974
transform 1 0 2192 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-975
transform 1 0 2412 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-976
transform 1 0 2430 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-977
transform 1 0 2464 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-978
transform 1 0 2447 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-979
transform 1 0 2453 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-980
transform 1 0 2211 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-981
transform 1 0 2228 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-982
transform 1 0 2226 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-983
transform 1 0 2230 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-984
transform 1 0 2228 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-985
transform 1 0 2236 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-986
transform 1 0 2266 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-987
transform 1 0 2492 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-988
transform 1 0 2577 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-989
transform 1 0 2585 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-990
transform 1 0 2482 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-991
transform 1 0 2504 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-992
transform 1 0 2513 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-993
transform 1 0 2503 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-994
transform 1 0 2427 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-995
transform 1 0 2370 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-996
transform 1 0 2387 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-997
transform 1 0 2368 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-998
transform 1 0 2380 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-999
transform 1 0 2417 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1000
transform 1 0 2435 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1001
transform 1 0 2137 0 1 2028
box 0 0 3 6
use FEEDTHRU  F-1002
transform 1 0 2134 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-1003
transform 1 0 2166 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-1004
transform 1 0 2207 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-1005
transform 1 0 2180 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1006
transform 1 0 2235 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1007
transform 1 0 2233 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1008
transform 1 0 2262 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1009
transform 1 0 2283 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1010
transform 1 0 2271 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1011
transform 1 0 2302 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1012
transform 1 0 2299 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1013
transform 1 0 2276 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1014
transform 1 0 2307 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1015
transform 1 0 2292 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1016
transform 1 0 2332 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1017
transform 1 0 2296 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1018
transform 1 0 2492 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1019
transform 1 0 2219 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-1020
transform 1 0 2190 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-1021
transform 1 0 2170 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-1022
transform 1 0 2385 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1023
transform 1 0 2587 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1024
transform 1 0 2289 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1025
transform 1 0 2257 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1026
transform 1 0 2301 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1027
transform 1 0 2498 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1028
transform 1 0 2512 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1029
transform 1 0 2312 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1030
transform 1 0 2421 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1031
transform 1 0 2463 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1032
transform 1 0 2473 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1033
transform 1 0 2318 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1034
transform 1 0 2318 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1035
transform 1 0 2299 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1036
transform 1 0 2290 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1037
transform 1 0 2300 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1038
transform 1 0 2289 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1039
transform 1 0 2237 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1040
transform 1 0 2319 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1041
transform 1 0 2295 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1042
transform 1 0 2230 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1043
transform 1 0 2202 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1044
transform 1 0 2232 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1045
transform 1 0 2398 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1046
transform 1 0 2429 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1047
transform 1 0 2192 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1048
transform 1 0 2183 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-1049
transform 1 0 2174 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1050
transform 1 0 2191 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1051
transform 1 0 2285 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1052
transform 1 0 2171 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1053
transform 1 0 2194 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1054
transform 1 0 2229 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1055
transform 1 0 2246 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1056
transform 1 0 2244 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1057
transform 1 0 2260 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1058
transform 1 0 2264 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1059
transform 1 0 2272 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1060
transform 1 0 2290 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1061
transform 1 0 2361 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1062
transform 1 0 2268 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1063
transform 1 0 2285 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1064
transform 1 0 2348 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1065
transform 1 0 2402 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1066
transform 1 0 2398 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1067
transform 1 0 2487 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1068
transform 1 0 2511 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1069
transform 1 0 2575 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1070
transform 1 0 2501 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1071
transform 1 0 2641 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1072
transform 1 0 2430 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1073
transform 1 0 2387 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1074
transform 1 0 2486 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1075
transform 1 0 2373 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1076
transform 1 0 2343 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1077
transform 1 0 2317 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1078
transform 1 0 2316 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1079
transform 1 0 2337 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1080
transform 1 0 2364 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1081
transform 1 0 2379 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1082
transform 1 0 2422 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1083
transform 1 0 2287 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1084
transform 1 0 2292 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1085
transform 1 0 2293 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1086
transform 1 0 2298 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1087
transform 1 0 2225 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1088
transform 1 0 2228 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-1089
transform 1 0 2229 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1090
transform 1 0 2519 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1091
transform 1 0 2503 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1092
transform 1 0 2503 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1093
transform 1 0 2525 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1094
transform 1 0 2712 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1095
transform 1 0 2524 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1096
transform 1 0 2472 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1097
transform 1 0 2602 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1098
transform 1 0 2512 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1099
transform 1 0 2558 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1100
transform 1 0 2447 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1101
transform 1 0 2632 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1102
transform 1 0 2711 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1103
transform 1 0 2659 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1104
transform 1 0 2392 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1105
transform 1 0 2193 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1106
transform 1 0 2232 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1107
transform 1 0 2256 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1108
transform 1 0 2220 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1109
transform 1 0 2251 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1110
transform 1 0 2406 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1111
transform 1 0 2465 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1112
transform 1 0 2331 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1113
transform 1 0 2331 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1114
transform 1 0 2422 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1115
transform 1 0 2472 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1116
transform 1 0 2484 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1117
transform 1 0 2433 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1118
transform 1 0 2456 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1119
transform 1 0 2476 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1120
transform 1 0 2419 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1121
transform 1 0 2469 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1122
transform 1 0 2481 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1123
transform 1 0 2430 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1124
transform 1 0 2236 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1125
transform 1 0 2380 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1126
transform 1 0 2349 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1127
transform 1 0 2252 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1128
transform 1 0 2601 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1129
transform 1 0 2609 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1130
transform 1 0 2473 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1131
transform 1 0 2260 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1132
transform 1 0 2248 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1133
transform 1 0 2234 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1134
transform 1 0 2348 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1135
transform 1 0 2394 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1136
transform 1 0 2423 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1137
transform 1 0 2419 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1138
transform 1 0 2254 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1139
transform 1 0 2236 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1140
transform 1 0 2458 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1141
transform 1 0 2459 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1142
transform 1 0 2447 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1143
transform 1 0 2425 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1144
transform 1 0 2407 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1145
transform 1 0 2203 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-1146
transform 1 0 2501 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1147
transform 1 0 2479 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1148
transform 1 0 2521 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1149
transform 1 0 2543 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1150
transform 1 0 2552 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1151
transform 1 0 2557 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1152
transform 1 0 2505 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1153
transform 1 0 2466 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1154
transform 1 0 2223 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1155
transform 1 0 2229 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1156
transform 1 0 2397 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1157
transform 1 0 2367 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1158
transform 1 0 2409 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1159
transform 1 0 2272 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1160
transform 1 0 2228 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1161
transform 1 0 2283 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1162
transform 1 0 2307 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1163
transform 1 0 2259 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1164
transform 1 0 2290 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1165
transform 1 0 2183 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1166
transform 1 0 2227 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1167
transform 1 0 2205 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1168
transform 1 0 2220 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-1169
transform 1 0 2282 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1170
transform 1 0 2345 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1171
transform 1 0 2385 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1172
transform 1 0 2393 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1173
transform 1 0 2386 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1174
transform 1 0 2404 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1175
transform 1 0 2315 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1176
transform 1 0 2271 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1177
transform 1 0 2306 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1178
transform 1 0 2308 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1179
transform 1 0 2277 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1180
transform 1 0 2312 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1181
transform 1 0 2314 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1182
transform 1 0 2311 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1183
transform 1 0 2312 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1184
transform 1 0 2342 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1185
transform 1 0 2106 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-1186
transform 1 0 2101 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-1187
transform 1 0 2381 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1188
transform 1 0 2374 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1189
transform 1 0 2392 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1190
transform 1 0 2399 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1191
transform 1 0 2261 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1192
transform 1 0 2264 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1193
transform 1 0 2211 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-1194
transform 1 0 2356 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1195
transform 1 0 2369 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1196
transform 1 0 2375 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1197
transform 1 0 2423 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1198
transform 1 0 2275 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1199
transform 1 0 2269 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1200
transform 1 0 2225 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1201
transform 1 0 2262 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1202
transform 1 0 2143 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-1203
transform 1 0 2372 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1204
transform 1 0 2412 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1205
transform 1 0 2465 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1206
transform 1 0 2443 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1207
transform 1 0 2485 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1208
transform 1 0 2507 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1209
transform 1 0 2516 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1210
transform 1 0 2378 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1211
transform 1 0 2418 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1212
transform 1 0 2471 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1213
transform 1 0 2449 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1214
transform 1 0 2491 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1215
transform 1 0 2513 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1216
transform 1 0 2522 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1217
transform 1 0 2662 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1218
transform 1 0 2396 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1219
transform 1 0 2430 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1220
transform 1 0 2483 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1221
transform 1 0 2455 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1222
transform 1 0 2497 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1223
transform 1 0 2519 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1224
transform 1 0 2528 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1225
transform 1 0 2518 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1226
transform 1 0 2243 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1227
transform 1 0 2300 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1228
transform 1 0 2352 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1229
transform 1 0 2399 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1230
transform 1 0 2325 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1231
transform 1 0 2277 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1232
transform 1 0 2331 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1233
transform 1 0 2208 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-1234
transform 1 0 2255 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1235
transform 1 0 2318 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1236
transform 1 0 2364 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1237
transform 1 0 2313 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1238
transform 1 0 2333 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1239
transform 1 0 2396 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1240
transform 1 0 2320 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1241
transform 1 0 2271 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1242
transform 1 0 2280 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1243
transform 1 0 2330 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1244
transform 1 0 2336 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1245
transform 1 0 2326 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1246
transform 1 0 2277 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1247
transform 1 0 2557 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1248
transform 1 0 2474 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1249
transform 1 0 2459 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1250
transform 1 0 2443 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1251
transform 1 0 2244 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-1252
transform 1 0 2279 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1253
transform 1 0 2345 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1254
transform 1 0 2362 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1255
transform 1 0 2387 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1256
transform 1 0 2381 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1257
transform 1 0 2365 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1258
transform 1 0 2334 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1259
transform 1 0 2337 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1260
transform 1 0 2288 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1261
transform 1 0 2332 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1262
transform 1 0 2317 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1263
transform 1 0 2289 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1264
transform 1 0 2343 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1265
transform 1 0 2307 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1266
transform 1 0 2269 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1267
transform 1 0 2365 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1268
transform 1 0 2374 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1269
transform 1 0 2312 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1270
transform 1 0 2451 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1271
transform 1 0 2737 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1272
transform 1 0 2441 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1273
transform 1 0 2354 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1274
transform 1 0 2164 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-1275
transform 1 0 2175 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-1276
transform 1 0 2216 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-1277
transform 1 0 2310 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1278
transform 1 0 2163 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-1279
transform 1 0 2204 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-1280
transform 1 0 2228 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1281
transform 1 0 2225 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1282
transform 1 0 2291 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1283
transform 1 0 2316 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1284
transform 1 0 2357 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1285
transform 1 0 2350 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1286
transform 1 0 2368 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1287
transform 1 0 2393 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1288
transform 1 0 2387 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1289
transform 1 0 2216 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1290
transform 1 0 2282 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1291
transform 1 0 2322 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1292
transform 1 0 2369 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1293
transform 1 0 2356 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1294
transform 1 0 2374 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1295
transform 1 0 2222 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1296
transform 1 0 2288 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1297
transform 1 0 2328 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1298
transform 1 0 2375 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1299
transform 1 0 2354 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1300
transform 1 0 2338 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1301
transform 1 0 2296 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1302
transform 1 0 2323 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1303
transform 1 0 2336 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1304
transform 1 0 2330 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1305
transform 1 0 2308 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1306
transform 1 0 2231 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1307
transform 1 0 2281 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1308
transform 1 0 2635 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1309
transform 1 0 2406 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1310
transform 1 0 2449 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1311
transform 1 0 2465 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1312
transform 1 0 2316 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1313
transform 1 0 2301 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1314
transform 1 0 2264 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1315
transform 1 0 2317 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1316
transform 1 0 2699 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1317
transform 1 0 2653 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1318
transform 1 0 2395 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1319
transform 1 0 2304 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1320
transform 1 0 2349 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1321
transform 1 0 2380 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1322
transform 1 0 2421 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1323
transform 1 0 2451 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1324
transform 1 0 2400 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1325
transform 1 0 2295 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1326
transform 1 0 2339 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1327
transform 1 0 2320 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1328
transform 1 0 2344 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1329
transform 1 0 2360 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1330
transform 1 0 2360 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1331
transform 1 0 2338 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1332
transform 1 0 2298 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1333
transform 1 0 2289 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1334
transform 1 0 2255 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1335
transform 1 0 2305 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1336
transform 1 0 2453 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1337
transform 1 0 2435 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1338
transform 1 0 2413 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1339
transform 1 0 2261 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1340
transform 1 0 2375 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1341
transform 1 0 2424 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1342
transform 1 0 2448 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1343
transform 1 0 2500 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1344
transform 1 0 2510 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1345
transform 1 0 2501 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1346
transform 1 0 2479 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1347
transform 1 0 2372 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1348
transform 1 0 2344 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1349
transform 1 0 2304 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1350
transform 1 0 2429 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1351
transform 1 0 2413 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1352
transform 1 0 2370 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1353
transform 1 0 2334 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1354
transform 1 0 2389 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1355
transform 1 0 2352 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1356
transform 1 0 2325 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1357
transform 1 0 2282 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1358
transform 1 0 2329 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1359
transform 1 0 2314 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1360
transform 1 0 2295 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1361
transform 1 0 2355 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1362
transform 1 0 2319 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1363
transform 1 0 2275 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1364
transform 1 0 2253 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1365
transform 1 0 2210 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1366
transform 1 0 2395 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1367
transform 1 0 2358 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1368
transform 1 0 2347 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1369
transform 1 0 2252 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1370
transform 1 0 2349 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1371
transform 1 0 2390 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1372
transform 1 0 2529 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1373
transform 1 0 2359 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1374
transform 1 0 2322 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1375
transform 1 0 2273 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1376
transform 1 0 2457 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1377
transform 1 0 2393 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1378
transform 1 0 2377 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1379
transform 1 0 2346 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1380
transform 1 0 2340 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1381
transform 1 0 2178 0 1 2316
box 0 0 3 6
use FEEDTHRU  F-1382
transform 1 0 2279 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1383
transform 1 0 2342 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1384
transform 1 0 2382 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1385
transform 1 0 2429 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1386
transform 1 0 2413 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1387
transform 1 0 2449 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1388
transform 1 0 2465 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1389
transform 1 0 2480 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1390
transform 1 0 2328 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1391
transform 1 0 2319 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1392
transform 1 0 2459 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1393
transform 1 0 2325 0 1 2304
box 0 0 3 6
use FEEDTHRU  F-1394
transform 1 0 2390 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1395
transform 1 0 2424 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1396
transform 1 0 2632 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1397
transform 1 0 2356 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1398
transform 1 0 2353 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1399
transform 1 0 2334 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1400
transform 1 0 2385 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1401
transform 1 0 2361 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1402
transform 1 0 2311 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1403
transform 1 0 2289 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1404
transform 1 0 2246 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1405
transform 1 0 2198 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-1406
transform 1 0 2154 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-1407
transform 1 0 2304 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1408
transform 1 0 2329 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1409
transform 1 0 2379 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1410
transform 1 0 2403 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1411
transform 1 0 2352 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1412
transform 1 0 2473 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1413
transform 1 0 2515 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1414
transform 1 0 2537 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1415
transform 1 0 2546 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1416
transform 1 0 2536 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1417
transform 1 0 2484 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1418
transform 1 0 2460 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1419
transform 1 0 2494 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1420
transform 1 0 2437 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1421
transform 1 0 2401 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1422
transform 1 0 2394 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1423
transform 1 0 2506 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1424
transform 1 0 2521 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1425
transform 1 0 2225 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-1426
transform 1 0 2187 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-1427
transform 1 0 2173 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-1428
transform 1 0 2322 0 1 2076
box 0 0 3 6
use FEEDTHRU  F-1429
transform 1 0 2370 0 1 2088
box 0 0 3 6
use FEEDTHRU  F-1430
transform 1 0 2401 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1431
transform 1 0 2451 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1432
transform 1 0 2461 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1433
transform 1 0 2477 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1434
transform 1 0 2492 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1435
transform 1 0 2476 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1436
transform 1 0 2298 0 1 2064
box 0 0 3 6
use FEEDTHRU  F-1437
transform 1 0 2248 0 1 2052
box 0 0 3 6
use FEEDTHRU  F-1438
transform 1 0 2240 0 1 2040
box 0 0 3 6
use FEEDTHRU  F-1439
transform 1 0 2381 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1440
transform 1 0 2399 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1441
transform 1 0 2383 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1442
transform 1 0 2496 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1443
transform 1 0 2482 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1444
transform 1 0 2436 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1445
transform 1 0 2406 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1446
transform 1 0 2384 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1447
transform 1 0 2404 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1448
transform 1 0 2396 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1449
transform 1 0 2483 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1450
transform 1 0 2447 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1451
transform 1 0 2356 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1452
transform 1 0 2279 0 1 2292
box 0 0 3 6
use FEEDTHRU  F-1453
transform 1 0 2310 0 1 2280
box 0 0 3 6
use FEEDTHRU  F-1454
transform 1 0 2363 0 1 2268
box 0 0 3 6
use FEEDTHRU  F-1455
transform 1 0 2344 0 1 2256
box 0 0 3 6
use FEEDTHRU  F-1456
transform 1 0 2386 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1457
transform 1 0 2405 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1458
transform 1 0 2417 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1459
transform 1 0 2407 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1460
transform 1 0 2307 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1461
transform 1 0 2548 0 1 2244
box 0 0 3 6
use FEEDTHRU  F-1462
transform 1 0 2570 0 1 2232
box 0 0 3 6
use FEEDTHRU  F-1463
transform 1 0 2579 0 1 2220
box 0 0 3 6
use FEEDTHRU  F-1464
transform 1 0 2572 0 1 2208
box 0 0 3 6
use FEEDTHRU  F-1465
transform 1 0 2526 0 1 2196
box 0 0 3 6
use FEEDTHRU  F-1466
transform 1 0 2496 0 1 2184
box 0 0 3 6
use FEEDTHRU  F-1467
transform 1 0 2439 0 1 2172
box 0 0 3 6
use FEEDTHRU  F-1468
transform 1 0 2488 0 1 2160
box 0 0 3 6
use FEEDTHRU  F-1469
transform 1 0 2483 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1470
transform 1 0 2463 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1471
transform 1 0 2514 0 1 2124
box 0 0 3 6
use FEEDTHRU  F-1472
transform 1 0 2499 0 1 2112
box 0 0 3 6
use FEEDTHRU  F-1473
transform 1 0 2446 0 1 2100
box 0 0 3 6
use FEEDTHRU  F-1474
transform 1 0 2313 0 1 2136
box 0 0 3 6
use FEEDTHRU  F-1475
transform 1 0 2438 0 1 2148
box 0 0 3 6
use FEEDTHRU  F-1476
transform 1 0 2160 0 1 2052
box 0 0 3 6
<< end >>
