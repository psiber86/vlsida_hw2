magic
tech scmos
timestamp 1395738639
<< m1p >>
use CELL  1
transform -1 0 493 0 1 276
box 0 0 6 6
use CELL  2
transform -1 0 614 0 1 258
box 0 0 6 6
use CELL  3
transform -1 0 505 0 1 249
box 0 0 6 6
use CELL  4
transform -1 0 533 0 1 348
box 0 0 6 6
use CELL  5
transform -1 0 498 0 1 330
box 0 0 6 6
use CELL  6
transform -1 0 699 0 -1 318
box 0 0 6 6
use CELL  7
transform -1 0 555 0 1 294
box 0 0 6 6
use CELL  8
transform -1 0 522 0 1 231
box 0 0 6 6
use CELL  9
transform -1 0 532 0 1 267
box 0 0 6 6
use CELL  10
transform -1 0 549 0 1 348
box 0 0 6 6
use CELL  11
transform -1 0 526 0 1 285
box 0 0 6 6
use CELL  12
transform 1 0 726 0 1 303
box 0 0 6 6
use CELL  13
transform 1 0 666 0 -1 327
box 0 0 6 6
use CELL  14
transform -1 0 524 0 1 249
box 0 0 6 6
use CELL  15
transform -1 0 517 0 1 321
box 0 0 6 6
use CELL  16
transform -1 0 668 0 1 276
box 0 0 6 6
use CELL  17
transform -1 0 726 0 1 303
box 0 0 6 6
use CELL  18
transform -1 0 599 0 -1 345
box 0 0 6 6
use CELL  19
transform -1 0 499 0 1 348
box 0 0 6 6
use CELL  20
transform -1 0 719 0 1 303
box 0 0 6 6
use CELL  21
transform -1 0 734 0 1 312
box 0 0 6 6
use CELL  22
transform -1 0 531 0 -1 237
box 0 0 6 6
use CELL  23
transform 1 0 511 0 -1 255
box 0 0 6 6
use CELL  24
transform 1 0 506 0 -1 282
box 0 0 6 6
use CELL  25
transform -1 0 513 0 -1 291
box 0 0 6 6
use CELL  26
transform -1 0 624 0 1 321
box 0 0 6 6
use CELL  27
transform -1 0 720 0 1 267
box 0 0 6 6
use CELL  28
transform -1 0 512 0 1 294
box 0 0 6 6
use CELL  29
transform -1 0 688 0 1 294
box 0 0 6 6
use CELL  30
transform -1 0 517 0 1 240
box 0 0 6 6
use CELL  31
transform -1 0 750 0 1 267
box 0 0 6 6
use CELL  32
transform 1 0 620 0 -1 336
box 0 0 6 6
use CELL  33
transform -1 0 492 0 1 267
box 0 0 6 6
use CELL  34
transform -1 0 651 0 1 258
box 0 0 6 6
use CELL  35
transform 1 0 618 0 1 312
box 0 0 6 6
use CELL  36
transform -1 0 626 0 1 258
box 0 0 6 6
use CELL  37
transform -1 0 505 0 1 276
box 0 0 6 6
use CELL  38
transform -1 0 474 0 1 303
box 0 0 6 6
use CELL  39
transform -1 0 528 0 1 357
box 0 0 6 6
use CELL  40
transform -1 0 592 0 1 339
box 0 0 6 6
use CELL  41
transform -1 0 682 0 -1 282
box 0 0 6 6
use CELL  42
transform -1 0 480 0 1 285
box 0 0 6 6
use CELL  43
transform -1 0 544 0 1 276
box 0 0 6 6
use CELL  44
transform -1 0 543 0 1 321
box 0 0 6 6
use CELL  45
transform -1 0 512 0 1 258
box 0 0 6 6
use CELL  46
transform -1 0 481 0 1 303
box 0 0 6 6
use CELL  47
transform -1 0 520 0 1 285
box 0 0 6 6
use CELL  48
transform 1 0 669 0 1 312
box 0 0 6 6
use CELL  49
transform -1 0 696 0 1 276
box 0 0 6 6
use CELL  50
transform -1 0 499 0 1 321
box 0 0 6 6
use CELL  51
transform -1 0 705 0 1 303
box 0 0 6 6
use CELL  52
transform 1 0 697 0 -1 282
box 0 0 6 6
use CELL  53
transform -1 0 617 0 1 249
box 0 0 6 6
use CELL  54
transform -1 0 713 0 1 267
box 0 0 6 6
use CELL  55
transform -1 0 732 0 1 285
box 0 0 6 6
use CELL  56
transform -1 0 533 0 1 303
box 0 0 6 6
use CELL  57
transform -1 0 727 0 1 312
box 0 0 6 6
use CELL  58
transform -1 0 583 0 -1 345
box 0 0 6 6
use CELL  59
transform -1 0 608 0 1 249
box 0 0 6 6
use CELL  60
transform -1 0 525 0 1 267
box 0 0 6 6
use CELL  61
transform 1 0 595 0 -1 255
box 0 0 6 6
use CELL  62
transform 1 0 721 0 1 267
box 0 0 6 6
use CELL  63
transform -1 0 540 0 1 348
box 0 0 6 6
use CELL  64
transform 1 0 706 0 1 303
box 0 0 6 6
use CELL  65
transform -1 0 536 0 1 321
box 0 0 6 6
use CELL  66
transform 1 0 673 0 1 321
box 0 0 6 6
use CELL  67
transform 1 0 645 0 1 321
box 0 0 6 6
use CELL  68
transform -1 0 669 0 1 303
box 0 0 6 6
use CELL  69
transform -1 0 494 0 1 285
box 0 0 6 6
use CELL  70
transform -1 0 504 0 1 267
box 0 0 6 6
use CELL  71
transform -1 0 720 0 1 312
box 0 0 6 6
use CELL  72
transform -1 0 515 0 -1 354
box 0 0 6 6
use CELL  73
transform -1 0 639 0 1 321
box 0 0 6 6
use CELL  74
transform 1 0 533 0 -1 273
box 0 0 6 6
use CELL  75
transform -1 0 523 0 1 339
box 0 0 6 6
use CELL  76
transform -1 0 617 0 1 330
box 0 0 6 6
use CELL  77
transform -1 0 665 0 1 285
box 0 0 6 6
use CELL  78
transform -1 0 507 0 1 330
box 0 0 6 6
use CELL  79
transform 1 0 480 0 1 276
box 0 0 6 6
use CELL  80
transform -1 0 526 0 1 276
box 0 0 6 6
use CELL  81
transform -1 0 524 0 1 258
box 0 0 6 6
use CELL  82
transform -1 0 537 0 1 294
box 0 0 6 6
use CELL  83
transform -1 0 552 0 1 231
box 0 0 6 6
use CELL  84
transform -1 0 642 0 1 330
box 0 0 6 6
use CELL  85
transform -1 0 521 0 -1 354
box 0 0 6 6
use CELL  86
transform -1 0 492 0 1 321
box 0 0 6 6
use CELL  87
transform -1 0 487 0 1 285
box 0 0 6 6
use CELL  88
transform -1 0 532 0 1 339
box 0 0 6 6
use CELL  89
transform -1 0 487 0 1 303
box 0 0 6 6
use CELL  90
transform -1 0 510 0 1 240
box 0 0 6 6
use CELL  91
transform -1 0 739 0 1 303
box 0 0 6 6
use CELL  92
transform -1 0 746 0 1 285
box 0 0 6 6
use CELL  93
transform -1 0 526 0 1 303
box 0 0 6 6
use CELL  94
transform 1 0 611 0 1 303
box 0 0 6 6
use CELL  95
transform -1 0 503 0 1 312
box 0 0 6 6
use CELL  96
transform -1 0 517 0 -1 372
box 0 0 6 6
use CELL  97
transform -1 0 675 0 1 276
box 0 0 6 6
use CELL  98
transform -1 0 489 0 1 312
box 0 0 6 6
use CELL  99
transform -1 0 508 0 1 348
box 0 0 6 6
use CELL  100
transform 1 0 551 0 -1 255
box 0 0 6 6
use CELL  101
transform -1 0 576 0 1 258
box 0 0 6 6
use CELL  102
transform -1 0 492 0 1 339
box 0 0 6 6
use CELL  103
transform -1 0 512 0 1 303
box 0 0 6 6
use CELL  104
transform -1 0 505 0 1 258
box 0 0 6 6
use CELL  105
transform 1 0 550 0 1 348
box 0 0 6 6
use CELL  106
transform 1 0 636 0 1 258
box 0 0 6 6
use CELL  107
transform -1 0 551 0 1 276
box 0 0 6 6
use CELL  108
transform 1 0 687 0 1 321
box 0 0 6 6
use CELL  109
transform 1 0 700 0 1 312
box 0 0 6 6
use CELL  110
transform 1 0 512 0 -1 273
box 0 0 6 6
use CELL  111
transform -1 0 528 0 1 294
box 0 0 6 6
use CELL  112
transform -1 0 578 0 1 249
box 0 0 6 6
use CELL  113
transform -1 0 686 0 1 267
box 0 0 6 6
use CELL  114
transform 1 0 504 0 1 366
box 0 0 6 6
use CELL  115
transform -1 0 533 0 -1 291
box 0 0 6 6
use CELL  116
transform -1 0 663 0 1 321
box 0 0 6 6
use CELL  117
transform -1 0 548 0 -1 246
box 0 0 6 6
use CELL  118
transform -1 0 757 0 1 267
box 0 0 6 6
use CELL  119
transform -1 0 493 0 1 294
box 0 0 6 6
use CELL  120
transform 1 0 740 0 -1 309
box 0 0 6 6
use CELL  121
transform -1 0 531 0 1 258
box 0 0 6 6
use CELL  122
transform -1 0 565 0 1 339
box 0 0 6 6
use CELL  123
transform 1 0 656 0 1 303
box 0 0 6 6
use CELL  124
transform -1 0 639 0 1 294
box 0 0 6 6
use CELL  125
transform 1 0 733 0 1 285
box 0 0 6 6
use CELL  126
transform -1 0 521 0 1 294
box 0 0 6 6
use CELL  127
transform 1 0 492 0 -1 264
box 0 0 6 6
use CELL  128
transform 1 0 586 0 -1 255
box 0 0 6 6
use CELL  129
transform -1 0 671 0 1 267
box 0 0 6 6
use CELL  130
transform -1 0 505 0 1 294
box 0 0 6 6
use CELL  131
transform 1 0 505 0 -1 273
box 0 0 6 6
use CELL  132
transform -1 0 635 0 1 285
box 0 0 6 6
use CELL  133
transform -1 0 681 0 1 294
box 0 0 6 6
use CELL  134
transform -1 0 724 0 1 294
box 0 0 6 6
use CELL  135
transform -1 0 663 0 1 312
box 0 0 6 6
use CELL  136
transform -1 0 498 0 1 249
box 0 0 6 6
use CELL  137
transform -1 0 607 0 1 258
box 0 0 6 6
use CELL  138
transform -1 0 506 0 1 285
box 0 0 6 6
use CELL  139
transform -1 0 496 0 1 303
box 0 0 6 6
use CELL  140
transform -1 0 524 0 1 240
box 0 0 6 6
use CELL  141
transform -1 0 492 0 1 348
box 0 0 6 6
use CELL  142
transform -1 0 533 0 -1 336
box 0 0 6 6
use CELL  143
transform -1 0 635 0 1 258
box 0 0 6 6
use CELL  144
transform -1 0 486 0 1 294
box 0 0 6 6
use CELL  145
transform -1 0 749 0 1 294
box 0 0 6 6
use CELL  146
transform -1 0 583 0 1 258
box 0 0 6 6
use CELL  147
transform 1 0 680 0 1 321
box 0 0 6 6
use CELL  148
transform -1 0 526 0 1 330
box 0 0 6 6
use CELL  149
transform -1 0 743 0 1 267
box 0 0 6 6
use CELL  150
transform -1 0 736 0 1 267
box 0 0 6 6
use CELL  151
transform -1 0 765 0 1 294
box 0 0 6 6
use CELL  152
transform -1 0 519 0 1 330
box 0 0 6 6
use CELL  153
transform -1 0 496 0 1 312
box 0 0 6 6
use CELL  154
transform -1 0 531 0 1 312
box 0 0 6 6
use CELL  155
transform 1 0 557 0 -1 354
box 0 0 6 6
use CELL  156
transform 1 0 591 0 -1 246
box 0 0 6 6
use CELL  157
transform 1 0 707 0 1 312
box 0 0 6 6
use CELL  158
transform -1 0 524 0 1 312
box 0 0 6 6
use CELL  159
transform -1 0 585 0 1 249
box 0 0 6 6
use CELL  160
transform -1 0 689 0 1 276
box 0 0 6 6
use CELL  161
transform -1 0 604 0 1 240
box 0 0 6 6
use CELL  162
transform -1 0 529 0 1 321
box 0 0 6 6
use CELL  163
transform -1 0 504 0 1 339
box 0 0 6 6
use CELL  164
transform 1 0 474 0 1 312
box 0 0 6 6
use CELL  165
transform -1 0 590 0 1 240
box 0 0 6 6
use CELL  166
transform -1 0 517 0 1 312
box 0 0 6 6
use CELL  167
transform 1 0 643 0 1 330
box 0 0 6 6
use CELL  168
transform -1 0 753 0 -1 291
box 0 0 6 6
use CELL  169
transform -1 0 620 0 1 276
box 0 0 6 6
use CELL  170
transform -1 0 519 0 1 276
box 0 0 6 6
use CELL  171
transform -1 0 635 0 1 330
box 0 0 6 6
use CELL  172
transform -1 0 758 0 1 294
box 0 0 6 6
use CELL  173
transform -1 0 505 0 1 303
box 0 0 6 6
use CELL  174
transform 1 0 513 0 1 303
box 0 0 6 6
use CELL  175
transform 1 0 641 0 1 285
box 0 0 6 6
use CELL  176
transform 1 0 529 0 -1 363
box 0 0 6 6
use CELL  177
transform -1 0 725 0 1 285
box 0 0 6 6
use CELL  178
transform -1 0 731 0 1 294
box 0 0 6 6
use CELL  179
transform -1 0 510 0 1 312
box 0 0 6 6
use CELL  180
transform -1 0 511 0 1 339
box 0 0 6 6
<< metal1 >>
rect 512 310 513 313
rect 487 310 513 311
rect 487 310 488 312
rect 756 283 757 295
rect 751 283 757 284
rect 751 283 752 285
rect 637 292 638 295
rect 637 292 657 293
rect 657 292 658 303
rect 528 301 529 304
rect 528 301 631 302
rect 631 292 632 302
rect 631 292 636 293
rect 636 265 637 293
rect 636 265 715 266
rect 715 265 716 267
rect 530 337 531 340
rect 524 337 531 338
rect 524 337 525 346
rect 519 346 525 347
rect 519 346 520 348
rect 673 310 674 313
rect 673 310 676 311
rect 676 310 677 319
rect 670 319 677 320
rect 670 317 671 320
rect 633 256 634 259
rect 466 256 634 257
rect 466 256 467 328
rect 466 328 534 329
rect 534 328 535 346
rect 531 346 535 347
rect 531 346 532 348
rect 731 265 732 268
rect 731 265 738 266
rect 738 265 739 267
rect 576 229 577 250
rect 526 229 577 230
rect 526 229 527 231
rect 741 274 742 286
rect 701 274 742 275
rect 701 274 702 276
rect 660 274 661 286
rect 660 274 666 275
rect 666 274 667 276
rect 630 328 631 331
rect 627 328 631 329
rect 627 328 628 337
rect 627 337 644 338
rect 644 335 645 338
rect 521 301 522 304
rect 513 301 522 302
rect 513 292 514 302
rect 507 292 514 293
rect 507 292 508 294
rect 533 355 534 358
rect 533 355 584 356
rect 584 337 585 356
rect 584 337 590 338
rect 590 337 591 339
rect 760 292 761 295
rect 760 292 766 293
rect 766 292 767 301
rect 724 301 767 302
rect 724 301 725 303
rect 494 292 495 304
rect 494 292 503 293
rect 503 292 504 294
rect 502 265 503 268
rect 490 265 503 266
rect 490 265 491 267
rect 485 283 486 286
rect 478 283 486 284
rect 478 265 479 284
rect 478 265 487 266
rect 487 265 488 267
rect 481 292 482 295
rect 469 292 482 293
rect 469 292 470 303
rect 602 238 603 241
rect 580 238 603 239
rect 580 238 581 249
rect 527 319 528 322
rect 527 319 538 320
rect 538 319 539 321
rect 563 319 564 340
rect 541 319 564 320
rect 541 319 542 321
rect 633 283 634 286
rect 553 283 634 284
rect 553 283 554 294
rect 503 346 504 349
rect 497 346 504 347
rect 497 346 498 348
rect 676 292 677 295
rect 670 292 677 293
rect 670 292 671 310
rect 664 310 671 311
rect 664 310 665 319
rect 661 319 665 320
rect 661 319 662 321
rect 755 256 756 268
rect 649 256 756 257
rect 649 256 650 258
rect 660 308 661 310
rect 655 310 661 311
rect 655 310 656 319
rect 655 319 658 320
rect 658 319 659 321
rect 612 227 613 250
rect 523 227 613 228
rect 523 227 524 238
rect 515 238 524 239
rect 515 238 516 240
rect 502 337 503 340
rect 502 337 512 338
rect 512 337 513 346
rect 510 346 513 347
rect 510 346 511 348
rect 718 310 719 313
rect 718 310 729 311
rect 729 310 730 312
<< metal2 >>
rect 478 317 479 319
rect 466 319 479 320
rect 466 301 467 320
rect 466 301 472 302
rect 472 301 473 303
rect 499 328 500 340
rect 499 328 514 329
rect 514 328 515 330
rect 615 274 616 277
rect 615 274 663 275
rect 663 274 664 276
rect 496 247 497 250
rect 496 247 506 248
rect 506 247 507 256
rect 503 256 507 257
rect 503 256 504 258
rect 515 310 516 313
rect 515 310 532 311
rect 532 310 533 319
rect 521 319 533 320
rect 521 319 522 328
rect 521 328 531 329
rect 531 328 532 330
rect 711 265 712 268
rect 552 265 712 266
rect 552 265 553 292
rect 544 292 553 293
rect 544 292 545 346
rect 523 346 545 347
rect 523 346 524 357
rect 574 256 575 259
rect 525 256 575 257
rect 525 247 526 257
rect 515 247 526 248
rect 515 247 516 249
rect 491 310 492 313
rect 481 310 492 311
rect 481 310 482 319
rect 481 319 490 320
rect 490 319 491 321
rect 578 256 579 259
rect 578 256 593 257
rect 593 247 594 257
rect 526 247 594 248
rect 526 238 527 248
rect 490 238 527 239
rect 490 238 491 265
rect 490 265 534 266
rect 534 265 535 267
rect 748 283 749 286
rect 748 283 763 284
rect 763 283 764 294
rect 737 301 738 304
rect 727 301 738 302
rect 727 301 728 303
rect 634 292 635 295
rect 566 292 635 293
rect 566 292 567 364
rect 464 364 567 365
rect 464 292 465 365
rect 464 292 535 293
rect 535 292 536 294
<< end >>
